/* Verilog module written by vlog2Verilog (qflow) */

module cpu(
    output [15:0] AB,
    input [7:0] DI,
    output [7:0] DO,
    input IRQ,
    input NMI,
    input RDY,
    output WE,
    input clk,
    input reset
);

wire vdd = 1'b1;
wire gnd = 1'b0;

wire C ;
wire D ;
wire I ;
wire N ;
wire V ;
wire Z ;
wire _1257_ ;
wire _588_ ;
wire _168_ ;
wire _800_ ;
wire _60_ ;
wire _1486_ ;
wire _1066_ ;
wire _397_ ;
wire _1295_ ;
wire _703_ ;
wire _1389_ ;
wire _19_ ;
wire _1601_ ;
wire _932_ ;
wire _512_ ;
wire _1198_ ;
wire _1410_ ;
wire _741_ ;
wire _321_ ;
wire _57_ ;
wire _970_ ;
wire _550_ ;
wire _130_ ;
wire _606_ ;
wire _1504_ ;
wire _835_ ;
wire _415_ ;
wire _95_ ;
wire _1313_ ;
wire _644_ ;
wire _224_ ;
wire _1542_ ;
wire _1122_ ;
wire _873_ ;
wire _453_ ;
wire _929_ ;
wire _509_ ;
wire _1351_ ;
wire _682_ ;
wire _262_ ;
wire _1407_ ;
wire _738_ ;
wire _318_ ;
wire _1580_ ;
wire _1160_ ;
wire _491_ ;
wire _1636_ ;
wire _1216_ ;
wire _967_ ;
wire _547_ ;
wire _127_ ;
wire _1445_ ;
wire _1025_ ;
wire _776_ ;
wire _356_ ;
wire _1254_ ;
wire _585_ ;
wire _165_ ;
wire _1483_ ;
wire _1063_ ;
wire _394_ ;
wire _1539_ ;
wire _1119_ ;
wire _1292_ ;
wire _1348_ ;
wire _679_ ;
wire _259_ ;
wire _1577_ ;
wire _1157_ ;
wire _488_ ;
wire _700_ ;
wire _1386_ ;
wire _297_ ;
wire _16_ ;
wire _1195_ ;
wire _54_ ;
wire _603_ ;
wire _1289_ ;
wire _1501_ ;
wire _832_ ;
wire _412_ ;
wire _92_ ;
wire _1098_ ;
wire _1310_ ;
wire _641_ ;
wire _221_ ;
wire _870_ ;
wire _450_ ;
wire _926_ ;
wire _506_ ;
wire _1404_ ;
wire _735_ ;
wire _315_ ;
wire _1633_ ;
wire _1213_ ;
wire _964_ ;
wire _544_ ;
wire _124_ ;
wire IRQ ;
wire _1442_ ;
wire _1022_ ;
wire _773_ ;
wire _353_ ;
wire _829_ ;
wire _409_ ;
wire _89_ ;
wire _1251_ ;
wire _582_ ;
wire _162_ ;
wire _1307_ ;
wire _638_ ;
wire _218_ ;
wire _1480_ ;
wire _1060_ ;
wire _391_ ;
wire _1536_ ;
wire _1116_ ;
wire _867_ ;
wire _447_ ;
wire _1345_ ;
wire _676_ ;
wire _256_ ;
wire _1__bF$buf10 ;
wire _1574_ ;
wire _1154_ ;
wire _485_ ;
wire WE ;
wire _1383_ ;
wire _294_ ;
wire _13_ ;
wire _1439_ ;
wire _1019_ ;
wire php ;
wire _1192_ ;
wire _1248_ ;
wire _999_ ;
wire _579_ ;
wire _159_ ;
wire _51_ ;
wire _1477_ ;
wire _1057_ ;
wire _388_ ;
wire _600_ ;
wire _1286_ ;
wire _197_ ;
wire _1095_ ;
wire _7_ ;
wire RDY ;
wire _923_ ;
wire _503_ ;
wire _1189_ ;
wire _1401_ ;
wire _732_ ;
wire _312_ ;
wire adc_sbc ;
wire _48_ ;
wire _1630_ ;
wire _1210_ ;
wire _961_ ;
wire _541_ ;
wire _121_ ;
wire _770_ ;
wire _350_ ;
wire _826_ ;
wire _406_ ;
wire _86_ ;
wire _1304_ ;
wire _635_ ;
wire _215_ ;
wire _1533_ ;
wire _1113_ ;
wire _864_ ;
wire _444_ ;
wire _1342_ ;
wire _673_ ;
wire _253_ ;
wire _729_ ;
wire _309_ ;
wire _1571_ ;
wire _1151_ ;
wire _482_ ;
wire _1627_ ;
wire _1207_ ;
wire _958_ ;
wire _538_ ;
wire _118_ ;
wire _1380_ ;
wire _291_ ;
wire _10_ ;
wire _1436_ ;
wire _1016_ ;
wire _767_ ;
wire _347_ ;
wire [15:0] _1665_ ;
wire _1245_ ;
wire _996_ ;
wire _576_ ;
wire _156_ ;
wire _1474_ ;
wire _1054_ ;
wire _385_ ;
wire _1283_ ;
wire _194_ ;
wire _1339_ ;
wire _1092_ ;
wire _1568_ ;
wire _1148_ ;
wire _899_ ;
wire _479_ ;
wire write_back ;
wire _1377_ ;
wire _288_ ;
wire _4_ ;
wire _920_ ;
wire _500_ ;
wire _1186_ ;
wire _45_ ;
wire _823_ ;
wire _403_ ;
wire _83_ ;
wire _1089_ ;
wire _1301_ ;
wire _632_ ;
wire _212_ ;
wire _1530_ ;
wire _1110_ ;
wire _861_ ;
wire _441_ ;
wire _917_ ;
wire _670_ ;
wire _250_ ;
wire _726_ ;
wire _306_ ;
wire \ALU.right  ;
wire _1624_ ;
wire _1204_ ;
wire _955_ ;
wire _535_ ;
wire _115_ ;
wire _1433_ ;
wire _1013_ ;
wire _764_ ;
wire _344_ ;
wire _1662_ ;
wire _1242_ ;
wire _993_ ;
wire _573_ ;
wire _153_ ;
wire _629_ ;
wire _209_ ;
wire _1471_ ;
wire _1051_ ;
wire _382_ ;
wire _1527_ ;
wire _1107_ ;
wire _858_ ;
wire _438_ ;
wire _1280_ ;
wire _191_ ;
wire _1336_ ;
wire _667_ ;
wire _247_ ;
wire _1565_ ;
wire _1145_ ;
wire _896_ ;
wire _476_ ;
wire clk_bF$buf0 ;
wire clk_bF$buf1 ;
wire clk_bF$buf2 ;
wire clk_bF$buf3 ;
wire clk_bF$buf4 ;
wire clk_bF$buf5 ;
wire clk_bF$buf6 ;
wire clk_bF$buf7 ;
wire clk_bF$buf8 ;
wire clk_bF$buf9 ;
wire _1374_ ;
wire _285_ ;
wire _1_ ;
wire index_y ;
wire _1183_ ;
wire _1659_ ;
wire _1239_ ;
wire _42_ ;
wire _1468_ ;
wire _1048_ ;
wire _799_ ;
wire _379_ ;
wire _1277_ ;
wire _188_ ;
wire _820_ ;
wire _400_ ;
wire _80_ ;
wire _1086_ ;
wire _914_ ;
wire _723_ ;
wire _303_ ;
wire _39_ ;
wire _1621_ ;
wire _1201_ ;
wire _952_ ;
wire _532_ ;
wire _112_ ;
wire _1430_ ;
wire _1010_ ;
wire _761_ ;
wire _341_ ;
wire clc ;
wire cld ;
wire cli ;
wire clk ;
wire clv ;
wire _817_ ;
wire _77_ ;
wire _990_ ;
wire _570_ ;
wire _150_ ;
wire _626_ ;
wire _206_ ;
wire _1524_ ;
wire _1104_ ;
wire _855_ ;
wire _435_ ;
wire _1333_ ;
wire _664_ ;
wire _244_ ;
wire _1562_ ;
wire _1142_ ;
wire _893_ ;
wire _473_ ;
wire _1618_ ;
wire _949_ ;
wire _529_ ;
wire _109_ ;
wire _1371_ ;
wire _282_ ;
wire _1427_ ;
wire _1007_ ;
wire _758_ ;
wire _338_ ;
wire _1180_ ;
wire _1656_ ;
wire _1236_ ;
wire _987_ ;
wire _567_ ;
wire _147_ ;
wire _1465_ ;
wire _1045_ ;
wire _796_ ;
wire _376_ ;
wire _1274_ ;
wire _185_ ;
wire _1083_ ;
wire _1559_ ;
wire _1139_ ;
wire _1368_ ;
wire _699_ ;
wire _279_ ;
wire _911_ ;
wire _1597_ ;
wire _1177_ ;
wire _720_ ;
wire _300_ ;
wire _36_ ;
wire _814_ ;
wire _74_ ;
wire _623_ ;
wire _203_ ;
wire _1521_ ;
wire _1101_ ;
wire _852_ ;
wire _432_ ;
wire _908_ ;
wire _1330_ ;
wire _661_ ;
wire _241_ ;
wire \ALU.CO  ;
wire _717_ ;
wire _890_ ;
wire _470_ ;
wire _1615_ ;
wire _946_ ;
wire _526_ ;
wire _106_ ;
wire _1424_ ;
wire _1004_ ;
wire _755_ ;
wire _335_ ;
wire _1653_ ;
wire _1233_ ;
wire _984_ ;
wire _564_ ;
wire _144_ ;
wire _1462_ ;
wire _1042_ ;
wire _793_ ;
wire _373_ ;
wire _1518_ ;
wire _849_ ;
wire _429_ ;
wire _1271_ ;
wire _182_ ;
wire _1327_ ;
wire _658_ ;
wire _238_ ;
wire _1080_ ;
wire _1556_ ;
wire _1136_ ;
wire _887_ ;
wire _467_ ;
wire _1365_ ;
wire _696_ ;
wire _276_ ;
wire _1594_ ;
wire _1174_ ;
wire _33_ ;
wire _1459_ ;
wire _1039_ ;
wire \ALU.HC  ;
wire _1268_ ;
wire _599_ ;
wire _179_ ;
wire _811_ ;
wire _71_ ;
wire _1497_ ;
wire _1077_ ;
wire _620_ ;
wire _200_ ;
wire _905_ ;
wire _714_ ;
wire [7:0] ADD ;
wire _1612_ ;
wire _943_ ;
wire _523_ ;
wire _103_ ;
wire _1421_ ;
wire _1001_ ;
wire _752_ ;
wire _332_ ;
wire _808_ ;
wire _68_ ;
wire _1650_ ;
wire _1230_ ;
wire _981_ ;
wire _561_ ;
wire _141_ ;
wire _617_ ;
wire _790_ ;
wire _370_ ;
wire _1515_ ;
wire _846_ ;
wire _426_ ;
wire _1324_ ;
wire _655_ ;
wire _235_ ;
wire _1553_ ;
wire _1133_ ;
wire _884_ ;
wire _464_ ;
wire _1609_ ;
wire _1362_ ;
wire RDY_bF$buf0 ;
wire RDY_bF$buf1 ;
wire RDY_bF$buf2 ;
wire RDY_bF$buf3 ;
wire RDY_bF$buf4 ;
wire RDY_bF$buf5 ;
wire RDY_bF$buf6 ;
wire RDY_bF$buf7 ;
wire RDY_bF$buf8 ;
wire _693_ ;
wire _273_ ;
wire _1418_ ;
wire _749_ ;
wire _329_ ;
wire _1591_ ;
wire _1171_ ;
wire _1647_ ;
wire _1227_ ;
wire _978_ ;
wire _558_ ;
wire _138_ ;
wire _30_ ;
wire _1456_ ;
wire _1036_ ;
wire res ;
wire _787_ ;
wire _367_ ;
wire rotate ;
wire _1265_ ;
wire _596_ ;
wire _176_ ;
wire _1494_ ;
wire _1074_ ;
wire _836__bF$buf0 ;
wire _836__bF$buf1 ;
wire _836__bF$buf2 ;
wire _836__bF$buf3 ;
wire _836__bF$buf4 ;
wire _836__bF$buf5 ;
wire _836__bF$buf6 ;
wire _836__bF$buf7 ;
wire _1359_ ;
wire _902_ ;
wire _1588_ ;
wire _1168_ ;
wire _499_ ;
wire \ALU.CI  ;
wire _711_ ;
wire _1397_ ;
wire _27_ ;
wire _940_ ;
wire _520_ ;
wire _100_ ;
wire [1:0] dst_reg ;
wire [7:0] DIHOLD ;
wire _805_ ;
wire _65_ ;
wire _614_ ;
wire _1512_ ;
wire _843_ ;
wire _423_ ;
wire _1321_ ;
wire _652_ ;
wire _232_ ;
wire _708_ ;
wire _1550_ ;
wire _1130_ ;
wire _881_ ;
wire _461_ ;
wire _1606_ ;
wire _937_ ;
wire _517_ ;
wire _690_ ;
wire _270_ ;
wire _1415_ ;
wire _746_ ;
wire _326_ ;
wire _1644_ ;
wire _1224_ ;
wire _975_ ;
wire _555_ ;
wire _135_ ;
wire _1453_ ;
wire _1033_ ;
wire _784_ ;
wire _364_ ;
wire _1509_ ;
wire _1262_ ;
wire _593_ ;
wire _173_ ;
wire _1318_ ;
wire _649_ ;
wire _229_ ;
wire _1491_ ;
wire _1071_ ;
wire _1547_ ;
wire _1127_ ;
wire _878_ ;
wire _458_ ;
wire _1356_ ;
wire _687_ ;
wire _267_ ;
wire _1585_ ;
wire _1165_ ;
wire _496_ ;
wire _1394_ ;
wire _24_ ;
wire _1259_ ;
wire _802_ ;
wire _62_ ;
wire _1488_ ;
wire _1068_ ;
wire _399_ ;
wire _611_ ;
wire _1297_ ;
wire _840_ ;
wire _420_ ;
wire _705_ ;
wire _1603_ ;
wire _934_ ;
wire _514_ ;
wire _1412_ ;
wire _743_ ;
wire _323_ ;
wire _59_ ;
wire _1641_ ;
wire _1221_ ;
wire _972_ ;
wire _552_ ;
wire _132_ ;
wire _608_ ;
wire _1450_ ;
wire _1030_ ;
wire _781_ ;
wire _361_ ;
wire _1506_ ;
wire _837_ ;
wire _417_ ;
wire _97_ ;
wire _590_ ;
wire _170_ ;
wire _1315_ ;
wire _646_ ;
wire _226_ ;
wire _1544_ ;
wire _1124_ ;
wire _875_ ;
wire _455_ ;
wire _1353_ ;
wire _684_ ;
wire _264_ ;
wire [3:0] \ALU.op  ;
wire _1409_ ;
wire _1582_ ;
wire _1162_ ;
wire _493_ ;
wire _1638_ ;
wire _1218_ ;
wire _969_ ;
wire _549_ ;
wire _129_ ;
wire _1391_ ;
wire _21_ ;
wire _1447_ ;
wire _1027_ ;
wire _778_ ;
wire _358_ ;
wire _1256_ ;
wire _587_ ;
wire _167_ ;
wire _1485_ ;
wire _1065_ ;
wire _396_ ;
wire _1294_ ;
wire [7:0] \AXYS[1]  ;
wire _1579_ ;
wire _1159_ ;
wire _702_ ;
wire _1388_ ;
wire _299_ ;
wire _18_ ;
wire _1600_ ;
wire _931_ ;
wire _511_ ;
wire _1197_ ;
wire _740_ ;
wire _320_ ;
wire _56_ ;
wire _605_ ;
wire _1503_ ;
wire _834_ ;
wire _414_ ;
wire _94_ ;
wire _1312_ ;
wire _643_ ;
wire _223_ ;
wire _1541_ ;
wire _1121_ ;
wire _872_ ;
wire _452_ ;
wire _928_ ;
wire _508_ ;
wire _1350_ ;
wire _681_ ;
wire _261_ ;
wire _1406_ ;
wire _737_ ;
wire _317_ ;
wire _490_ ;
wire _1635_ ;
wire _1215_ ;
wire _966_ ;
wire _546_ ;
wire _126_ ;
wire _1444_ ;
wire _1024_ ;
wire _775_ ;
wire _355_ ;
wire _1253_ ;
wire _584_ ;
wire _164_ ;
wire _1309_ ;
wire _1482_ ;
wire _1062_ ;
wire _393_ ;
wire _1538_ ;
wire _1118_ ;
wire _869_ ;
wire _449_ ;
wire _1291_ ;
wire _1347_ ;
wire _678_ ;
wire _258_ ;
wire _1576_ ;
wire _1156_ ;
wire _487_ ;
wire _1385_ ;
wire _296_ ;
wire _15_ ;
wire _1194_ ;
wire _53_ ;
wire _1479_ ;
wire _1059_ ;
wire store ;
wire _602_ ;
wire _1288_ ;
wire _199_ ;
wire _1500_ ;
wire _831_ ;
wire _411_ ;
wire _91_ ;
wire _1097_ ;
wire _640_ ;
wire _220_ ;
wire _9_ ;
wire _925_ ;
wire _505_ ;
wire IRHOLD_valid ;
wire _1403_ ;
wire _734_ ;
wire _314_ ;
wire _1632_ ;
wire _1212_ ;
wire _963_ ;
wire _543_ ;
wire _123_ ;
wire _1441_ ;
wire _1021_ ;
wire _772_ ;
wire _352_ ;
wire _828_ ;
wire _408_ ;
wire _88_ ;
wire _1250_ ;
wire _581_ ;
wire _161_ ;
wire _1306_ ;
wire _637_ ;
wire _217_ ;
wire _390_ ;
wire _1535_ ;
wire _1115_ ;
wire _866_ ;
wire _446_ ;
wire _1344_ ;
wire _675_ ;
wire _255_ ;
wire _1573_ ;
wire _1153_ ;
wire _484_ ;
wire _1629_ ;
wire _1209_ ;
wire _1382_ ;
wire _293_ ;
wire _12_ ;
wire _1438_ ;
wire _1018_ ;
wire _769_ ;
wire _349_ ;
wire _1191_ ;
wire _1667_ ;
wire _1247_ ;
wire _998_ ;
wire _578_ ;
wire _158_ ;
wire _50_ ;
wire _1476_ ;
wire _1056_ ;
wire _387_ ;
wire _1285_ ;
wire _196_ ;
wire _1094_ ;
wire _856__bF$buf0 ;
wire _856__bF$buf1 ;
wire _856__bF$buf2 ;
wire _856__bF$buf3 ;
wire _860__bF$buf0 ;
wire _860__bF$buf1 ;
wire _860__bF$buf2 ;
wire _860__bF$buf3 ;
wire _860__bF$buf4 ;
wire _1379_ ;
wire _6_ ;
wire _922_ ;
wire _502_ ;
wire _1188_ ;
wire _1400_ ;
wire _731_ ;
wire _311_ ;
wire _47_ ;
wire _960_ ;
wire _540_ ;
wire _120_ ;
wire _825_ ;
wire _405_ ;
wire _85_ ;
wire _1303_ ;
wire _634_ ;
wire _214_ ;
wire _1532_ ;
wire _1112_ ;
wire _863_ ;
wire _443_ ;
wire _1__bF$buf0 ;
wire _1__bF$buf1 ;
wire _1__bF$buf2 ;
wire _1__bF$buf3 ;
wire _1__bF$buf4 ;
wire _1__bF$buf5 ;
wire _1__bF$buf6 ;
wire _1__bF$buf7 ;
wire _1__bF$buf8 ;
wire _1__bF$buf9 ;
wire _919_ ;
wire _1341_ ;
wire _672_ ;
wire _252_ ;
wire _728_ ;
wire _308_ ;
wire _1570_ ;
wire _1150_ ;
wire _481_ ;
wire _1626_ ;
wire _1206_ ;
wire _957_ ;
wire _537_ ;
wire _117_ ;
wire _290_ ;
wire _1435_ ;
wire _1015_ ;
wire _766_ ;
wire _346_ ;
wire _1664_ ;
wire _1244_ ;
wire _995_ ;
wire _575_ ;
wire _155_ ;
wire backwards ;
wire _1473_ ;
wire _1053_ ;
wire _384_ ;
wire _1529_ ;
wire _1109_ ;
wire _1282_ ;
wire _193_ ;
wire _1338_ ;
wire _669_ ;
wire _249_ ;
wire _1091_ ;
wire _1567_ ;
wire _1147_ ;
wire _898_ ;
wire _478_ ;
wire _1376_ ;
wire _287_ ;
wire _3_ ;
wire _1185_ ;
wire _859__bF$buf0 ;
wire _859__bF$buf1 ;
wire _859__bF$buf2 ;
wire _859__bF$buf3 ;
wire _44_ ;
wire _1279_ ;
wire _822_ ;
wire _402_ ;
wire _82_ ;
wire _1088_ ;
wire _1300_ ;
wire _631_ ;
wire _211_ ;
wire _860_ ;
wire _440_ ;
wire _916_ ;
wire _725_ ;
wire _305_ ;
wire [15:0] PC ;
wire _1623_ ;
wire _1203_ ;
wire _954_ ;
wire _534_ ;
wire _114_ ;
wire _1432_ ;
wire _1012_ ;
wire _763_ ;
wire _343_ ;
wire _819_ ;
wire _79_ ;
wire _1661_ ;
wire _1241_ ;
wire _992_ ;
wire _572_ ;
wire _152_ ;
wire _628_ ;
wire _208_ ;
wire _1470_ ;
wire _1050_ ;
wire _381_ ;
wire _1526_ ;
wire _1106_ ;
wire _857_ ;
wire _437_ ;
wire _190_ ;
wire _1335_ ;
wire _666_ ;
wire _246_ ;
wire _1564_ ;
wire _1144_ ;
wire _895_ ;
wire _475_ ;
wire _1373_ ;
wire _284_ ;
wire _0_ ;
wire _1429_ ;
wire _1009_ ;
wire _1182_ ;
wire _1658_ ;
wire _1238_ ;
wire _989_ ;
wire _569_ ;
wire _149_ ;
wire adj_bcd ;
wire _41_ ;
wire _1467_ ;
wire _1047_ ;
wire _798_ ;
wire _378_ ;
wire _1276_ ;
wire _187_ ;
wire _1085_ ;
wire _913_ ;
wire [7:0] \AXYS[3]  ;
wire _1599_ ;
wire _1179_ ;
wire _722_ ;
wire _302_ ;
wire _38_ ;
wire _1620_ ;
wire _1200_ ;
wire _951_ ;
wire _531_ ;
wire _111_ ;
wire _760_ ;
wire _340_ ;
wire compare ;
wire _816_ ;
wire _76_ ;
wire _625_ ;
wire _205_ ;
wire load_only ;
wire clk_bF$buf10 ;
wire shift ;
wire _1523_ ;
wire _1103_ ;
wire _854_ ;
wire _434_ ;
wire _1332_ ;
wire _663_ ;
wire _243_ ;
wire _719_ ;
wire _1561_ ;
wire _1141_ ;
wire _892_ ;
wire _472_ ;
wire _1617_ ;
wire _948_ ;
wire _528_ ;
wire _108_ ;
wire _1370_ ;
wire _281_ ;
wire _1426_ ;
wire _1006_ ;
wire _757_ ;
wire _337_ ;
wire _1655_ ;
wire _1235_ ;
wire _986_ ;
wire _566_ ;
wire _146_ ;
wire [1:0] src_reg ;
wire _1464_ ;
wire _1044_ ;
wire _795_ ;
wire _375_ ;
wire _1273_ ;
wire _184_ ;
wire _1329_ ;
wire _1082_ ;
wire _1558_ ;
wire _1138_ ;
wire _889_ ;
wire _469_ ;
wire _1367_ ;
wire _698_ ;
wire _278_ ;
wire _910_ ;
wire _1596_ ;
wire _1176_ ;
wire _35_ ;
wire _813_ ;
wire _73_ ;
wire _1499_ ;
wire _1079_ ;
wire _622_ ;
wire _202_ ;
wire _1520_ ;
wire _1100_ ;
wire _851_ ;
wire _431_ ;
wire _907_ ;
wire _660_ ;
wire _240_ ;
wire _716_ ;
wire _1614_ ;
wire _945_ ;
wire _525_ ;
wire _105_ ;
wire _1423_ ;
wire _1003_ ;
wire _754_ ;
wire _334_ ;
wire _1652_ ;
wire _1232_ ;
wire _983_ ;
wire _563_ ;
wire _143_ ;
wire _619_ ;
wire _1461_ ;
wire _1041_ ;
wire _792_ ;
wire _372_ ;
wire _1517_ ;
wire _848_ ;
wire _428_ ;
wire _1270_ ;
wire _181_ ;
wire _1326_ ;
wire _657_ ;
wire _237_ ;
wire _1555_ ;
wire _1135_ ;
wire _886_ ;
wire _466_ ;
wire _1364_ ;
wire _695_ ;
wire _275_ ;
wire _1593_ ;
wire _1173_ ;
wire _1649_ ;
wire _1229_ ;
wire \ALU.Z  ;
wire _32_ ;
wire _1458_ ;
wire _1038_ ;
wire [2:0] cond_code ;
wire _789_ ;
wire _369_ ;
wire _1267_ ;
wire _598_ ;
wire _178_ ;
wire _810_ ;
wire _70_ ;
wire _1496_ ;
wire _1076_ ;
wire _904_ ;
wire _713_ ;
wire _1399_ ;
wire _29_ ;
wire _1611_ ;
wire _942_ ;
wire _522_ ;
wire _102_ ;
wire _1420_ ;
wire _1000_ ;
wire _751_ ;
wire _331_ ;
wire _807_ ;
wire _67_ ;
wire _980_ ;
wire _560_ ;
wire _140_ ;
wire _616_ ;
wire [5:0] state ;
wire _1514_ ;
wire _845_ ;
wire _425_ ;
wire _1323_ ;
wire _654_ ;
wire _234_ ;
wire bit_ins ;
wire _1552_ ;
wire _1132_ ;
wire _883_ ;
wire _463_ ;
wire _1608_ ;
wire _939_ ;
wire _519_ ;
wire _1361_ ;
wire _692_ ;
wire _272_ ;
wire _1417_ ;
wire _748_ ;
wire _328_ ;
wire _1590_ ;
wire _1170_ ;
wire _1646_ ;
wire _1226_ ;
wire _977_ ;
wire _557_ ;
wire _137_ ;
wire [7:0] DI ;
wire [7:0] DO ;
wire _1455_ ;
wire _1035_ ;
wire _786_ ;
wire _366_ ;
wire _1264_ ;
wire _595_ ;
wire _175_ ;
wire _1493_ ;
wire _1073_ ;
wire _1549_ ;
wire _1129_ ;
wire _1358_ ;
wire _689_ ;
wire _269_ ;
wire _901_ ;
wire _1587_ ;
wire _1167_ ;
wire _498_ ;
wire _710_ ;
wire _1396_ ;
wire _26_ ;
wire \ALU.BI7  ;
wire _804_ ;
wire _64_ ;
wire _613_ ;
wire _1299_ ;
wire _1511_ ;
wire _842_ ;
wire _422_ ;
wire _1320_ ;
wire _651_ ;
wire _231_ ;
wire _707_ ;
wire _880_ ;
wire _460_ ;
wire _1605_ ;
wire _936_ ;
wire _516_ ;
wire _1414_ ;
wire _745_ ;
wire _325_ ;
wire _1643_ ;
wire _1223_ ;
wire _974_ ;
wire _554_ ;
wire _134_ ;
wire [15:0] AB ;
wire [7:0] AI ;
wire _1452_ ;
wire _1032_ ;
wire _783_ ;
wire _363_ ;
wire _1508_ ;
wire _839_ ;
wire _419_ ;
wire _99_ ;
wire _1261_ ;
wire _592_ ;
wire _172_ ;
wire _1317_ ;
wire _648_ ;
wire _228_ ;
wire _1490_ ;
wire _1070_ ;
wire _1546_ ;
wire _1126_ ;
wire _877_ ;
wire _457_ ;
wire _1355_ ;
wire _686_ ;
wire _266_ ;
wire _1584_ ;
wire _1164_ ;
wire _495_ ;
wire _1393_ ;
wire _23_ ;
wire _1449_ ;
wire _1029_ ;
wire _1258_ ;
wire _589_ ;
wire _169_ ;
wire _801_ ;
wire _61_ ;
wire _1487_ ;
wire _1067_ ;
wire _398_ ;
wire _610_ ;
wire _1296_ ;
wire \ALU.AI7  ;
wire _704_ ;
wire _815__bF$buf0 ;
wire _815__bF$buf1 ;
wire _815__bF$buf2 ;
wire _815__bF$buf3 ;
wire _815__bF$buf4 ;
wire _1602_ ;
wire _933_ ;
wire _513_ ;
wire _1199_ ;
wire _1411_ ;
wire _742_ ;
wire _322_ ;
wire _58_ ;
wire _1640_ ;
wire _1220_ ;
wire _971_ ;
wire _551_ ;
wire _131_ ;
wire _607_ ;
wire _780_ ;
wire _360_ ;
wire _1505_ ;
wire _836_ ;
wire _416_ ;
wire _96_ ;
wire NMI ;
wire _1314_ ;
wire _645_ ;
wire _225_ ;
wire \ALU.BCD  ;
wire _1543_ ;
wire _1123_ ;
wire _874_ ;
wire _454_ ;
wire _1352_ ;
wire _683_ ;
wire _263_ ;
wire _1408_ ;
wire _739_ ;
wire _319_ ;
wire _1581_ ;
wire _1161_ ;
wire _492_ ;
wire _1637_ ;
wire _1217_ ;
wire _968_ ;
wire _548_ ;
wire _128_ ;
wire _1390_ ;
wire _20_ ;
wire _1446_ ;
wire _1026_ ;
wire _777_ ;
wire _357_ ;
wire _1255_ ;
wire _586_ ;
wire _166_ ;
wire _1484_ ;
wire _1064_ ;
wire _395_ ;
wire _1293_ ;
wire _1349_ ;
wire _1578_ ;
wire _1158_ ;
wire _489_ ;
wire [7:0] \ALU.BI  ;
wire _701_ ;
wire _1387_ ;
wire _298_ ;
wire _17_ ;
wire _930_ ;
wire _510_ ;
wire plp ;
wire _1196_ ;
wire _55_ ;
wire \ALU.N  ;
wire _604_ ;
wire _1502_ ;
wire _833_ ;
wire _413_ ;
wire _93_ ;
wire _1099_ ;
wire _1311_ ;
wire _642_ ;
wire _222_ ;
wire _1540_ ;
wire _1120_ ;
wire _871_ ;
wire _451_ ;
wire _927_ ;
wire _507_ ;
wire _680_ ;
wire _260_ ;
wire _1405_ ;
wire _736_ ;
wire _316_ ;
wire _1634_ ;
wire _1214_ ;
wire _965_ ;
wire _545_ ;
wire _125_ ;
wire _1443_ ;
wire _1023_ ;
wire _774_ ;
wire _354_ ;
wire _1252_ ;
wire _583_ ;
wire _163_ ;
wire _1308_ ;
wire _639_ ;
wire _219_ ;
wire _1481_ ;
wire _1061_ ;
wire _392_ ;
wire _1537_ ;
wire _1117_ ;
wire _868_ ;
wire _448_ ;
wire _1290_ ;
wire _1346_ ;
wire _677_ ;
wire _257_ ;
wire _1575_ ;
wire _1155_ ;
wire _486_ ;
wire _1384_ ;
wire _295_ ;
wire _14_ ;
wire _1193_ ;
wire _1249_ ;
wire _52_ ;
wire _1478_ ;
wire _1058_ ;
wire _389_ ;
wire _1629__bF$buf0 ;
wire _1629__bF$buf1 ;
wire _1629__bF$buf2 ;
wire _1629__bF$buf3 ;
wire _601_ ;
wire _1287_ ;
wire _198_ ;
wire _830_ ;
wire _410_ ;
wire _90_ ;
wire _1096_ ;
wire _8_ ;
wire _924_ ;
wire _504_ ;
wire _1402_ ;
wire _733_ ;
wire _313_ ;
wire _923__bF$buf0 ;
wire _923__bF$buf1 ;
wire _923__bF$buf2 ;
wire _923__bF$buf3 ;
wire _49_ ;
wire _1631_ ;
wire _1211_ ;
wire _962_ ;
wire _542_ ;
wire _122_ ;
wire _1440_ ;
wire _1020_ ;
wire _771_ ;
wire _351_ ;
wire _827_ ;
wire _407_ ;
wire _87_ ;
wire _580_ ;
wire _160_ ;
wire _1305_ ;
wire _636_ ;
wire _216_ ;
wire _1534_ ;
wire _1114_ ;
wire _865_ ;
wire _445_ ;
wire _1343_ ;
wire _674_ ;
wire _254_ ;
wire _1572_ ;
wire _1152_ ;
wire _483_ ;
wire _1628_ ;
wire _1208_ ;
wire _959_ ;
wire _539_ ;
wire _119_ ;
wire _1381_ ;
wire _292_ ;
wire _11_ ;
wire _1437_ ;
wire _1017_ ;
wire _768_ ;
wire _348_ ;
wire _1190_ ;
wire [7:0] _1666_ ;
wire _1246_ ;
wire _997_ ;
wire _577_ ;
wire _157_ ;
wire _1475_ ;
wire _1055_ ;
wire _386_ ;
wire _1284_ ;
wire _195_ ;
wire _1093_ ;
wire [7:0] \AXYS[0]  ;
wire _1569_ ;
wire _1149_ ;
wire _1378_ ;
wire _289_ ;
wire _5_ ;
wire _921_ ;
wire _501_ ;
wire _1187_ ;
wire _730_ ;
wire _310_ ;
wire _899__bF$buf0 ;
wire _899__bF$buf1 ;
wire _899__bF$buf2 ;
wire _899__bF$buf3 ;
wire _899__bF$buf4 ;
wire _46_ ;
wire _824_ ;
wire _404_ ;
wire _84_ ;
wire _1302_ ;
wire _633_ ;
wire _213_ ;
wire _1531_ ;
wire _1111_ ;
wire _862_ ;
wire _442_ ;
wire _918_ ;
wire _1340_ ;
wire _671_ ;
wire _251_ ;
wire _727_ ;
wire _307_ ;
wire _480_ ;
wire _1625_ ;
wire _1205_ ;
wire _956_ ;
wire _536_ ;
wire _116_ ;
wire _1434_ ;
wire _1014_ ;
wire _765_ ;
wire _345_ ;
wire _1663_ ;
wire _1243_ ;
wire _994_ ;
wire _574_ ;
wire _154_ ;
wire _1472_ ;
wire _1052_ ;
wire _383_ ;
wire _1528_ ;
wire _1108_ ;
wire shift_right ;
wire _859_ ;
wire _439_ ;
wire _1281_ ;
wire _192_ ;
wire _1337_ ;
wire _668_ ;
wire _248_ ;
wire _1090_ ;
wire _1566_ ;
wire _1146_ ;
wire _897_ ;
wire _477_ ;
wire _1375_ ;
wire _286_ ;
wire _2_ ;
wire _1184_ ;
wire _43_ ;
wire _1469_ ;
wire _1049_ ;
wire [7:0] DIMUX ;
wire _1278_ ;
wire _189_ ;
wire _821_ ;
wire _401_ ;
wire _81_ ;
wire _1087_ ;
wire [3:0] op ;
wire _630_ ;
wire _210_ ;
wire _915_ ;
wire _724_ ;
wire _304_ ;
wire _1622_ ;
wire _1202_ ;
wire _953_ ;
wire _533_ ;
wire _113_ ;
wire _1431_ ;
wire _1011_ ;
wire _762_ ;
wire _342_ ;
wire _818_ ;
wire _78_ ;
wire _1660_ ;
wire _1240_ ;
wire _991_ ;
wire _571_ ;
wire _151_ ;
wire _627_ ;
wire _207_ ;
wire _380_ ;
wire _1525_ ;
wire _1105_ ;
wire _856_ ;
wire _436_ ;
wire _1334_ ;
wire _665_ ;
wire _245_ ;
wire _1563_ ;
wire _1143_ ;
wire _894_ ;
wire _474_ ;
wire _1619_ ;
wire _854__bF$buf0 ;
wire _854__bF$buf1 ;
wire _854__bF$buf2 ;
wire _854__bF$buf3 ;
wire _1372_ ;
wire _283_ ;
wire _1428_ ;
wire _1008_ ;
wire _759_ ;
wire _339_ ;
wire _1181_ ;
wire _1657_ ;
wire _1237_ ;
wire _988_ ;
wire _568_ ;
wire _148_ ;
wire _40_ ;
wire sec ;
wire sed ;
wire sei ;
wire _1466_ ;
wire _1046_ ;
wire _797_ ;
wire _377_ ;
wire [7:0] IRHOLD ;
wire _1275_ ;
wire _186_ ;
wire _1084_ ;
wire _917__bF$buf0 ;
wire _917__bF$buf1 ;
wire _917__bF$buf2 ;
wire _917__bF$buf3 ;
wire _917__bF$buf4 ;
wire _1369_ ;
wire _912_ ;
wire _1598_ ;
wire _1178_ ;
wire _721_ ;
wire _301_ ;
wire _37_ ;
wire _950_ ;
wire _530_ ;
wire _110_ ;
wire _815_ ;
wire _75_ ;
wire _624_ ;
wire _204_ ;
wire _1522_ ;
wire _1102_ ;
wire _853_ ;
wire _433_ ;
wire _1074__bF$buf0 ;
wire _1074__bF$buf1 ;
wire _1074__bF$buf2 ;
wire _1074__bF$buf3 ;
wire _909_ ;
wire _1331_ ;
wire _662_ ;
wire _242_ ;
wire _718_ ;
wire _1560_ ;
wire _1140_ ;
wire _891_ ;
wire _471_ ;
wire _1616_ ;
wire _947_ ;
wire _527_ ;
wire _107_ ;
wire _280_ ;
wire _1425_ ;
wire _1005_ ;
wire _756_ ;
wire _336_ ;
wire _1654_ ;
wire _1234_ ;
wire _985_ ;
wire _565_ ;
wire _145_ ;
wire [5:0] _1463_ ;
wire _1043_ ;
wire _794_ ;
wire _374_ ;
wire _1519_ ;
wire _1272_ ;
wire _861__bF$buf0 ;
wire _861__bF$buf1 ;
wire _861__bF$buf2 ;
wire _183_ ;
wire _861__bF$buf3 ;
wire _1328_ ;
wire _659_ ;
wire _239_ ;
wire _1081_ ;
wire _1557_ ;
wire _1137_ ;
wire _888_ ;
wire _468_ ;
wire _1366_ ;
wire _697_ ;
wire _277_ ;
wire _1595_ ;
wire _1175_ ;
wire _34_ ;
wire _1269_ ;
wire NMI_1 ;
wire _812_ ;
wire _72_ ;
wire _1498_ ;
wire _1078_ ;
wire _621_ ;
wire _201_ ;
wire _850_ ;
wire _430_ ;
wire _906_ ;
wire _715_ ;
wire _1613_ ;
wire _944_ ;
wire _524_ ;
wire _104_ ;
wire adc_bcd ;
wire _1422_ ;
wire _1002_ ;
wire _753_ ;
wire _333_ ;
wire _809_ ;
wire _69_ ;
wire _1651_ ;
wire _1231_ ;
wire _982_ ;
wire _562_ ;
wire _142_ ;
wire _618_ ;
wire _1460_ ;
wire _1040_ ;
wire _791_ ;
wire _371_ ;
wire _1516_ ;
wire _847_ ;
wire _427_ ;
wire _180_ ;
wire _1325_ ;
wire _656_ ;
wire _236_ ;
wire _1554_ ;
wire _1134_ ;
wire _885_ ;
wire _465_ ;
wire _1363_ ;
wire _694_ ;
wire _274_ ;
wire _1419_ ;
wire _1592_ ;
wire _1172_ ;
wire _1648_ ;
wire _1228_ ;
wire _979_ ;
wire _559_ ;
wire _139_ ;
wire _31_ ;
wire _1457_ ;
wire _1037_ ;
wire _788_ ;
wire _368_ ;
wire _1266_ ;
wire _597_ ;
wire _177_ ;
wire _1495_ ;
wire _1075_ ;
wire _903_ ;
wire [7:0] \AXYS[2]  ;
wire _1589_ ;
wire _1169_ ;
wire _712_ ;
wire [7:0] ABH ;
wire [7:0] ABL ;
wire _1398_ ;
wire _28_ ;
wire _1610_ ;
wire _941_ ;
wire _521_ ;
wire _101_ ;
wire _750_ ;
wire _330_ ;
wire NMI_edge ;
wire _806_ ;
wire _66_ ;
wire _615_ ;
wire _1513_ ;
wire _844_ ;
wire _424_ ;
wire _1322_ ;
wire _653_ ;
wire _233_ ;
wire load_reg ;
wire _709_ ;
wire _1551_ ;
wire _1131_ ;
wire _882_ ;
wire _462_ ;
wire _1607_ ;
wire _938_ ;
wire _518_ ;
wire _1360_ ;
wire _691_ ;
wire _271_ ;
wire _1416_ ;
wire _747_ ;
wire _327_ ;
wire _1645_ ;
wire _1225_ ;
wire _976_ ;
wire _556_ ;
wire _136_ ;
wire \ALU.V  ;
wire _1454_ ;
wire _1034_ ;
wire _785_ ;
wire _365_ ;
wire _1263_ ;
wire _594_ ;
wire _174_ ;
wire _1319_ ;
wire _1492_ ;
wire _1072_ ;
wire inc ;
wire _1548_ ;
wire _1128_ ;
wire _879_ ;
wire _459_ ;
wire _1357_ ;
wire _688_ ;
wire _268_ ;
wire _900_ ;
wire _1586_ ;
wire _1166_ ;
wire _497_ ;
wire _1395_ ;
wire _25_ ;
wire _803_ ;
wire _63_ ;
wire _1489_ ;
wire _1069_ ;
wire _612_ ;
wire _1298_ ;
wire reset ;
wire _1510_ ;
wire _841_ ;
wire _421_ ;
wire _650_ ;
wire _230_ ;
wire _706_ ;
wire _1604_ ;
wire _935_ ;
wire _515_ ;
wire _1413_ ;
wire _744_ ;
wire _324_ ;
wire _1642_ ;
wire _1222_ ;
wire _973_ ;
wire _553_ ;
wire _133_ ;
wire _609_ ;
wire _1451_ ;
wire _1031_ ;
wire _782_ ;
wire _362_ ;
wire _1507_ ;
wire _838_ ;
wire _418_ ;
wire _98_ ;
wire _1260_ ;
wire _591_ ;
wire _171_ ;
wire _1316_ ;
wire _647_ ;
wire _227_ ;
wire _1545_ ;
wire _1125_ ;
wire _876_ ;
wire _456_ ;
wire _1354_ ;
wire _685_ ;
wire _265_ ;
wire _1583_ ;
wire _1163_ ;
wire _494_ ;
wire _1639_ ;
wire _1219_ ;
wire _1392_ ;
wire _22_ ;
wire _1448_ ;
wire _1028_ ;
wire _779_ ;
wire _359_ ;

BUFX2 BUFX2_insert86 (
    .A(_815_),
    .Y(_815__bF$buf0)
);

BUFX2 BUFX2_insert85 (
    .A(_815_),
    .Y(_815__bF$buf1)
);

BUFX2 BUFX2_insert84 (
    .A(_815_),
    .Y(_815__bF$buf2)
);

BUFX2 BUFX2_insert83 (
    .A(_815_),
    .Y(_815__bF$buf3)
);

BUFX2 BUFX2_insert82 (
    .A(_815_),
    .Y(_815__bF$buf4)
);

BUFX2 BUFX2_insert81 (
    .A(_856_),
    .Y(_856__bF$buf0)
);

BUFX2 BUFX2_insert80 (
    .A(_856_),
    .Y(_856__bF$buf1)
);

BUFX2 BUFX2_insert79 (
    .A(_856_),
    .Y(_856__bF$buf2)
);

BUFX2 BUFX2_insert78 (
    .A(_856_),
    .Y(_856__bF$buf3)
);

BUFX2 BUFX2_insert77 (
    .A(_859_),
    .Y(_859__bF$buf0)
);

BUFX2 BUFX2_insert76 (
    .A(_859_),
    .Y(_859__bF$buf1)
);

BUFX2 BUFX2_insert75 (
    .A(_859_),
    .Y(_859__bF$buf2)
);

BUFX2 BUFX2_insert74 (
    .A(_859_),
    .Y(_859__bF$buf3)
);

BUFX2 BUFX2_insert73 (
    .A(_836_),
    .Y(_836__bF$buf0)
);

BUFX2 BUFX2_insert72 (
    .A(_836_),
    .Y(_836__bF$buf1)
);

BUFX2 BUFX2_insert71 (
    .A(_836_),
    .Y(_836__bF$buf2)
);

BUFX2 BUFX2_insert70 (
    .A(_836_),
    .Y(_836__bF$buf3)
);

BUFX2 BUFX2_insert69 (
    .A(_836_),
    .Y(_836__bF$buf4)
);

BUFX2 BUFX2_insert68 (
    .A(_836_),
    .Y(_836__bF$buf5)
);

BUFX2 BUFX2_insert67 (
    .A(_836_),
    .Y(_836__bF$buf6)
);

BUFX2 BUFX2_insert66 (
    .A(_836_),
    .Y(_836__bF$buf7)
);

BUFX2 BUFX2_insert65 (
    .A(_854_),
    .Y(_854__bF$buf0)
);

BUFX2 BUFX2_insert64 (
    .A(_854_),
    .Y(_854__bF$buf1)
);

BUFX2 BUFX2_insert63 (
    .A(_854_),
    .Y(_854__bF$buf2)
);

BUFX2 BUFX2_insert62 (
    .A(_854_),
    .Y(_854__bF$buf3)
);

BUFX2 BUFX2_insert61 (
    .A(_860_),
    .Y(_860__bF$buf0)
);

BUFX2 BUFX2_insert60 (
    .A(_860_),
    .Y(_860__bF$buf1)
);

BUFX2 BUFX2_insert59 (
    .A(_860_),
    .Y(_860__bF$buf2)
);

BUFX2 BUFX2_insert58 (
    .A(_860_),
    .Y(_860__bF$buf3)
);

BUFX2 BUFX2_insert57 (
    .A(_860_),
    .Y(_860__bF$buf4)
);

BUFX2 BUFX2_insert56 (
    .A(_1629_),
    .Y(_1629__bF$buf0)
);

BUFX2 BUFX2_insert55 (
    .A(_1629_),
    .Y(_1629__bF$buf1)
);

BUFX2 BUFX2_insert54 (
    .A(_1629_),
    .Y(_1629__bF$buf2)
);

BUFX2 BUFX2_insert53 (
    .A(_1629_),
    .Y(_1629__bF$buf3)
);

BUFX2 BUFX2_insert52 (
    .A(_1074_),
    .Y(_1074__bF$buf0)
);

BUFX2 BUFX2_insert51 (
    .A(_1074_),
    .Y(_1074__bF$buf1)
);

BUFX2 BUFX2_insert50 (
    .A(_1074_),
    .Y(_1074__bF$buf2)
);

BUFX2 BUFX2_insert49 (
    .A(_1074_),
    .Y(_1074__bF$buf3)
);

CLKBUF1 CLKBUF1_insert48 (
    .A(clk),
    .Y(clk_bF$buf0)
);

CLKBUF1 CLKBUF1_insert47 (
    .A(clk),
    .Y(clk_bF$buf1)
);

CLKBUF1 CLKBUF1_insert46 (
    .A(clk),
    .Y(clk_bF$buf2)
);

CLKBUF1 CLKBUF1_insert45 (
    .A(clk),
    .Y(clk_bF$buf3)
);

CLKBUF1 CLKBUF1_insert44 (
    .A(clk),
    .Y(clk_bF$buf4)
);

CLKBUF1 CLKBUF1_insert43 (
    .A(clk),
    .Y(clk_bF$buf5)
);

CLKBUF1 CLKBUF1_insert42 (
    .A(clk),
    .Y(clk_bF$buf6)
);

CLKBUF1 CLKBUF1_insert41 (
    .A(clk),
    .Y(clk_bF$buf7)
);

CLKBUF1 CLKBUF1_insert40 (
    .A(clk),
    .Y(clk_bF$buf8)
);

CLKBUF1 CLKBUF1_insert39 (
    .A(clk),
    .Y(clk_bF$buf9)
);

CLKBUF1 CLKBUF1_insert38 (
    .A(clk),
    .Y(clk_bF$buf10)
);

BUFX2 BUFX2_insert37 (
    .A(_1_),
    .Y(_1__bF$buf0)
);

BUFX2 BUFX2_insert36 (
    .A(_1_),
    .Y(_1__bF$buf1)
);

BUFX2 BUFX2_insert35 (
    .A(_1_),
    .Y(_1__bF$buf2)
);

BUFX2 BUFX2_insert34 (
    .A(_1_),
    .Y(_1__bF$buf3)
);

BUFX2 BUFX2_insert33 (
    .A(_1_),
    .Y(_1__bF$buf4)
);

BUFX2 BUFX2_insert32 (
    .A(_1_),
    .Y(_1__bF$buf5)
);

BUFX2 BUFX2_insert31 (
    .A(_1_),
    .Y(_1__bF$buf6)
);

BUFX2 BUFX2_insert30 (
    .A(_1_),
    .Y(_1__bF$buf7)
);

BUFX2 BUFX2_insert29 (
    .A(_1_),
    .Y(_1__bF$buf8)
);

BUFX2 BUFX2_insert28 (
    .A(_1_),
    .Y(_1__bF$buf9)
);

BUFX2 BUFX2_insert27 (
    .A(_1_),
    .Y(_1__bF$buf10)
);

BUFX2 BUFX2_insert26 (
    .A(_917_),
    .Y(_917__bF$buf0)
);

BUFX2 BUFX2_insert25 (
    .A(_917_),
    .Y(_917__bF$buf1)
);

BUFX2 BUFX2_insert24 (
    .A(_917_),
    .Y(_917__bF$buf2)
);

BUFX2 BUFX2_insert23 (
    .A(_917_),
    .Y(_917__bF$buf3)
);

BUFX2 BUFX2_insert22 (
    .A(_917_),
    .Y(_917__bF$buf4)
);

BUFX2 BUFX2_insert21 (
    .A(_861_),
    .Y(_861__bF$buf0)
);

BUFX2 BUFX2_insert20 (
    .A(_861_),
    .Y(_861__bF$buf1)
);

BUFX2 BUFX2_insert19 (
    .A(_861_),
    .Y(_861__bF$buf2)
);

BUFX2 BUFX2_insert18 (
    .A(_861_),
    .Y(_861__bF$buf3)
);

BUFX2 BUFX2_insert17 (
    .A(_899_),
    .Y(_899__bF$buf0)
);

BUFX2 BUFX2_insert16 (
    .A(_899_),
    .Y(_899__bF$buf1)
);

BUFX2 BUFX2_insert15 (
    .A(_899_),
    .Y(_899__bF$buf2)
);

BUFX2 BUFX2_insert14 (
    .A(_899_),
    .Y(_899__bF$buf3)
);

BUFX2 BUFX2_insert13 (
    .A(_899_),
    .Y(_899__bF$buf4)
);

BUFX2 BUFX2_insert12 (
    .A(_923_),
    .Y(_923__bF$buf0)
);

BUFX2 BUFX2_insert11 (
    .A(_923_),
    .Y(_923__bF$buf1)
);

BUFX2 BUFX2_insert10 (
    .A(_923_),
    .Y(_923__bF$buf2)
);

BUFX2 BUFX2_insert9 (
    .A(_923_),
    .Y(_923__bF$buf3)
);

BUFX2 BUFX2_insert8 (
    .A(RDY),
    .Y(RDY_bF$buf0)
);

BUFX2 BUFX2_insert7 (
    .A(RDY),
    .Y(RDY_bF$buf1)
);

BUFX2 BUFX2_insert6 (
    .A(RDY),
    .Y(RDY_bF$buf2)
);

BUFX2 BUFX2_insert5 (
    .A(RDY),
    .Y(RDY_bF$buf3)
);

BUFX2 BUFX2_insert4 (
    .A(RDY),
    .Y(RDY_bF$buf4)
);

BUFX2 BUFX2_insert3 (
    .A(RDY),
    .Y(RDY_bF$buf5)
);

BUFX2 BUFX2_insert2 (
    .A(RDY),
    .Y(RDY_bF$buf6)
);

BUFX2 BUFX2_insert1 (
    .A(RDY),
    .Y(RDY_bF$buf7)
);

BUFX2 BUFX2_insert0 (
    .A(RDY),
    .Y(RDY_bF$buf8)
);

INVX1 _1668_ (
    .A(DIHOLD[0]),
    .Y(_832_)
);

NAND2X1 _1669_ (
    .A(RDY_bF$buf8),
    .B(DI[0]),
    .Y(_833_)
);

OAI21X1 _1670_ (
    .A(RDY_bF$buf7),
    .B(_832_),
    .C(_833_),
    .Y(DIMUX[0])
);

INVX1 _1671_ (
    .A(DIHOLD[1]),
    .Y(_834_)
);

NAND2X1 _1672_ (
    .A(RDY_bF$buf6),
    .B(DI[1]),
    .Y(_835_)
);

OAI21X1 _1673_ (
    .A(RDY_bF$buf5),
    .B(_834_),
    .C(_835_),
    .Y(DIMUX[1])
);

INVX8 _1674_ (
    .A(RDY_bF$buf4),
    .Y(_836_)
);

OR2X2 _1675_ (
    .A(RDY_bF$buf3),
    .B(DIHOLD[2]),
    .Y(_837_)
);

OAI21X1 _1676_ (
    .A(_836__bF$buf7),
    .B(DI[2]),
    .C(_837_),
    .Y(_838_)
);

INVX1 _1677_ (
    .A(_838_),
    .Y(DIMUX[2])
);

INVX1 _1678_ (
    .A(DIHOLD[3]),
    .Y(_839_)
);

NAND2X1 _1679_ (
    .A(RDY_bF$buf2),
    .B(DI[3]),
    .Y(_840_)
);

OAI21X1 _1680_ (
    .A(RDY_bF$buf1),
    .B(_839_),
    .C(_840_),
    .Y(DIMUX[3])
);

INVX1 _1681_ (
    .A(DIHOLD[4]),
    .Y(_841_)
);

NAND2X1 _1682_ (
    .A(RDY_bF$buf0),
    .B(DI[4]),
    .Y(_842_)
);

OAI21X1 _1683_ (
    .A(RDY_bF$buf8),
    .B(_841_),
    .C(_842_),
    .Y(DIMUX[4])
);

OR2X2 _1684_ (
    .A(RDY_bF$buf7),
    .B(DIHOLD[5]),
    .Y(_843_)
);

OAI21X1 _1685_ (
    .A(_836__bF$buf6),
    .B(DI[5]),
    .C(_843_),
    .Y(_844_)
);

INVX1 _1686_ (
    .A(_844_),
    .Y(DIMUX[5])
);

OR2X2 _1687_ (
    .A(RDY_bF$buf6),
    .B(DIHOLD[6]),
    .Y(_845_)
);

OAI21X1 _1688_ (
    .A(_836__bF$buf5),
    .B(DI[6]),
    .C(_845_),
    .Y(_846_)
);

INVX1 _1689_ (
    .A(_846_),
    .Y(DIMUX[6])
);

MUX2X1 _1690_ (
    .A(DI[7]),
    .B(DIHOLD[7]),
    .S(RDY_bF$buf5),
    .Y(_847_)
);

INVX1 _1691_ (
    .A(_847_),
    .Y(DIMUX[7])
);

INVX1 _1692_ (
    .A(state[1]),
    .Y(_848_)
);

NAND2X1 _1693_ (
    .A(state[0]),
    .B(_848_),
    .Y(_849_)
);

INVX1 _1694_ (
    .A(state[3]),
    .Y(_850_)
);

NAND2X1 _1695_ (
    .A(state[2]),
    .B(_850_),
    .Y(_851_)
);

NOR2X1 _1696_ (
    .A(_849_),
    .B(_851_),
    .Y(_852_)
);

INVX2 _1697_ (
    .A(state[5]),
    .Y(_853_)
);

NOR2X1 _1698_ (
    .A(state[4]),
    .B(_853_),
    .Y(_854_)
);

NAND2X1 _1699_ (
    .A(_854__bF$buf3),
    .B(_852_),
    .Y(_855_)
);

NOR2X1 _1700_ (
    .A(state[5]),
    .B(state[4]),
    .Y(_856_)
);

AND2X2 _1701_ (
    .A(state[3]),
    .B(state[2]),
    .Y(_857_)
);

NOR2X1 _1702_ (
    .A(state[1]),
    .B(state[0]),
    .Y(_858_)
);

NAND3X1 _1703_ (
    .A(_856__bF$buf3),
    .B(_857_),
    .C(_858_),
    .Y(_859_)
);

NOR2X1 _1704_ (
    .A(_836__bF$buf4),
    .B(_859__bF$buf3),
    .Y(_860_)
);

INVX4 _1705_ (
    .A(_860__bF$buf4),
    .Y(_861_)
);

NOR2X1 _1706_ (
    .A(IRHOLD_valid),
    .B(DIMUX[3]),
    .Y(_862_)
);

INVX1 _1707_ (
    .A(IRHOLD_valid),
    .Y(_863_)
);

INVX1 _1708_ (
    .A(I),
    .Y(_864_)
);

INVX1 _1709_ (
    .A(IRQ),
    .Y(_865_)
);

INVX1 _1710_ (
    .A(NMI_edge),
    .Y(_866_)
);

NAND2X1 _1711_ (
    .A(_865_),
    .B(_866_),
    .Y(_867_)
);

OAI21X1 _1712_ (
    .A(_864_),
    .B(NMI_edge),
    .C(_867_),
    .Y(_868_)
);

OAI21X1 _1713_ (
    .A(_863_),
    .B(IRHOLD[3]),
    .C(_868_),
    .Y(_869_)
);

NAND2X1 _1714_ (
    .A(IRHOLD_valid),
    .B(IRHOLD[2]),
    .Y(_870_)
);

OAI21X1 _1715_ (
    .A(IRHOLD_valid),
    .B(_838_),
    .C(_870_),
    .Y(_871_)
);

NAND2X1 _1716_ (
    .A(_868_),
    .B(_871_),
    .Y(_872_)
);

OAI21X1 _1717_ (
    .A(_862_),
    .B(_869_),
    .C(_872_),
    .Y(_873_)
);

OAI21X1 _1718_ (
    .A(I),
    .B(_865_),
    .C(_866_),
    .Y(_874_)
);

INVX1 _1719_ (
    .A(IRHOLD[1]),
    .Y(_875_)
);

AOI21X1 _1720_ (
    .A(IRHOLD_valid),
    .B(_875_),
    .C(_874_),
    .Y(_876_)
);

OAI21X1 _1721_ (
    .A(IRHOLD_valid),
    .B(DIMUX[1]),
    .C(_876_),
    .Y(_877_)
);

MUX2X1 _1722_ (
    .A(DIMUX[0]),
    .B(IRHOLD[0]),
    .S(_863_),
    .Y(_878_)
);

OAI21X1 _1723_ (
    .A(_874_),
    .B(_878_),
    .C(_877_),
    .Y(_879_)
);

NOR2X1 _1724_ (
    .A(_879_),
    .B(_873_),
    .Y(_880_)
);

INVX1 _1725_ (
    .A(IRHOLD[4]),
    .Y(_881_)
);

AOI21X1 _1726_ (
    .A(IRHOLD_valid),
    .B(_881_),
    .C(_874_),
    .Y(_882_)
);

OAI21X1 _1727_ (
    .A(IRHOLD_valid),
    .B(DIMUX[4]),
    .C(_882_),
    .Y(_883_)
);

NAND2X1 _1728_ (
    .A(IRHOLD_valid),
    .B(IRHOLD[5]),
    .Y(_884_)
);

OAI21X1 _1729_ (
    .A(IRHOLD_valid),
    .B(_844_),
    .C(_884_),
    .Y(_885_)
);

NAND2X1 _1730_ (
    .A(_868_),
    .B(_885_),
    .Y(_886_)
);

NAND2X1 _1731_ (
    .A(_883_),
    .B(_886_),
    .Y(_887_)
);

NAND2X1 _1732_ (
    .A(IRHOLD[7]),
    .B(IRHOLD_valid),
    .Y(_888_)
);

OAI21X1 _1733_ (
    .A(IRHOLD_valid),
    .B(_847_),
    .C(_888_),
    .Y(_889_)
);

NAND2X1 _1734_ (
    .A(_868_),
    .B(_889_),
    .Y(_890_)
);

NAND2X1 _1735_ (
    .A(IRHOLD_valid),
    .B(IRHOLD[6]),
    .Y(_891_)
);

OAI21X1 _1736_ (
    .A(IRHOLD_valid),
    .B(_846_),
    .C(_891_),
    .Y(_892_)
);

AND2X2 _1737_ (
    .A(_892_),
    .B(_868_),
    .Y(_893_)
);

NAND2X1 _1738_ (
    .A(_890_),
    .B(_893_),
    .Y(_894_)
);

NOR2X1 _1739_ (
    .A(_887_),
    .B(_894_),
    .Y(_895_)
);

NAND2X1 _1740_ (
    .A(_880_),
    .B(_895_),
    .Y(_896_)
);

OAI22X1 _1741_ (
    .A(RDY_bF$buf4),
    .B(_855_),
    .C(_861__bF$buf3),
    .D(_896_),
    .Y(_897_)
);

INVX1 _1742_ (
    .A(_897_),
    .Y(_898_)
);

NAND2X1 _1743_ (
    .A(state[4]),
    .B(_853_),
    .Y(_899_)
);

INVX4 _1744_ (
    .A(_899__bF$buf4),
    .Y(_900_)
);

NAND2X1 _1745_ (
    .A(_900_),
    .B(_852_),
    .Y(_901_)
);

NOR2X1 _1746_ (
    .A(\ALU.CO ),
    .B(store),
    .Y(_902_)
);

INVX1 _1747_ (
    .A(state[2]),
    .Y(_903_)
);

NOR2X1 _1748_ (
    .A(state[3]),
    .B(_903_),
    .Y(_904_)
);

NAND2X1 _1749_ (
    .A(_858_),
    .B(_904_),
    .Y(_905_)
);

NOR2X1 _1750_ (
    .A(_899__bF$buf3),
    .B(_905_),
    .Y(_906_)
);

NAND2X1 _1751_ (
    .A(RDY_bF$buf3),
    .B(_906_),
    .Y(_907_)
);

OAI22X1 _1752_ (
    .A(RDY_bF$buf2),
    .B(_901_),
    .C(_902_),
    .D(_907_),
    .Y(_908_)
);

INVX1 _1753_ (
    .A(_908_),
    .Y(_909_)
);

INVX1 _1754_ (
    .A(state[0]),
    .Y(_910_)
);

NOR2X1 _1755_ (
    .A(state[1]),
    .B(_910_),
    .Y(_911_)
);

NOR2X1 _1756_ (
    .A(state[3]),
    .B(state[2]),
    .Y(_912_)
);

NAND2X1 _1757_ (
    .A(_912_),
    .B(_911_),
    .Y(_913_)
);

INVX2 _1758_ (
    .A(state[4]),
    .Y(_914_)
);

NOR2X1 _1759_ (
    .A(_853_),
    .B(_914_),
    .Y(_915_)
);

INVX1 _1760_ (
    .A(_915_),
    .Y(_916_)
);

INVX8 _1761_ (
    .A(_854__bF$buf2),
    .Y(_917_)
);

NAND2X1 _1762_ (
    .A(state[3]),
    .B(state[2]),
    .Y(_918_)
);

NAND2X1 _1763_ (
    .A(state[1]),
    .B(state[0]),
    .Y(_919_)
);

NOR2X1 _1764_ (
    .A(_918_),
    .B(_919_),
    .Y(_920_)
);

INVX1 _1765_ (
    .A(_920_),
    .Y(_921_)
);

NOR2X1 _1766_ (
    .A(_917__bF$buf4),
    .B(_921_),
    .Y(_922_)
);

INVX8 _1767_ (
    .A(_856__bF$buf2),
    .Y(_923_)
);

NAND2X1 _1768_ (
    .A(_848_),
    .B(_910_),
    .Y(_924_)
);

NOR2X1 _1769_ (
    .A(_851_),
    .B(_924_),
    .Y(_925_)
);

NAND2X1 _1770_ (
    .A(_856__bF$buf1),
    .B(_925_),
    .Y(_926_)
);

OAI21X1 _1771_ (
    .A(_923__bF$buf3),
    .B(_913_),
    .C(_926_),
    .Y(_927_)
);

NOR2X1 _1772_ (
    .A(_922_),
    .B(_927_),
    .Y(_928_)
);

OAI21X1 _1773_ (
    .A(_913_),
    .B(_916_),
    .C(_928_),
    .Y(_929_)
);

AOI21X1 _1774_ (
    .A(_929_),
    .B(write_back),
    .C(_836__bF$buf3),
    .Y(_930_)
);

NAND2X1 _1775_ (
    .A(state[1]),
    .B(_910_),
    .Y(_931_)
);

NOR2X1 _1776_ (
    .A(_918_),
    .B(_931_),
    .Y(_932_)
);

INVX2 _1777_ (
    .A(_932_),
    .Y(_933_)
);

NOR2X1 _1778_ (
    .A(_917__bF$buf3),
    .B(_933_),
    .Y(_934_)
);

INVX2 _1779_ (
    .A(_934_),
    .Y(_935_)
);

OAI21X1 _1780_ (
    .A(_899__bF$buf2),
    .B(_913_),
    .C(_935_),
    .Y(_936_)
);

INVX1 _1781_ (
    .A(_852_),
    .Y(_937_)
);

NOR2X1 _1782_ (
    .A(_918_),
    .B(_849_),
    .Y(_938_)
);

OAI21X1 _1783_ (
    .A(_854__bF$buf1),
    .B(_900_),
    .C(_938_),
    .Y(_939_)
);

OAI21X1 _1784_ (
    .A(_899__bF$buf1),
    .B(_937_),
    .C(_939_),
    .Y(_940_)
);

OR2X2 _1785_ (
    .A(_936_),
    .B(_940_),
    .Y(_941_)
);

OAI21X1 _1786_ (
    .A(_929_),
    .B(_941_),
    .C(_930_),
    .Y(_942_)
);

INVX1 _1787_ (
    .A(_902_),
    .Y(_943_)
);

NOR2X1 _1788_ (
    .A(write_back),
    .B(_943_),
    .Y(_944_)
);

INVX1 _1789_ (
    .A(_912_),
    .Y(_945_)
);

NOR2X1 _1790_ (
    .A(_919_),
    .B(_945_),
    .Y(_946_)
);

NAND2X1 _1791_ (
    .A(_856__bF$buf0),
    .B(_946_),
    .Y(_947_)
);

NOR2X1 _1792_ (
    .A(_836__bF$buf2),
    .B(_947_),
    .Y(_948_)
);

NAND2X1 _1793_ (
    .A(_944_),
    .B(_948_),
    .Y(_949_)
);

AND2X2 _1794_ (
    .A(_857_),
    .B(_858_),
    .Y(_950_)
);

NAND2X1 _1795_ (
    .A(_900_),
    .B(_950_),
    .Y(_951_)
);

AOI21X1 _1796_ (
    .A(_938_),
    .B(_900_),
    .C(RDY_bF$buf1),
    .Y(_952_)
);

AOI21X1 _1797_ (
    .A(RDY_bF$buf0),
    .B(_951_),
    .C(_952_),
    .Y(_953_)
);

NAND2X1 _1798_ (
    .A(_857_),
    .B(_911_),
    .Y(_954_)
);

NOR2X1 _1799_ (
    .A(_923__bF$buf2),
    .B(_954_),
    .Y(_955_)
);

AOI21X1 _1800_ (
    .A(_836__bF$buf1),
    .B(_955_),
    .C(_953_),
    .Y(_956_)
);

NAND2X1 _1801_ (
    .A(_858_),
    .B(_857_),
    .Y(_957_)
);

NOR2X1 _1802_ (
    .A(_957_),
    .B(_917__bF$buf2),
    .Y(_958_)
);

OAI21X1 _1803_ (
    .A(_917__bF$buf1),
    .B(_954_),
    .C(_836__bF$buf0),
    .Y(_959_)
);

OAI21X1 _1804_ (
    .A(_836__bF$buf7),
    .B(_958_),
    .C(_959_),
    .Y(_960_)
);

INVX1 _1805_ (
    .A(_960_),
    .Y(_961_)
);

NOR2X1 _1806_ (
    .A(_943_),
    .B(_907_),
    .Y(_962_)
);

NOR2X1 _1807_ (
    .A(_961_),
    .B(_962_),
    .Y(_963_)
);

NAND3X1 _1808_ (
    .A(_949_),
    .B(_956_),
    .C(_963_),
    .Y(_964_)
);

INVX2 _1809_ (
    .A(_883_),
    .Y(_965_)
);

NOR2X1 _1810_ (
    .A(_861__bF$buf2),
    .B(_965_),
    .Y(_966_)
);

NOR2X1 _1811_ (
    .A(_862_),
    .B(_869_),
    .Y(_967_)
);

NAND2X1 _1812_ (
    .A(_872_),
    .B(_967_),
    .Y(_968_)
);

INVX1 _1813_ (
    .A(_968_),
    .Y(_969_)
);

NOR2X1 _1814_ (
    .A(_874_),
    .B(_878_),
    .Y(_970_)
);

NAND2X1 _1815_ (
    .A(_877_),
    .B(_970_),
    .Y(_971_)
);

INVX2 _1816_ (
    .A(_971_),
    .Y(_972_)
);

NAND2X1 _1817_ (
    .A(_972_),
    .B(_969_),
    .Y(_973_)
);

INVX1 _1818_ (
    .A(_890_),
    .Y(_974_)
);

OAI21X1 _1819_ (
    .A(_874_),
    .B(_878_),
    .C(_974_),
    .Y(_975_)
);

OAI21X1 _1820_ (
    .A(_873_),
    .B(_975_),
    .C(_973_),
    .Y(_976_)
);

AOI21X1 _1821_ (
    .A(_966_),
    .B(_976_),
    .C(_964_),
    .Y(_977_)
);

AND2X2 _1822_ (
    .A(_977_),
    .B(_942_),
    .Y(_978_)
);

NAND3X1 _1823_ (
    .A(_898_),
    .B(_909_),
    .C(_978_),
    .Y(_979_)
);

NOR2X1 _1824_ (
    .A(_917__bF$buf0),
    .B(_913_),
    .Y(_980_)
);

NAND2X1 _1825_ (
    .A(_836__bF$buf6),
    .B(_980_),
    .Y(_981_)
);

INVX1 _1826_ (
    .A(_887_),
    .Y(_982_)
);

NOR2X1 _1827_ (
    .A(_879_),
    .B(_968_),
    .Y(_983_)
);

NAND3X1 _1828_ (
    .A(_982_),
    .B(_890_),
    .C(_983_),
    .Y(_984_)
);

OAI21X1 _1829_ (
    .A(_861__bF$buf1),
    .B(_984_),
    .C(_981_),
    .Y(_985_)
);

NAND2X1 _1830_ (
    .A(_856__bF$buf3),
    .B(_852_),
    .Y(_986_)
);

NAND2X1 _1831_ (
    .A(_965_),
    .B(_880_),
    .Y(_987_)
);

OAI22X1 _1832_ (
    .A(RDY_bF$buf8),
    .B(_986_),
    .C(_861__bF$buf0),
    .D(_987_),
    .Y(_988_)
);

NOR2X1 _1833_ (
    .A(state[2]),
    .B(_850_),
    .Y(_989_)
);

NAND2X1 _1834_ (
    .A(_858_),
    .B(_989_),
    .Y(_990_)
);

NOR2X1 _1835_ (
    .A(_899__bF$buf0),
    .B(_990_),
    .Y(_991_)
);

NAND2X1 _1836_ (
    .A(_911_),
    .B(_989_),
    .Y(_992_)
);

OAI21X1 _1837_ (
    .A(_899__bF$buf4),
    .B(_992_),
    .C(_836__bF$buf5),
    .Y(_993_)
);

OAI21X1 _1838_ (
    .A(_836__bF$buf4),
    .B(_991_),
    .C(_993_),
    .Y(_994_)
);

NAND2X1 _1839_ (
    .A(state[3]),
    .B(_903_),
    .Y(_995_)
);

NOR2X1 _1840_ (
    .A(_849_),
    .B(_995_),
    .Y(_996_)
);

NAND2X1 _1841_ (
    .A(_854__bF$buf0),
    .B(_996_),
    .Y(_997_)
);

NOR2X1 _1842_ (
    .A(_917__bF$buf4),
    .B(_990_),
    .Y(_998_)
);

NAND2X1 _1843_ (
    .A(RDY_bF$buf7),
    .B(_998_),
    .Y(_999_)
);

OAI21X1 _1844_ (
    .A(RDY_bF$buf6),
    .B(_997_),
    .C(_999_),
    .Y(_1000_)
);

NOR2X1 _1845_ (
    .A(_923__bF$buf1),
    .B(_990_),
    .Y(_1001_)
);

NAND2X1 _1846_ (
    .A(RDY_bF$buf5),
    .B(_1001_),
    .Y(_1002_)
);

NAND2X1 _1847_ (
    .A(_856__bF$buf2),
    .B(_996_),
    .Y(_1003_)
);

OAI21X1 _1848_ (
    .A(RDY_bF$buf4),
    .B(_1003_),
    .C(_1002_),
    .Y(_1004_)
);

NOR2X1 _1849_ (
    .A(_1004_),
    .B(_1000_),
    .Y(_1005_)
);

NAND2X1 _1850_ (
    .A(_858_),
    .B(_912_),
    .Y(_1006_)
);

INVX2 _1851_ (
    .A(_1006_),
    .Y(_1007_)
);

NAND2X1 _1852_ (
    .A(_915_),
    .B(_1007_),
    .Y(_1008_)
);

NOR2X1 _1853_ (
    .A(_849_),
    .B(_945_),
    .Y(_1009_)
);

AOI21X1 _1854_ (
    .A(_1009_),
    .B(_915_),
    .C(RDY_bF$buf3),
    .Y(_1010_)
);

AOI21X1 _1855_ (
    .A(RDY_bF$buf2),
    .B(_1008_),
    .C(_1010_),
    .Y(_1011_)
);

OAI21X1 _1856_ (
    .A(_899__bF$buf3),
    .B(_1006_),
    .C(RDY_bF$buf1),
    .Y(_1012_)
);

OAI21X1 _1857_ (
    .A(_899__bF$buf2),
    .B(_913_),
    .C(_836__bF$buf3),
    .Y(_1013_)
);

AOI21X1 _1858_ (
    .A(_1012_),
    .B(_1013_),
    .C(_1011_),
    .Y(_1014_)
);

NOR2X1 _1859_ (
    .A(_923__bF$buf0),
    .B(_913_),
    .Y(_1015_)
);

OAI21X1 _1860_ (
    .A(_923__bF$buf3),
    .B(_1006_),
    .C(RDY_bF$buf0),
    .Y(_1016_)
);

OAI21X1 _1861_ (
    .A(RDY_bF$buf8),
    .B(_1015_),
    .C(_1016_),
    .Y(_1017_)
);

AND2X2 _1862_ (
    .A(_1014_),
    .B(_1017_),
    .Y(_1018_)
);

NAND3X1 _1863_ (
    .A(_994_),
    .B(_1005_),
    .C(_1018_),
    .Y(_1019_)
);

NOR3X1 _1864_ (
    .A(_988_),
    .B(_985_),
    .C(_1019_),
    .Y(_1020_)
);

NOR2X1 _1865_ (
    .A(_872_),
    .B(_967_),
    .Y(_1021_)
);

AOI22X1 _1866_ (
    .A(_836__bF$buf2),
    .B(_922_),
    .C(_966_),
    .D(_1021_),
    .Y(_1022_)
);

NAND2X1 _1867_ (
    .A(_856__bF$buf1),
    .B(_920_),
    .Y(_1023_)
);

INVX1 _1868_ (
    .A(_1023_),
    .Y(_1024_)
);

OAI21X1 _1869_ (
    .A(_923__bF$buf2),
    .B(_933_),
    .C(RDY_bF$buf7),
    .Y(_1025_)
);

OAI21X1 _1870_ (
    .A(RDY_bF$buf6),
    .B(_1024_),
    .C(_1025_),
    .Y(_1026_)
);

AND2X2 _1871_ (
    .A(_1022_),
    .B(_1026_),
    .Y(_1027_)
);

NOR2X1 _1872_ (
    .A(_851_),
    .B(_931_),
    .Y(_1028_)
);

INVX2 _1873_ (
    .A(_1028_),
    .Y(_1029_)
);

OAI21X1 _1874_ (
    .A(_899__bF$buf1),
    .B(_1029_),
    .C(RDY_bF$buf5),
    .Y(_1030_)
);

NOR3X1 _1875_ (
    .A(_919_),
    .B(_851_),
    .C(_899__bF$buf0),
    .Y(_1031_)
);

OAI21X1 _1876_ (
    .A(RDY_bF$buf4),
    .B(_1031_),
    .C(_1030_),
    .Y(_1032_)
);

NOR2X1 _1877_ (
    .A(_917__bF$buf3),
    .B(_1029_),
    .Y(_1033_)
);

INVX1 _1878_ (
    .A(_919_),
    .Y(_1034_)
);

NAND2X1 _1879_ (
    .A(_1034_),
    .B(_904_),
    .Y(_1035_)
);

OAI21X1 _1880_ (
    .A(_917__bF$buf2),
    .B(_1035_),
    .C(_836__bF$buf1),
    .Y(_1036_)
);

OAI21X1 _1881_ (
    .A(_836__bF$buf0),
    .B(_1033_),
    .C(_1036_),
    .Y(_1037_)
);

NOR3X1 _1882_ (
    .A(_919_),
    .B(_851_),
    .C(_923__bF$buf1),
    .Y(_1038_)
);

NOR3X1 _1883_ (
    .A(_851_),
    .B(_931_),
    .C(_923__bF$buf0),
    .Y(_1039_)
);

XOR2X1 _1884_ (
    .A(\ALU.CO ),
    .B(backwards),
    .Y(_1040_)
);

AND2X2 _1885_ (
    .A(_1040_),
    .B(RDY_bF$buf3),
    .Y(_1041_)
);

AOI22X1 _1886_ (
    .A(_836__bF$buf7),
    .B(_1038_),
    .C(_1041_),
    .D(_1039_),
    .Y(_1042_)
);

AND2X2 _1887_ (
    .A(_1037_),
    .B(_1042_),
    .Y(_1043_)
);

NAND3X1 _1888_ (
    .A(_1032_),
    .B(_1043_),
    .C(_1027_),
    .Y(_1044_)
);

NAND2X1 _1889_ (
    .A(_900_),
    .B(_946_),
    .Y(_1045_)
);

INVX1 _1890_ (
    .A(_931_),
    .Y(_1046_)
);

NAND2X1 _1891_ (
    .A(_912_),
    .B(_1046_),
    .Y(_1047_)
);

NOR2X1 _1892_ (
    .A(_899__bF$buf4),
    .B(_1047_),
    .Y(_1048_)
);

NAND2X1 _1893_ (
    .A(RDY_bF$buf2),
    .B(_1048_),
    .Y(_1049_)
);

OAI21X1 _1894_ (
    .A(RDY_bF$buf1),
    .B(_1045_),
    .C(_1049_),
    .Y(_1050_)
);

INVX2 _1895_ (
    .A(_1047_),
    .Y(_1051_)
);

NAND2X1 _1896_ (
    .A(_856__bF$buf0),
    .B(_1051_),
    .Y(_1052_)
);

INVX1 _1897_ (
    .A(_947_),
    .Y(_1053_)
);

NAND2X1 _1898_ (
    .A(_836__bF$buf6),
    .B(_1053_),
    .Y(_1054_)
);

OAI21X1 _1899_ (
    .A(_836__bF$buf5),
    .B(_1052_),
    .C(_1054_),
    .Y(_1055_)
);

NOR2X1 _1900_ (
    .A(_1050_),
    .B(_1055_),
    .Y(_1056_)
);

NAND2X1 _1901_ (
    .A(_900_),
    .B(_932_),
    .Y(_1057_)
);

INVX1 _1902_ (
    .A(_1057_),
    .Y(_1058_)
);

OAI21X1 _1903_ (
    .A(_899__bF$buf3),
    .B(_921_),
    .C(_836__bF$buf4),
    .Y(_1059_)
);

OAI21X1 _1904_ (
    .A(_836__bF$buf3),
    .B(_1058_),
    .C(_1059_),
    .Y(_1060_)
);

NAND2X1 _1905_ (
    .A(_1060_),
    .B(_1056_),
    .Y(_1061_)
);

INVX1 _1906_ (
    .A(_946_),
    .Y(_1062_)
);

NOR2X1 _1907_ (
    .A(_917__bF$buf1),
    .B(_1062_),
    .Y(_1063_)
);

INVX1 _1908_ (
    .A(write_back),
    .Y(_1064_)
);

NOR2X1 _1909_ (
    .A(_1064_),
    .B(_836__bF$buf2),
    .Y(_1065_)
);

AOI22X1 _1910_ (
    .A(_836__bF$buf1),
    .B(_1063_),
    .C(_929_),
    .D(_1065_),
    .Y(_1066_)
);

NOR2X1 _1911_ (
    .A(_931_),
    .B(_995_),
    .Y(_1067_)
);

NAND2X1 _1912_ (
    .A(_854__bF$buf3),
    .B(_1067_),
    .Y(_1068_)
);

NOR2X1 _1913_ (
    .A(_919_),
    .B(_995_),
    .Y(_1069_)
);

NAND2X1 _1914_ (
    .A(_854__bF$buf2),
    .B(_1069_),
    .Y(_1070_)
);

INVX1 _1915_ (
    .A(_1070_),
    .Y(_1071_)
);

NAND2X1 _1916_ (
    .A(_836__bF$buf0),
    .B(_1071_),
    .Y(_1072_)
);

OAI21X1 _1917_ (
    .A(_836__bF$buf7),
    .B(_1068_),
    .C(_1072_),
    .Y(_1073_)
);

NAND2X1 _1918_ (
    .A(_856__bF$buf3),
    .B(_1067_),
    .Y(_1074_)
);

NAND2X1 _1919_ (
    .A(_856__bF$buf2),
    .B(_1069_),
    .Y(_1075_)
);

INVX1 _1920_ (
    .A(_1075_),
    .Y(_1076_)
);

NAND2X1 _1921_ (
    .A(_836__bF$buf6),
    .B(_1076_),
    .Y(_1077_)
);

OAI21X1 _1922_ (
    .A(_836__bF$buf5),
    .B(_1074__bF$buf3),
    .C(_1077_),
    .Y(_1078_)
);

NOR2X1 _1923_ (
    .A(_1073_),
    .B(_1078_),
    .Y(_1079_)
);

NAND2X1 _1924_ (
    .A(_900_),
    .B(_1067_),
    .Y(_1080_)
);

INVX1 _1925_ (
    .A(_1080_),
    .Y(_1081_)
);

NAND2X1 _1926_ (
    .A(_1034_),
    .B(_989_),
    .Y(_1082_)
);

OAI21X1 _1927_ (
    .A(_899__bF$buf2),
    .B(_1082_),
    .C(_836__bF$buf4),
    .Y(_1083_)
);

OAI21X1 _1928_ (
    .A(_836__bF$buf3),
    .B(_1081_),
    .C(_1083_),
    .Y(_1084_)
);

NAND3X1 _1929_ (
    .A(_1079_),
    .B(_1084_),
    .C(_1066_),
    .Y(_1085_)
);

NOR3X1 _1930_ (
    .A(_1061_),
    .B(_1085_),
    .C(_1044_),
    .Y(_1086_)
);

NAND2X1 _1931_ (
    .A(_1020_),
    .B(_1086_),
    .Y(_1087_)
);

NOR2X1 _1932_ (
    .A(_979_),
    .B(_1087_),
    .Y(_1088_)
);

INVX1 _1933_ (
    .A(_1088_),
    .Y(_1463_[0])
);

NAND2X1 _1934_ (
    .A(_836__bF$buf2),
    .B(_1081_),
    .Y(_1089_)
);

INVX1 _1935_ (
    .A(_880_),
    .Y(_1090_)
);

NAND2X1 _1936_ (
    .A(_868_),
    .B(_892_),
    .Y(_1091_)
);

NAND2X1 _1937_ (
    .A(_890_),
    .B(_883_),
    .Y(_1092_)
);

NOR2X1 _1938_ (
    .A(_886_),
    .B(_1092_),
    .Y(_1093_)
);

NAND2X1 _1939_ (
    .A(_1091_),
    .B(_1093_),
    .Y(_1094_)
);

NOR2X1 _1940_ (
    .A(_1094_),
    .B(_1090_),
    .Y(_1095_)
);

NAND2X1 _1941_ (
    .A(_860__bF$buf3),
    .B(_1095_),
    .Y(_1096_)
);

INVX1 _1942_ (
    .A(_1068_),
    .Y(_1097_)
);

NOR2X1 _1943_ (
    .A(_1091_),
    .B(_974_),
    .Y(_1098_)
);

NOR2X1 _1944_ (
    .A(_886_),
    .B(_965_),
    .Y(_1099_)
);

NAND2X1 _1945_ (
    .A(_1098_),
    .B(_1099_),
    .Y(_1100_)
);

NOR2X1 _1946_ (
    .A(_1100_),
    .B(_1090_),
    .Y(_1101_)
);

AOI22X1 _1947_ (
    .A(_836__bF$buf1),
    .B(_1097_),
    .C(_1101_),
    .D(_860__bF$buf2),
    .Y(_1102_)
);

NAND3X1 _1948_ (
    .A(_1089_),
    .B(_1096_),
    .C(_1102_),
    .Y(_1103_)
);

NAND2X1 _1949_ (
    .A(_836__bF$buf0),
    .B(_1058_),
    .Y(_1104_)
);

NAND3X1 _1950_ (
    .A(_860__bF$buf1),
    .B(_1093_),
    .C(_983_),
    .Y(_1105_)
);

NAND2X1 _1951_ (
    .A(_914_),
    .B(_932_),
    .Y(_1106_)
);

NAND2X1 _1952_ (
    .A(RDY_bF$buf0),
    .B(_1063_),
    .Y(_1107_)
);

OAI21X1 _1953_ (
    .A(RDY_bF$buf8),
    .B(_1106_),
    .C(_1107_),
    .Y(_1108_)
);

INVX1 _1954_ (
    .A(_873_),
    .Y(_1109_)
);

NAND2X1 _1955_ (
    .A(_972_),
    .B(_1109_),
    .Y(_1110_)
);

INVX1 _1956_ (
    .A(_1110_),
    .Y(_1111_)
);

AOI21X1 _1957_ (
    .A(_1111_),
    .B(_966_),
    .C(_1108_),
    .Y(_1112_)
);

NAND3X1 _1958_ (
    .A(_1104_),
    .B(_1105_),
    .C(_1112_),
    .Y(_1113_)
);

INVX1 _1959_ (
    .A(_941_),
    .Y(_1114_)
);

NOR2X1 _1960_ (
    .A(_836__bF$buf7),
    .B(_929_),
    .Y(_1115_)
);

OAI21X1 _1961_ (
    .A(_899__bF$buf1),
    .B(_992_),
    .C(_1075_),
    .Y(_1116_)
);

NAND3X1 _1962_ (
    .A(_1115_),
    .B(_1116_),
    .C(_1114_),
    .Y(_1117_)
);

NOR2X1 _1963_ (
    .A(_899__bF$buf0),
    .B(_1029_),
    .Y(_1118_)
);

INVX2 _1964_ (
    .A(_872_),
    .Y(_1119_)
);

NAND2X1 _1965_ (
    .A(_967_),
    .B(_1119_),
    .Y(_1120_)
);

NOR2X1 _1966_ (
    .A(_879_),
    .B(_1120_),
    .Y(_1121_)
);

AND2X2 _1967_ (
    .A(_1121_),
    .B(_895_),
    .Y(_1122_)
);

AOI22X1 _1968_ (
    .A(_836__bF$buf6),
    .B(_1118_),
    .C(_1122_),
    .D(_860__bF$buf0),
    .Y(_1123_)
);

OAI21X1 _1969_ (
    .A(_917__bF$buf0),
    .B(_937_),
    .C(RDY_bF$buf7),
    .Y(_1124_)
);

OAI21X1 _1970_ (
    .A(state[4]),
    .B(_1029_),
    .C(_836__bF$buf5),
    .Y(_1125_)
);

AND2X2 _1971_ (
    .A(cond_code[2]),
    .B(Z),
    .Y(_1126_)
);

INVX1 _1972_ (
    .A(V),
    .Y(_1127_)
);

NOR2X1 _1973_ (
    .A(cond_code[2]),
    .B(_1127_),
    .Y(_1128_)
);

OAI21X1 _1974_ (
    .A(_1126_),
    .B(_1128_),
    .C(cond_code[1]),
    .Y(_1129_)
);

MUX2X1 _1975_ (
    .A(C),
    .B(N),
    .S(cond_code[2]),
    .Y(_1130_)
);

OAI21X1 _1976_ (
    .A(cond_code[1]),
    .B(_1130_),
    .C(_1129_),
    .Y(_1131_)
);

XOR2X1 _1977_ (
    .A(_1131_),
    .B(cond_code[0]),
    .Y(_1132_)
);

NOR2X1 _1978_ (
    .A(_836__bF$buf4),
    .B(_986_),
    .Y(_1133_)
);

INVX1 _1979_ (
    .A(_1133_),
    .Y(_1134_)
);

NOR2X1 _1980_ (
    .A(_1134_),
    .B(_1132_),
    .Y(_1135_)
);

AOI21X1 _1981_ (
    .A(_1124_),
    .B(_1125_),
    .C(_1135_),
    .Y(_1136_)
);

NAND3X1 _1982_ (
    .A(_1136_),
    .B(_1117_),
    .C(_1123_),
    .Y(_1137_)
);

NOR3X1 _1983_ (
    .A(_1113_),
    .B(_1103_),
    .C(_1137_),
    .Y(_1138_)
);

NOR2X1 _1984_ (
    .A(_883_),
    .B(_1110_),
    .Y(_1139_)
);

AOI22X1 _1985_ (
    .A(_836__bF$buf3),
    .B(_1048_),
    .C(_1139_),
    .D(_860__bF$buf4),
    .Y(_1140_)
);

OAI21X1 _1986_ (
    .A(_968_),
    .B(_971_),
    .C(_1120_),
    .Y(_1141_)
);

NAND2X1 _1987_ (
    .A(_860__bF$buf3),
    .B(_965_),
    .Y(_1142_)
);

INVX1 _1988_ (
    .A(_1142_),
    .Y(_1143_)
);

INVX1 _1989_ (
    .A(_1074__bF$buf2),
    .Y(_1144_)
);

OAI21X1 _1990_ (
    .A(_923__bF$buf3),
    .B(_992_),
    .C(RDY_bF$buf6),
    .Y(_1145_)
);

OAI21X1 _1991_ (
    .A(RDY_bF$buf5),
    .B(_1144_),
    .C(_1145_),
    .Y(_1146_)
);

OAI21X1 _1992_ (
    .A(_917__bF$buf4),
    .B(_1047_),
    .C(_836__bF$buf2),
    .Y(_1147_)
);

OAI21X1 _1993_ (
    .A(_836__bF$buf1),
    .B(_980_),
    .C(_1147_),
    .Y(_1148_)
);

NAND3X1 _1994_ (
    .A(_856__bF$buf1),
    .B(_1051_),
    .C(_1145_),
    .Y(_1149_)
);

NAND3X1 _1995_ (
    .A(_1148_),
    .B(_1149_),
    .C(_1146_),
    .Y(_1150_)
);

AOI21X1 _1996_ (
    .A(_1141_),
    .B(_1143_),
    .C(_1150_),
    .Y(_1151_)
);

AND2X2 _1997_ (
    .A(_1140_),
    .B(_1151_),
    .Y(_1152_)
);

NAND3X1 _1998_ (
    .A(_1086_),
    .B(_1152_),
    .C(_1138_),
    .Y(_1463_[1])
);

INVX1 _1999_ (
    .A(_979_),
    .Y(_1153_)
);

NOR2X1 _2000_ (
    .A(_1113_),
    .B(_1137_),
    .Y(_1154_)
);

AND2X2 _2001_ (
    .A(_1114_),
    .B(_1115_),
    .Y(_1155_)
);

OAI21X1 _2002_ (
    .A(_925_),
    .B(_1007_),
    .C(_854__bF$buf1),
    .Y(_1156_)
);

NOR2X1 _2003_ (
    .A(_919_),
    .B(_851_),
    .Y(_1157_)
);

AOI21X1 _2004_ (
    .A(_853_),
    .B(_1157_),
    .C(_955_),
    .Y(_1158_)
);

OAI21X1 _2005_ (
    .A(_996_),
    .B(_1051_),
    .C(_854__bF$buf0),
    .Y(_1159_)
);

NAND3X1 _2006_ (
    .A(_1156_),
    .B(_1158_),
    .C(_1159_),
    .Y(_1160_)
);

NAND2X1 _2007_ (
    .A(_1133_),
    .B(_1132_),
    .Y(_1161_)
);

NAND3X1 _2008_ (
    .A(_856__bF$buf0),
    .B(_904_),
    .C(_1046_),
    .Y(_1162_)
);

NOR2X1 _2009_ (
    .A(_1040_),
    .B(_1162_),
    .Y(_1163_)
);

OAI21X1 _2010_ (
    .A(RDY_bF$buf4),
    .B(_958_),
    .C(_1163_),
    .Y(_1164_)
);

INVX1 _2011_ (
    .A(_951_),
    .Y(_1165_)
);

OAI21X1 _2012_ (
    .A(_899__bF$buf4),
    .B(_1082_),
    .C(RDY_bF$buf3),
    .Y(_1166_)
);

OAI21X1 _2013_ (
    .A(RDY_bF$buf2),
    .B(_1165_),
    .C(_1166_),
    .Y(_1167_)
);

INVX1 _2014_ (
    .A(_1167_),
    .Y(_1168_)
);

OAI21X1 _2015_ (
    .A(_917__bF$buf3),
    .B(_1082_),
    .C(RDY_bF$buf1),
    .Y(_1169_)
);

OAI21X1 _2016_ (
    .A(RDY_bF$buf0),
    .B(_958_),
    .C(_1169_),
    .Y(_1170_)
);

OAI21X1 _2017_ (
    .A(RDY_bF$buf8),
    .B(_859__bF$buf2),
    .C(_1170_),
    .Y(_1171_)
);

NOR2X1 _2018_ (
    .A(_1171_),
    .B(_1168_),
    .Y(_1172_)
);

NAND3X1 _2019_ (
    .A(_1161_),
    .B(_1164_),
    .C(_1172_),
    .Y(_1173_)
);

AOI21X1 _2020_ (
    .A(_1155_),
    .B(_1160_),
    .C(_1173_),
    .Y(_1174_)
);

NAND2X1 _2021_ (
    .A(_883_),
    .B(_976_),
    .Y(_1175_)
);

NAND2X1 _2022_ (
    .A(_965_),
    .B(_1141_),
    .Y(_1176_)
);

INVX1 _2023_ (
    .A(_877_),
    .Y(_1177_)
);

OAI21X1 _2024_ (
    .A(_874_),
    .B(_878_),
    .C(_1177_),
    .Y(_1178_)
);

NOR2X1 _2025_ (
    .A(_968_),
    .B(_1178_),
    .Y(_1179_)
);

AOI21X1 _2026_ (
    .A(_1092_),
    .B(_983_),
    .C(_1179_),
    .Y(_1180_)
);

NAND3X1 _2027_ (
    .A(_1176_),
    .B(_1180_),
    .C(_1175_),
    .Y(_1181_)
);

INVX1 _2028_ (
    .A(_1181_),
    .Y(_1182_)
);

NAND2X1 _2029_ (
    .A(_895_),
    .B(_1121_),
    .Y(_1183_)
);

NOR2X1 _2030_ (
    .A(_861__bF$buf3),
    .B(_1021_),
    .Y(_1184_)
);

NAND3X1 _2031_ (
    .A(_987_),
    .B(_1184_),
    .C(_1183_),
    .Y(_1185_)
);

INVX1 _2032_ (
    .A(_879_),
    .Y(_1186_)
);

OR2X2 _2033_ (
    .A(_869_),
    .B(_862_),
    .Y(_1187_)
);

NOR2X1 _2034_ (
    .A(_872_),
    .B(_1187_),
    .Y(_1188_)
);

NAND2X1 _2035_ (
    .A(_1186_),
    .B(_1188_),
    .Y(_1189_)
);

NAND2X1 _2036_ (
    .A(_890_),
    .B(_1091_),
    .Y(_1190_)
);

NOR2X1 _2037_ (
    .A(_887_),
    .B(_1190_),
    .Y(_1191_)
);

NAND2X1 _2038_ (
    .A(_880_),
    .B(_1191_),
    .Y(_1192_)
);

OAI21X1 _2039_ (
    .A(_1100_),
    .B(_1189_),
    .C(_1192_),
    .Y(_1193_)
);

NOR3X1 _2040_ (
    .A(_1111_),
    .B(_1193_),
    .C(_1185_),
    .Y(_1194_)
);

OAI21X1 _2041_ (
    .A(_965_),
    .B(_890_),
    .C(_1094_),
    .Y(_1195_)
);

NAND2X1 _2042_ (
    .A(_971_),
    .B(_1178_),
    .Y(_1196_)
);

NOR2X1 _2043_ (
    .A(_965_),
    .B(_1120_),
    .Y(_1197_)
);

AOI22X1 _2044_ (
    .A(_1196_),
    .B(_1197_),
    .C(_1195_),
    .D(_1121_),
    .Y(_1198_)
);

AND2X2 _2045_ (
    .A(_896_),
    .B(_984_),
    .Y(_1199_)
);

OAI21X1 _2046_ (
    .A(_880_),
    .B(_983_),
    .C(_1093_),
    .Y(_1200_)
);

NAND3X1 _2047_ (
    .A(_1200_),
    .B(_1198_),
    .C(_1199_),
    .Y(_1201_)
);

INVX1 _2048_ (
    .A(_1201_),
    .Y(_1202_)
);

NAND3X1 _2049_ (
    .A(_1182_),
    .B(_1194_),
    .C(_1202_),
    .Y(_1203_)
);

NOR2X1 _2050_ (
    .A(_917__bF$buf2),
    .B(_905_),
    .Y(_1204_)
);

INVX1 _2051_ (
    .A(_1204_),
    .Y(_1205_)
);

OAI22X1 _2052_ (
    .A(RDY_bF$buf7),
    .B(_1205_),
    .C(_861__bF$buf2),
    .D(_1180_),
    .Y(_1206_)
);

OAI21X1 _2053_ (
    .A(write_back),
    .B(_943_),
    .C(_948_),
    .Y(_1207_)
);

OAI21X1 _2054_ (
    .A(_899__bF$buf3),
    .B(_1062_),
    .C(RDY_bF$buf6),
    .Y(_1208_)
);

OAI21X1 _2055_ (
    .A(RDY_bF$buf5),
    .B(_906_),
    .C(_1208_),
    .Y(_1209_)
);

NOR2X1 _2056_ (
    .A(_923__bF$buf2),
    .B(_905_),
    .Y(_1210_)
);

NAND2X1 _2057_ (
    .A(_836__bF$buf0),
    .B(_1210_),
    .Y(_1211_)
);

NAND3X1 _2058_ (
    .A(_1211_),
    .B(_1209_),
    .C(_1207_),
    .Y(_1212_)
);

NOR2X1 _2059_ (
    .A(_1212_),
    .B(_1206_),
    .Y(_1213_)
);

NAND3X1 _2060_ (
    .A(_1174_),
    .B(_1213_),
    .C(_1203_),
    .Y(_1214_)
);

INVX1 _2061_ (
    .A(_1060_),
    .Y(_1215_)
);

OR2X2 _2062_ (
    .A(_988_),
    .B(_1215_),
    .Y(_1216_)
);

OR2X2 _2063_ (
    .A(_1216_),
    .B(_1044_),
    .Y(_1217_)
);

NOR2X1 _2064_ (
    .A(_1217_),
    .B(_1214_),
    .Y(_1218_)
);

NAND3X1 _2065_ (
    .A(_1153_),
    .B(_1154_),
    .C(_1218_),
    .Y(_1463_[2])
);

NOR2X1 _2066_ (
    .A(_861__bF$buf1),
    .B(_1198_),
    .Y(_1219_)
);

NOR2X1 _2067_ (
    .A(_1100_),
    .B(_1189_),
    .Y(_1220_)
);

AOI22X1 _2068_ (
    .A(_836__bF$buf7),
    .B(_991_),
    .C(_1220_),
    .D(_860__bF$buf2),
    .Y(_1221_)
);

OAI21X1 _2069_ (
    .A(_917__bF$buf1),
    .B(_1035_),
    .C(RDY_bF$buf4),
    .Y(_1222_)
);

OAI21X1 _2070_ (
    .A(RDY_bF$buf3),
    .B(_998_),
    .C(_1222_),
    .Y(_1223_)
);

NAND2X1 _2071_ (
    .A(_1223_),
    .B(_1221_),
    .Y(_1224_)
);

OAI21X1 _2072_ (
    .A(_862_),
    .B(_869_),
    .C(_1119_),
    .Y(_1225_)
);

OAI22X1 _2073_ (
    .A(RDY_bF$buf2),
    .B(_1008_),
    .C(_1142_),
    .D(_1225_),
    .Y(_1226_)
);

NOR2X1 _2074_ (
    .A(_899__bF$buf2),
    .B(_1006_),
    .Y(_1227_)
);

NAND2X1 _2075_ (
    .A(_836__bF$buf6),
    .B(_1227_),
    .Y(_1228_)
);

OAI21X1 _2076_ (
    .A(_836__bF$buf5),
    .B(_1023_),
    .C(_1228_),
    .Y(_1229_)
);

OR2X2 _2077_ (
    .A(_1226_),
    .B(_1229_),
    .Y(_1230_)
);

NAND2X1 _2078_ (
    .A(_856__bF$buf3),
    .B(_1007_),
    .Y(_1231_)
);

NAND2X1 _2079_ (
    .A(_920_),
    .B(_900_),
    .Y(_1232_)
);

OAI21X1 _2080_ (
    .A(_1006_),
    .B(_917__bF$buf0),
    .C(_836__bF$buf4),
    .Y(_1233_)
);

INVX1 _2081_ (
    .A(_1233_),
    .Y(_1234_)
);

AOI22X1 _2082_ (
    .A(RDY_bF$buf1),
    .B(_1232_),
    .C(_1234_),
    .D(_1231_),
    .Y(_1235_)
);

NOR2X1 _2083_ (
    .A(_1235_),
    .B(_1230_),
    .Y(_1236_)
);

NAND3X1 _2084_ (
    .A(_1140_),
    .B(_1151_),
    .C(_1236_),
    .Y(_1237_)
);

NOR3X1 _2085_ (
    .A(_1219_),
    .B(_1224_),
    .C(_1237_),
    .Y(_1238_)
);

NAND3X1 _2086_ (
    .A(_1138_),
    .B(_1238_),
    .C(_1088_),
    .Y(_1239_)
);

NAND2X1 _2087_ (
    .A(_1174_),
    .B(_1203_),
    .Y(_1240_)
);

INVX1 _2088_ (
    .A(_1224_),
    .Y(_1241_)
);

NOR2X1 _2089_ (
    .A(_1113_),
    .B(_1103_),
    .Y(_1242_)
);

NAND2X1 _2090_ (
    .A(_942_),
    .B(_977_),
    .Y(_1243_)
);

NAND2X1 _2091_ (
    .A(_1084_),
    .B(_1079_),
    .Y(_1244_)
);

NOR2X1 _2092_ (
    .A(_1215_),
    .B(_1244_),
    .Y(_1245_)
);

NAND3X1 _2093_ (
    .A(_994_),
    .B(_1146_),
    .C(_1005_),
    .Y(_1246_)
);

INVX1 _2094_ (
    .A(_1246_),
    .Y(_1247_)
);

NAND3X1 _2095_ (
    .A(_1027_),
    .B(_1247_),
    .C(_1245_),
    .Y(_1248_)
);

NOR2X1 _2096_ (
    .A(_1243_),
    .B(_1248_),
    .Y(_1249_)
);

NAND3X1 _2097_ (
    .A(_1241_),
    .B(_1249_),
    .C(_1242_),
    .Y(_1250_)
);

NOR2X1 _2098_ (
    .A(_1240_),
    .B(_1250_),
    .Y(_1251_)
);

OAI21X1 _2099_ (
    .A(_1214_),
    .B(_1239_),
    .C(_1251_),
    .Y(_1463_[3])
);

NAND2X1 _2100_ (
    .A(_1117_),
    .B(_1123_),
    .Y(_1252_)
);

INVX1 _2101_ (
    .A(_1252_),
    .Y(_1253_)
);

OAI21X1 _2102_ (
    .A(RDY_bF$buf0),
    .B(_1057_),
    .C(_1105_),
    .Y(_1254_)
);

NAND2X1 _2103_ (
    .A(_1221_),
    .B(_1140_),
    .Y(_1255_)
);

NOR2X1 _2104_ (
    .A(_1254_),
    .B(_1255_),
    .Y(_1256_)
);

NOR2X1 _2105_ (
    .A(_953_),
    .B(_1050_),
    .Y(_1257_)
);

NAND3X1 _2106_ (
    .A(_1032_),
    .B(_909_),
    .C(_1257_),
    .Y(_1258_)
);

NAND2X1 _2107_ (
    .A(_1060_),
    .B(_1084_),
    .Y(_1259_)
);

NAND3X1 _2108_ (
    .A(_1167_),
    .B(_994_),
    .C(_1209_),
    .Y(_1260_)
);

NOR2X1 _2109_ (
    .A(_1259_),
    .B(_1260_),
    .Y(_1261_)
);

NAND2X1 _2110_ (
    .A(_1014_),
    .B(_1261_),
    .Y(_1262_)
);

NOR2X1 _2111_ (
    .A(_1258_),
    .B(_1262_),
    .Y(_1263_)
);

NAND3X1 _2112_ (
    .A(_1089_),
    .B(_1096_),
    .C(_1263_),
    .Y(_1264_)
);

NOR2X1 _2113_ (
    .A(_1230_),
    .B(_1264_),
    .Y(_1265_)
);

NAND3X1 _2114_ (
    .A(_1253_),
    .B(_1256_),
    .C(_1265_),
    .Y(_1463_[4])
);

AND2X2 _2115_ (
    .A(_898_),
    .B(_1102_),
    .Y(_1266_)
);

INVX1 _2116_ (
    .A(_1232_),
    .Y(_1267_)
);

OAI21X1 _2117_ (
    .A(_836__bF$buf3),
    .B(_1267_),
    .C(_1233_),
    .Y(_1268_)
);

NAND3X1 _2118_ (
    .A(_1170_),
    .B(_1223_),
    .C(_1268_),
    .Y(_1269_)
);

NOR2X1 _2119_ (
    .A(_1269_),
    .B(_1226_),
    .Y(_1270_)
);

NAND2X1 _2120_ (
    .A(_1022_),
    .B(_1270_),
    .Y(_1271_)
);

NOR2X1 _2121_ (
    .A(_985_),
    .B(_1271_),
    .Y(_1272_)
);

INVX1 _2122_ (
    .A(_1037_),
    .Y(_1273_)
);

NOR2X1 _2123_ (
    .A(_1011_),
    .B(_1273_),
    .Y(_1274_)
);

NAND3X1 _2124_ (
    .A(_960_),
    .B(_1148_),
    .C(_1274_),
    .Y(_1275_)
);

OAI21X1 _2125_ (
    .A(RDY_bF$buf8),
    .B(_935_),
    .C(_1107_),
    .Y(_1276_)
);

OAI21X1 _2126_ (
    .A(_917__bF$buf4),
    .B(_1029_),
    .C(_836__bF$buf2),
    .Y(_1277_)
);

AOI21X1 _2127_ (
    .A(_1124_),
    .B(_1277_),
    .C(_1276_),
    .Y(_1278_)
);

NOR2X1 _2128_ (
    .A(_1000_),
    .B(_1073_),
    .Y(_1279_)
);

NAND2X1 _2129_ (
    .A(_1279_),
    .B(_1278_),
    .Y(_1280_)
);

NOR2X1 _2130_ (
    .A(_1275_),
    .B(_1280_),
    .Y(_1281_)
);

NAND2X1 _2131_ (
    .A(_1066_),
    .B(_1281_),
    .Y(_1282_)
);

NOR2X1 _2132_ (
    .A(_1206_),
    .B(_1282_),
    .Y(_1283_)
);

NAND3X1 _2133_ (
    .A(_1266_),
    .B(_1272_),
    .C(_1283_),
    .Y(_1463_[5])
);

OAI21X1 _2134_ (
    .A(_899__bF$buf1),
    .B(_905_),
    .C(_1162_),
    .Y(_1284_)
);

OAI21X1 _2135_ (
    .A(_1284_),
    .B(_1053_),
    .C(\ALU.CO ),
    .Y(_1285_)
);

INVX1 _2136_ (
    .A(_1048_),
    .Y(_1286_)
);

NAND3X1 _2137_ (
    .A(_1070_),
    .B(_1057_),
    .C(_1286_),
    .Y(_1287_)
);

OAI21X1 _2138_ (
    .A(_852_),
    .B(_1067_),
    .C(_854__bF$buf3),
    .Y(_1288_)
);

OAI21X1 _2139_ (
    .A(_917__bF$buf3),
    .B(_1035_),
    .C(_1023_),
    .Y(_1289_)
);

NOR2X1 _2140_ (
    .A(_1289_),
    .B(_1033_),
    .Y(_1290_)
);

NAND2X1 _2141_ (
    .A(_1288_),
    .B(_1290_),
    .Y(_1291_)
);

NOR2X1 _2142_ (
    .A(_1287_),
    .B(_1291_),
    .Y(_1292_)
);

INVX1 _2143_ (
    .A(rotate),
    .Y(_1293_)
);

OAI21X1 _2144_ (
    .A(_925_),
    .B(_946_),
    .C(_854__bF$buf2),
    .Y(_1294_)
);

INVX1 _2145_ (
    .A(shift),
    .Y(_1295_)
);

AOI21X1 _2146_ (
    .A(_1295_),
    .B(inc),
    .C(rotate),
    .Y(_1296_)
);

INVX1 _2147_ (
    .A(compare),
    .Y(_1297_)
);

NAND2X1 _2148_ (
    .A(C),
    .B(_1295_),
    .Y(_1298_)
);

OAI21X1 _2149_ (
    .A(load_only),
    .B(_1298_),
    .C(_1297_),
    .Y(_1299_)
);

OAI21X1 _2150_ (
    .A(rotate),
    .B(_1299_),
    .C(_955_),
    .Y(_1300_)
);

OAI21X1 _2151_ (
    .A(_1294_),
    .B(_1296_),
    .C(_1300_),
    .Y(_1301_)
);

OAI21X1 _2152_ (
    .A(C),
    .B(_1293_),
    .C(_1301_),
    .Y(_1302_)
);

NAND3X1 _2153_ (
    .A(_1285_),
    .B(_1302_),
    .C(_1292_),
    .Y(\ALU.CI )
);

INVX2 _2154_ (
    .A(PC[0]),
    .Y(_1303_)
);

INVX2 _2155_ (
    .A(DIMUX[0]),
    .Y(_1304_)
);

OAI21X1 _2156_ (
    .A(_917__bF$buf2),
    .B(_913_),
    .C(_1057_),
    .Y(_1305_)
);

NOR2X1 _2157_ (
    .A(_1001_),
    .B(_1305_),
    .Y(_1306_)
);

OAI21X1 _2158_ (
    .A(_917__bF$buf1),
    .B(_905_),
    .C(_951_),
    .Y(_1307_)
);

OAI21X1 _2159_ (
    .A(_923__bF$buf1),
    .B(_992_),
    .C(_986_),
    .Y(_1308_)
);

NOR2X1 _2160_ (
    .A(_1307_),
    .B(_1308_),
    .Y(_1309_)
);

INVX1 _2161_ (
    .A(_1015_),
    .Y(_1310_)
);

INVX1 _2162_ (
    .A(_1063_),
    .Y(_1311_)
);

OAI21X1 _2163_ (
    .A(_923__bF$buf0),
    .B(_957_),
    .C(_855_),
    .Y(_1312_)
);

INVX2 _2164_ (
    .A(_1067_),
    .Y(_1313_)
);

OAI22X1 _2165_ (
    .A(state[4]),
    .B(_1029_),
    .C(state[5]),
    .D(_1313_),
    .Y(_1314_)
);

NOR2X1 _2166_ (
    .A(_1312_),
    .B(_1314_),
    .Y(_1315_)
);

NAND3X1 _2167_ (
    .A(_1310_),
    .B(_1311_),
    .C(_1315_),
    .Y(_1316_)
);

NAND2X1 _2168_ (
    .A(_854__bF$buf1),
    .B(_1051_),
    .Y(_1317_)
);

OAI21X1 _2169_ (
    .A(_899__bF$buf0),
    .B(_1082_),
    .C(_1070_),
    .Y(_1318_)
);

NOR2X1 _2170_ (
    .A(_1289_),
    .B(_1318_),
    .Y(_1319_)
);

NAND3X1 _2171_ (
    .A(_1068_),
    .B(_1317_),
    .C(_1319_),
    .Y(_1320_)
);

NOR2X1 _2172_ (
    .A(_1320_),
    .B(_1316_),
    .Y(_1321_)
);

NAND3X1 _2173_ (
    .A(_1306_),
    .B(_1309_),
    .C(_1321_),
    .Y(_1322_)
);

OAI22X1 _2174_ (
    .A(_1303_),
    .B(_986_),
    .C(_1304_),
    .D(_1322_),
    .Y(\ALU.BI [0])
);

INVX2 _2175_ (
    .A(PC[1]),
    .Y(_1323_)
);

INVX2 _2176_ (
    .A(DIMUX[1]),
    .Y(_1324_)
);

OAI22X1 _2177_ (
    .A(_1323_),
    .B(_986_),
    .C(_1324_),
    .D(_1322_),
    .Y(\ALU.BI [1])
);

INVX1 _2178_ (
    .A(PC[2]),
    .Y(_1325_)
);

OAI22X1 _2179_ (
    .A(_1325_),
    .B(_986_),
    .C(_838_),
    .D(_1322_),
    .Y(\ALU.BI [2])
);

INVX2 _2180_ (
    .A(PC[3]),
    .Y(_1326_)
);

INVX2 _2181_ (
    .A(DIMUX[3]),
    .Y(_1327_)
);

OAI22X1 _2182_ (
    .A(_1326_),
    .B(_986_),
    .C(_1327_),
    .D(_1322_),
    .Y(\ALU.BI [3])
);

INVX1 _2183_ (
    .A(PC[4]),
    .Y(_1328_)
);

INVX1 _2184_ (
    .A(DIMUX[4]),
    .Y(_1329_)
);

OAI22X1 _2185_ (
    .A(_1328_),
    .B(_986_),
    .C(_1329_),
    .D(_1322_),
    .Y(\ALU.BI [4])
);

INVX2 _2186_ (
    .A(PC[5]),
    .Y(_1330_)
);

OAI22X1 _2187_ (
    .A(_1330_),
    .B(_986_),
    .C(_844_),
    .D(_1322_),
    .Y(\ALU.BI [5])
);

INVX2 _2188_ (
    .A(PC[6]),
    .Y(_1331_)
);

OAI22X1 _2189_ (
    .A(_1331_),
    .B(_986_),
    .C(_846_),
    .D(_1322_),
    .Y(\ALU.BI [6])
);

INVX1 _2190_ (
    .A(PC[7]),
    .Y(_1332_)
);

OAI22X1 _2191_ (
    .A(_1332_),
    .B(_986_),
    .C(_847_),
    .D(_1322_),
    .Y(\ALU.BI [7])
);

INVX1 _2192_ (
    .A(src_reg[1]),
    .Y(_1333_)
);

OAI21X1 _2193_ (
    .A(_854__bF$buf0),
    .B(_900_),
    .C(_950_),
    .Y(_1334_)
);

INVX1 _2194_ (
    .A(_1334_),
    .Y(_1335_)
);

NAND3X1 _2195_ (
    .A(_1232_),
    .B(_1075_),
    .C(_1080_),
    .Y(_1336_)
);

NOR2X1 _2196_ (
    .A(_1335_),
    .B(_1336_),
    .Y(_1337_)
);

OAI21X1 _2197_ (
    .A(_917__bF$buf0),
    .B(_1047_),
    .C(_1068_),
    .Y(_1338_)
);

NOR2X1 _2198_ (
    .A(_995_),
    .B(_924_),
    .Y(_1339_)
);

NAND2X1 _2199_ (
    .A(_914_),
    .B(_1339_),
    .Y(_1340_)
);

NAND3X1 _2200_ (
    .A(_1057_),
    .B(_855_),
    .C(_1340_),
    .Y(_1341_)
);

NOR2X1 _2201_ (
    .A(_1338_),
    .B(_1341_),
    .Y(_1342_)
);

INVX4 _2202_ (
    .A(_859__bF$buf1),
    .Y(_1343_)
);

OAI21X1 _2203_ (
    .A(_923__bF$buf3),
    .B(_933_),
    .C(_1045_),
    .Y(_1344_)
);

OAI21X1 _2204_ (
    .A(_923__bF$buf2),
    .B(_1047_),
    .C(_1008_),
    .Y(_1345_)
);

NOR3X1 _2205_ (
    .A(_1343_),
    .B(_1345_),
    .C(_1344_),
    .Y(_1346_)
);

NAND3X1 _2206_ (
    .A(_1337_),
    .B(_1342_),
    .C(_1346_),
    .Y(_1347_)
);

OR2X2 _2207_ (
    .A(_1344_),
    .B(_1345_),
    .Y(_1348_)
);

AOI21X1 _2208_ (
    .A(dst_reg[1]),
    .B(_1343_),
    .C(_1348_),
    .Y(_1349_)
);

OAI21X1 _2209_ (
    .A(_1333_),
    .B(_1347_),
    .C(_1349_),
    .Y(_1350_)
);

INVX2 _2210_ (
    .A(_1350_),
    .Y(_1351_)
);

OAI21X1 _2211_ (
    .A(_1345_),
    .B(_1344_),
    .C(index_y),
    .Y(_1352_)
);

NAND2X1 _2212_ (
    .A(_1337_),
    .B(_1342_),
    .Y(_1353_)
);

AOI21X1 _2213_ (
    .A(dst_reg[0]),
    .B(_1343_),
    .C(_1353_),
    .Y(_1354_)
);

NAND3X1 _2214_ (
    .A(_1347_),
    .B(_1352_),
    .C(_1354_),
    .Y(_1355_)
);

OAI21X1 _2215_ (
    .A(src_reg[0]),
    .B(_1347_),
    .C(_1355_),
    .Y(_1356_)
);

NAND3X1 _2216_ (
    .A(\AXYS[0] [0]),
    .B(_1351_),
    .C(_1356_),
    .Y(_1357_)
);

AND2X2 _2217_ (
    .A(_1354_),
    .B(_1352_),
    .Y(_1358_)
);

INVX1 _2218_ (
    .A(src_reg[0]),
    .Y(_1359_)
);

OR2X2 _2219_ (
    .A(_1347_),
    .B(_1359_),
    .Y(_1360_)
);

AOI21X1 _2220_ (
    .A(_1358_),
    .B(_1360_),
    .C(_1350_),
    .Y(_1361_)
);

NAND2X1 _2221_ (
    .A(\AXYS[1] [0]),
    .B(_1361_),
    .Y(_1362_)
);

OR2X2 _2222_ (
    .A(_1347_),
    .B(_1333_),
    .Y(_1363_)
);

OR2X2 _2223_ (
    .A(_1347_),
    .B(src_reg[0]),
    .Y(_1364_)
);

AOI22X1 _2224_ (
    .A(_1363_),
    .B(_1349_),
    .C(_1355_),
    .D(_1364_),
    .Y(_1365_)
);

AOI22X1 _2225_ (
    .A(_1363_),
    .B(_1349_),
    .C(_1358_),
    .D(_1360_),
    .Y(_1366_)
);

AOI22X1 _2226_ (
    .A(_1365_),
    .B(\AXYS[2] [0]),
    .C(\AXYS[3] [0]),
    .D(_1366_),
    .Y(_1367_)
);

NAND3X1 _2227_ (
    .A(_1357_),
    .B(_1362_),
    .C(_1367_),
    .Y(_1368_)
);

INVX1 _2228_ (
    .A(_1368_),
    .Y(_1369_)
);

OAI21X1 _2229_ (
    .A(state[4]),
    .B(_1047_),
    .C(_855_),
    .Y(_1370_)
);

OR2X2 _2230_ (
    .A(_1370_),
    .B(_1305_),
    .Y(_1371_)
);

NOR2X1 _2231_ (
    .A(_1307_),
    .B(_1371_),
    .Y(_1372_)
);

OAI21X1 _2232_ (
    .A(_854__bF$buf3),
    .B(_900_),
    .C(_1067_),
    .Y(_1373_)
);

AOI21X1 _2233_ (
    .A(_915_),
    .B(_1007_),
    .C(_1001_),
    .Y(_1374_)
);

AND2X2 _2234_ (
    .A(_1374_),
    .B(_1373_),
    .Y(_1375_)
);

INVX1 _2235_ (
    .A(load_only),
    .Y(_1376_)
);

AOI21X1 _2236_ (
    .A(_955_),
    .B(_1376_),
    .C(_1344_),
    .Y(_1377_)
);

NAND3X1 _2237_ (
    .A(_1375_),
    .B(_1377_),
    .C(_1372_),
    .Y(_1378_)
);

INVX2 _2238_ (
    .A(_1378_),
    .Y(_1379_)
);

NOR2X1 _2239_ (
    .A(_1144_),
    .B(_1033_),
    .Y(_1380_)
);

NAND2X1 _2240_ (
    .A(_854__bF$buf2),
    .B(_1157_),
    .Y(_1381_)
);

OAI21X1 _2241_ (
    .A(_917__bF$buf4),
    .B(_1082_),
    .C(_1381_),
    .Y(_1382_)
);

OAI21X1 _2242_ (
    .A(_899__bF$buf4),
    .B(_1082_),
    .C(_1003_),
    .Y(_1383_)
);

NOR2X1 _2243_ (
    .A(_1382_),
    .B(_1383_),
    .Y(_1384_)
);

NAND3X1 _2244_ (
    .A(_1023_),
    .B(_1384_),
    .C(_1380_),
    .Y(_1385_)
);

INVX1 _2245_ (
    .A(ABH[0]),
    .Y(_1386_)
);

AOI21X1 _2246_ (
    .A(_852_),
    .B(_856__bF$buf2),
    .C(_1063_),
    .Y(_1387_)
);

OAI22X1 _2247_ (
    .A(_1386_),
    .B(_1162_),
    .C(_1304_),
    .D(_1387_),
    .Y(_1388_)
);

AOI21X1 _2248_ (
    .A(_1385_),
    .B(ADD[0]),
    .C(_1388_),
    .Y(_1389_)
);

OAI21X1 _2249_ (
    .A(_1379_),
    .B(_1369_),
    .C(_1389_),
    .Y(AI[0])
);

NAND2X1 _2250_ (
    .A(\AXYS[1] [1]),
    .B(_1361_),
    .Y(_1390_)
);

AOI22X1 _2251_ (
    .A(_1365_),
    .B(\AXYS[2] [1]),
    .C(\AXYS[3] [1]),
    .D(_1366_),
    .Y(_1391_)
);

NAND3X1 _2252_ (
    .A(\AXYS[0] [1]),
    .B(_1351_),
    .C(_1356_),
    .Y(_1392_)
);

NAND3X1 _2253_ (
    .A(_1390_),
    .B(_1392_),
    .C(_1391_),
    .Y(_1393_)
);

INVX1 _2254_ (
    .A(_1393_),
    .Y(_1394_)
);

NAND2X1 _2255_ (
    .A(ABH[1]),
    .B(_1039_),
    .Y(_1395_)
);

OAI21X1 _2256_ (
    .A(_1324_),
    .B(_1387_),
    .C(_1395_),
    .Y(_1396_)
);

AOI21X1 _2257_ (
    .A(_1385_),
    .B(ADD[1]),
    .C(_1396_),
    .Y(_1397_)
);

OAI21X1 _2258_ (
    .A(_1379_),
    .B(_1394_),
    .C(_1397_),
    .Y(AI[1])
);

NAND2X1 _2259_ (
    .A(\AXYS[1] [2]),
    .B(_1361_),
    .Y(_1398_)
);

AOI22X1 _2260_ (
    .A(_1365_),
    .B(\AXYS[2] [2]),
    .C(\AXYS[3] [2]),
    .D(_1366_),
    .Y(_1399_)
);

NAND3X1 _2261_ (
    .A(\AXYS[0] [2]),
    .B(_1351_),
    .C(_1356_),
    .Y(_1400_)
);

NAND3X1 _2262_ (
    .A(_1398_),
    .B(_1400_),
    .C(_1399_),
    .Y(_1401_)
);

INVX1 _2263_ (
    .A(_1401_),
    .Y(_1402_)
);

INVX1 _2264_ (
    .A(ABH[2]),
    .Y(_1403_)
);

NOR2X1 _2265_ (
    .A(_1403_),
    .B(_1162_),
    .Y(_1404_)
);

INVX1 _2266_ (
    .A(_1404_),
    .Y(_1405_)
);

OAI21X1 _2267_ (
    .A(_838_),
    .B(_1387_),
    .C(_1405_),
    .Y(_1406_)
);

AOI21X1 _2268_ (
    .A(_1385_),
    .B(ADD[2]),
    .C(_1406_),
    .Y(_1407_)
);

OAI21X1 _2269_ (
    .A(_1379_),
    .B(_1402_),
    .C(_1407_),
    .Y(AI[2])
);

NAND2X1 _2270_ (
    .A(\AXYS[1] [3]),
    .B(_1361_),
    .Y(_1408_)
);

AOI22X1 _2271_ (
    .A(_1365_),
    .B(\AXYS[2] [3]),
    .C(\AXYS[3] [3]),
    .D(_1366_),
    .Y(_1409_)
);

NAND3X1 _2272_ (
    .A(\AXYS[0] [3]),
    .B(_1351_),
    .C(_1356_),
    .Y(_1410_)
);

NAND3X1 _2273_ (
    .A(_1408_),
    .B(_1410_),
    .C(_1409_),
    .Y(_1411_)
);

INVX1 _2274_ (
    .A(_1411_),
    .Y(_1412_)
);

NAND2X1 _2275_ (
    .A(ABH[3]),
    .B(_1039_),
    .Y(_1413_)
);

OAI21X1 _2276_ (
    .A(_1327_),
    .B(_1387_),
    .C(_1413_),
    .Y(_1414_)
);

AOI21X1 _2277_ (
    .A(_1385_),
    .B(ADD[3]),
    .C(_1414_),
    .Y(_1415_)
);

OAI21X1 _2278_ (
    .A(_1379_),
    .B(_1412_),
    .C(_1415_),
    .Y(AI[3])
);

NAND2X1 _2279_ (
    .A(\AXYS[1] [4]),
    .B(_1361_),
    .Y(_1416_)
);

AOI22X1 _2280_ (
    .A(_1365_),
    .B(\AXYS[2] [4]),
    .C(\AXYS[3] [4]),
    .D(_1366_),
    .Y(_1417_)
);

NAND3X1 _2281_ (
    .A(\AXYS[0] [4]),
    .B(_1351_),
    .C(_1356_),
    .Y(_1418_)
);

NAND3X1 _2282_ (
    .A(_1416_),
    .B(_1418_),
    .C(_1417_),
    .Y(_1419_)
);

INVX1 _2283_ (
    .A(_1419_),
    .Y(_1420_)
);

NAND2X1 _2284_ (
    .A(ABH[4]),
    .B(_1039_),
    .Y(_1421_)
);

OAI21X1 _2285_ (
    .A(_1329_),
    .B(_1387_),
    .C(_1421_),
    .Y(_1422_)
);

AOI21X1 _2286_ (
    .A(_1385_),
    .B(ADD[4]),
    .C(_1422_),
    .Y(_1423_)
);

OAI21X1 _2287_ (
    .A(_1379_),
    .B(_1420_),
    .C(_1423_),
    .Y(AI[4])
);

NAND2X1 _2288_ (
    .A(\AXYS[1] [5]),
    .B(_1361_),
    .Y(_1424_)
);

AOI22X1 _2289_ (
    .A(_1365_),
    .B(\AXYS[2] [5]),
    .C(\AXYS[3] [5]),
    .D(_1366_),
    .Y(_1425_)
);

NAND3X1 _2290_ (
    .A(\AXYS[0] [5]),
    .B(_1351_),
    .C(_1356_),
    .Y(_1426_)
);

NAND3X1 _2291_ (
    .A(_1424_),
    .B(_1426_),
    .C(_1425_),
    .Y(_1427_)
);

INVX1 _2292_ (
    .A(_1427_),
    .Y(_1428_)
);

NAND2X1 _2293_ (
    .A(ABH[5]),
    .B(_1039_),
    .Y(_1429_)
);

OAI21X1 _2294_ (
    .A(_844_),
    .B(_1387_),
    .C(_1429_),
    .Y(_1430_)
);

AOI21X1 _2295_ (
    .A(_1385_),
    .B(ADD[5]),
    .C(_1430_),
    .Y(_1431_)
);

OAI21X1 _2296_ (
    .A(_1379_),
    .B(_1428_),
    .C(_1431_),
    .Y(AI[5])
);

NAND2X1 _2297_ (
    .A(\AXYS[1] [6]),
    .B(_1361_),
    .Y(_1432_)
);

AOI22X1 _2298_ (
    .A(_1365_),
    .B(\AXYS[2] [6]),
    .C(\AXYS[3] [6]),
    .D(_1366_),
    .Y(_1433_)
);

NAND3X1 _2299_ (
    .A(\AXYS[0] [6]),
    .B(_1351_),
    .C(_1356_),
    .Y(_1434_)
);

NAND3X1 _2300_ (
    .A(_1432_),
    .B(_1434_),
    .C(_1433_),
    .Y(_1435_)
);

INVX1 _2301_ (
    .A(_1435_),
    .Y(_1436_)
);

INVX1 _2302_ (
    .A(ABH[6]),
    .Y(_1437_)
);

NOR2X1 _2303_ (
    .A(_1437_),
    .B(_1162_),
    .Y(_1438_)
);

INVX1 _2304_ (
    .A(_1438_),
    .Y(_1439_)
);

OAI21X1 _2305_ (
    .A(_846_),
    .B(_1387_),
    .C(_1439_),
    .Y(_1440_)
);

AOI21X1 _2306_ (
    .A(_1385_),
    .B(ADD[6]),
    .C(_1440_),
    .Y(_1441_)
);

OAI21X1 _2307_ (
    .A(_1379_),
    .B(_1436_),
    .C(_1441_),
    .Y(AI[6])
);

NAND2X1 _2308_ (
    .A(\AXYS[1] [7]),
    .B(_1361_),
    .Y(_1442_)
);

AOI22X1 _2309_ (
    .A(_1365_),
    .B(\AXYS[2] [7]),
    .C(\AXYS[3] [7]),
    .D(_1366_),
    .Y(_1443_)
);

NAND3X1 _2310_ (
    .A(\AXYS[0] [7]),
    .B(_1351_),
    .C(_1356_),
    .Y(_1444_)
);

NAND3X1 _2311_ (
    .A(_1442_),
    .B(_1444_),
    .C(_1443_),
    .Y(_1445_)
);

INVX1 _2312_ (
    .A(_1445_),
    .Y(_1446_)
);

INVX1 _2313_ (
    .A(ABH[7]),
    .Y(_1447_)
);

NOR2X1 _2314_ (
    .A(_1447_),
    .B(_1162_),
    .Y(_1448_)
);

INVX1 _2315_ (
    .A(_1448_),
    .Y(_1449_)
);

OAI21X1 _2316_ (
    .A(_847_),
    .B(_1387_),
    .C(_1449_),
    .Y(_1450_)
);

AOI21X1 _2317_ (
    .A(_1385_),
    .B(\ALU.N ),
    .C(_1450_),
    .Y(_1451_)
);

OAI21X1 _2318_ (
    .A(_1379_),
    .B(_1446_),
    .C(_1451_),
    .Y(AI[7])
);

INVX1 _2319_ (
    .A(op[0]),
    .Y(_1452_)
);

OAI21X1 _2320_ (
    .A(_923__bF$buf1),
    .B(_954_),
    .C(_1294_),
    .Y(_1453_)
);

INVX2 _2321_ (
    .A(_1453_),
    .Y(_1454_)
);

NAND3X1 _2322_ (
    .A(_859__bF$buf0),
    .B(_1310_),
    .C(_1454_),
    .Y(_1455_)
);

OAI21X1 _2323_ (
    .A(_1452_),
    .B(_1454_),
    .C(_1455_),
    .Y(\ALU.op [0])
);

INVX1 _2324_ (
    .A(op[1]),
    .Y(_1456_)
);

OAI21X1 _2325_ (
    .A(_1456_),
    .B(_1454_),
    .C(_1455_),
    .Y(\ALU.op [1])
);

INVX1 _2326_ (
    .A(_1001_),
    .Y(_1457_)
);

OAI21X1 _2327_ (
    .A(state[5]),
    .B(_1313_),
    .C(_1457_),
    .Y(_1458_)
);

INVX2 _2328_ (
    .A(_1383_),
    .Y(_1459_)
);

OAI21X1 _2329_ (
    .A(_917__bF$buf3),
    .B(_1047_),
    .C(_1459_),
    .Y(_1460_)
);

NOR2X1 _2330_ (
    .A(_1458_),
    .B(_1460_),
    .Y(_1461_)
);

AOI22X1 _2331_ (
    .A(backwards),
    .B(_1039_),
    .C(_1453_),
    .D(op[2]),
    .Y(_1462_)
);

NAND2X1 _2332_ (
    .A(_1462_),
    .B(_1461_),
    .Y(\ALU.op [2])
);

INVX1 _2333_ (
    .A(op[3]),
    .Y(_117_)
);

NOR2X1 _2334_ (
    .A(_117_),
    .B(_1454_),
    .Y(\ALU.op [3])
);

OAI21X1 _2335_ (
    .A(_917__bF$buf2),
    .B(_933_),
    .C(_1461_),
    .Y(_118_)
);

INVX1 _2336_ (
    .A(_118_),
    .Y(_119_)
);

INVX1 _2337_ (
    .A(_901_),
    .Y(_120_)
);

OAI21X1 _2338_ (
    .A(_914_),
    .B(_913_),
    .C(_928_),
    .Y(_121_)
);

OAI21X1 _2339_ (
    .A(_120_),
    .B(_121_),
    .C(store),
    .Y(_122_)
);

NAND2X1 _2340_ (
    .A(_122_),
    .B(_119_),
    .Y(_1667_)
);

INVX1 _2341_ (
    .A(PC[8]),
    .Y(_123_)
);

OAI21X1 _2342_ (
    .A(_923__bF$buf0),
    .B(_990_),
    .C(_1080_),
    .Y(_124_)
);

INVX2 _2343_ (
    .A(_124_),
    .Y(_125_)
);

OAI21X1 _2344_ (
    .A(php),
    .B(_1317_),
    .C(_935_),
    .Y(_126_)
);

INVX1 _2345_ (
    .A(php),
    .Y(_127_)
);

OAI21X1 _2346_ (
    .A(_127_),
    .B(_1317_),
    .C(_1074__bF$buf1),
    .Y(_128_)
);

NAND2X1 _2347_ (
    .A(C),
    .B(_128_),
    .Y(_129_)
);

OAI21X1 _2348_ (
    .A(_1303_),
    .B(_1459_),
    .C(_129_),
    .Y(_130_)
);

AOI21X1 _2349_ (
    .A(ADD[0]),
    .B(_126_),
    .C(_130_),
    .Y(_131_)
);

OAI21X1 _2350_ (
    .A(_123_),
    .B(_125_),
    .C(_131_),
    .Y(_132_)
);

INVX1 _2351_ (
    .A(_132_),
    .Y(_133_)
);

OAI21X1 _2352_ (
    .A(_118_),
    .B(_1369_),
    .C(_133_),
    .Y(_1666_[0])
);

INVX1 _2353_ (
    .A(PC[9]),
    .Y(_134_)
);

NAND2X1 _2354_ (
    .A(Z),
    .B(_128_),
    .Y(_135_)
);

OAI21X1 _2355_ (
    .A(_134_),
    .B(_125_),
    .C(_135_),
    .Y(_136_)
);

AOI21X1 _2356_ (
    .A(ADD[1]),
    .B(_126_),
    .C(_136_),
    .Y(_137_)
);

OAI21X1 _2357_ (
    .A(_1323_),
    .B(_1459_),
    .C(_137_),
    .Y(_138_)
);

INVX1 _2358_ (
    .A(_138_),
    .Y(_139_)
);

OAI21X1 _2359_ (
    .A(_118_),
    .B(_1394_),
    .C(_139_),
    .Y(_1666_[1])
);

INVX1 _2360_ (
    .A(PC[10]),
    .Y(_140_)
);

NAND2X1 _2361_ (
    .A(I),
    .B(_128_),
    .Y(_141_)
);

OAI21X1 _2362_ (
    .A(_140_),
    .B(_125_),
    .C(_141_),
    .Y(_142_)
);

AOI21X1 _2363_ (
    .A(ADD[2]),
    .B(_126_),
    .C(_142_),
    .Y(_143_)
);

OAI21X1 _2364_ (
    .A(_1325_),
    .B(_1459_),
    .C(_143_),
    .Y(_144_)
);

INVX1 _2365_ (
    .A(_144_),
    .Y(_145_)
);

OAI21X1 _2366_ (
    .A(_118_),
    .B(_1402_),
    .C(_145_),
    .Y(_1666_[2])
);

INVX1 _2367_ (
    .A(PC[11]),
    .Y(_146_)
);

NAND2X1 _2368_ (
    .A(D),
    .B(_128_),
    .Y(_147_)
);

OAI21X1 _2369_ (
    .A(_146_),
    .B(_125_),
    .C(_147_),
    .Y(_148_)
);

AOI21X1 _2370_ (
    .A(ADD[3]),
    .B(_126_),
    .C(_148_),
    .Y(_149_)
);

OAI21X1 _2371_ (
    .A(_1326_),
    .B(_1459_),
    .C(_149_),
    .Y(_150_)
);

INVX1 _2372_ (
    .A(_150_),
    .Y(_151_)
);

OAI21X1 _2373_ (
    .A(_118_),
    .B(_1412_),
    .C(_151_),
    .Y(_1666_[3])
);

INVX1 _2374_ (
    .A(PC[12]),
    .Y(_152_)
);

OAI21X1 _2375_ (
    .A(_917__bF$buf1),
    .B(_933_),
    .C(_1317_),
    .Y(_153_)
);

OAI22X1 _2376_ (
    .A(_867_),
    .B(_1074__bF$buf0),
    .C(_127_),
    .D(_1317_),
    .Y(_154_)
);

AOI21X1 _2377_ (
    .A(ADD[4]),
    .B(_153_),
    .C(_154_),
    .Y(_155_)
);

OAI21X1 _2378_ (
    .A(_1328_),
    .B(_1459_),
    .C(_155_),
    .Y(_156_)
);

AOI21X1 _2379_ (
    .A(_1419_),
    .B(_119_),
    .C(_156_),
    .Y(_157_)
);

OAI21X1 _2380_ (
    .A(_152_),
    .B(_125_),
    .C(_157_),
    .Y(_1666_[4])
);

AOI22X1 _2381_ (
    .A(PC[13]),
    .B(_124_),
    .C(_153_),
    .D(ADD[5]),
    .Y(_158_)
);

OAI21X1 _2382_ (
    .A(_1330_),
    .B(_1459_),
    .C(_158_),
    .Y(_159_)
);

NOR2X1 _2383_ (
    .A(_128_),
    .B(_159_),
    .Y(_160_)
);

OAI21X1 _2384_ (
    .A(_118_),
    .B(_1428_),
    .C(_160_),
    .Y(_1666_[5])
);

INVX1 _2385_ (
    .A(PC[14]),
    .Y(_161_)
);

NAND2X1 _2386_ (
    .A(V),
    .B(_128_),
    .Y(_162_)
);

OAI21X1 _2387_ (
    .A(_1331_),
    .B(_1459_),
    .C(_162_),
    .Y(_163_)
);

AOI21X1 _2388_ (
    .A(ADD[6]),
    .B(_126_),
    .C(_163_),
    .Y(_164_)
);

OAI21X1 _2389_ (
    .A(_161_),
    .B(_125_),
    .C(_164_),
    .Y(_165_)
);

INVX1 _2390_ (
    .A(_165_),
    .Y(_166_)
);

OAI21X1 _2391_ (
    .A(_118_),
    .B(_1436_),
    .C(_166_),
    .Y(_1666_[6])
);

INVX1 _2392_ (
    .A(PC[15]),
    .Y(_167_)
);

NAND2X1 _2393_ (
    .A(N),
    .B(_128_),
    .Y(_168_)
);

OAI21X1 _2394_ (
    .A(_1332_),
    .B(_1459_),
    .C(_168_),
    .Y(_169_)
);

AOI21X1 _2395_ (
    .A(\ALU.N ),
    .B(_126_),
    .C(_169_),
    .Y(_170_)
);

OAI21X1 _2396_ (
    .A(_167_),
    .B(_125_),
    .C(_170_),
    .Y(_171_)
);

INVX1 _2397_ (
    .A(_171_),
    .Y(_172_)
);

OAI21X1 _2398_ (
    .A(_118_),
    .B(_1446_),
    .C(_172_),
    .Y(_1666_[7])
);

OAI21X1 _2399_ (
    .A(_917__bF$buf0),
    .B(_1047_),
    .C(_1288_),
    .Y(_173_)
);

NOR2X1 _2400_ (
    .A(_124_),
    .B(_173_),
    .Y(_174_)
);

INVX2 _2401_ (
    .A(_174_),
    .Y(_175_)
);

OAI21X1 _2402_ (
    .A(_950_),
    .B(_1339_),
    .C(_854__bF$buf1),
    .Y(_176_)
);

AND2X2 _2403_ (
    .A(_176_),
    .B(_1232_),
    .Y(_177_)
);

NAND3X1 _2404_ (
    .A(_1384_),
    .B(_177_),
    .C(_1380_),
    .Y(_178_)
);

AOI21X1 _2405_ (
    .A(_1009_),
    .B(_915_),
    .C(_1227_),
    .Y(_179_)
);

NAND3X1 _2406_ (
    .A(_1023_),
    .B(_1045_),
    .C(_179_),
    .Y(_180_)
);

NOR2X1 _2407_ (
    .A(_180_),
    .B(_178_),
    .Y(_181_)
);

AOI21X1 _2408_ (
    .A(_853_),
    .B(_1009_),
    .C(_906_),
    .Y(_182_)
);

OAI21X1 _2409_ (
    .A(_923__bF$buf3),
    .B(_1062_),
    .C(_182_),
    .Y(_183_)
);

OAI21X1 _2410_ (
    .A(_854__bF$buf0),
    .B(_900_),
    .C(_996_),
    .Y(_184_)
);

OAI21X1 _2411_ (
    .A(_899__bF$buf3),
    .B(_1035_),
    .C(_184_),
    .Y(_185_)
);

NOR2X1 _2412_ (
    .A(_185_),
    .B(_183_),
    .Y(_186_)
);

OAI21X1 _2413_ (
    .A(_923__bF$buf2),
    .B(_1029_),
    .C(_186_),
    .Y(_187_)
);

OAI21X1 _2414_ (
    .A(_917__bF$buf4),
    .B(_933_),
    .C(_1294_),
    .Y(_188_)
);

INVX2 _2415_ (
    .A(_188_),
    .Y(_189_)
);

INVX1 _2416_ (
    .A(_922_),
    .Y(_190_)
);

OAI21X1 _2417_ (
    .A(_899__bF$buf2),
    .B(_1047_),
    .C(_190_),
    .Y(_191_)
);

NAND2X1 _2418_ (
    .A(_856__bF$buf1),
    .B(_1157_),
    .Y(_192_)
);

NAND3X1 _2419_ (
    .A(_192_),
    .B(_901_),
    .C(_926_),
    .Y(_193_)
);

NOR2X1 _2420_ (
    .A(_193_),
    .B(_191_),
    .Y(_194_)
);

NAND3X1 _2421_ (
    .A(_174_),
    .B(_189_),
    .C(_194_),
    .Y(_195_)
);

NOR2X1 _2422_ (
    .A(_195_),
    .B(_187_),
    .Y(_196_)
);

NAND2X1 _2423_ (
    .A(_181_),
    .B(_196_),
    .Y(_197_)
);

NAND2X1 _2424_ (
    .A(_186_),
    .B(_181_),
    .Y(_198_)
);

INVX1 _2425_ (
    .A(ABL[0]),
    .Y(_199_)
);

NOR2X1 _2426_ (
    .A(_193_),
    .B(_188_),
    .Y(_200_)
);

AOI22X1 _2427_ (
    .A(ADD[0]),
    .B(_1039_),
    .C(_191_),
    .D(DIMUX[0]),
    .Y(_201_)
);

OAI21X1 _2428_ (
    .A(_199_),
    .B(_200_),
    .C(_201_),
    .Y(_202_)
);

AOI21X1 _2429_ (
    .A(_198_),
    .B(ADD[0]),
    .C(_202_),
    .Y(_203_)
);

OAI21X1 _2430_ (
    .A(_1303_),
    .B(_197_),
    .C(_203_),
    .Y(_204_)
);

AOI21X1 _2431_ (
    .A(_1368_),
    .B(_175_),
    .C(_204_),
    .Y(_205_)
);

INVX1 _2432_ (
    .A(_205_),
    .Y(_1665_[0])
);

OR2X2 _2433_ (
    .A(_198_),
    .B(_1039_),
    .Y(_206_)
);

INVX2 _2434_ (
    .A(_191_),
    .Y(_207_)
);

OAI21X1 _2435_ (
    .A(_193_),
    .B(_188_),
    .C(ABL[1]),
    .Y(_208_)
);

OAI21X1 _2436_ (
    .A(_1324_),
    .B(_207_),
    .C(_208_),
    .Y(_209_)
);

AOI21X1 _2437_ (
    .A(_206_),
    .B(ADD[1]),
    .C(_209_),
    .Y(_210_)
);

OAI21X1 _2438_ (
    .A(_1323_),
    .B(_197_),
    .C(_210_),
    .Y(_211_)
);

AOI21X1 _2439_ (
    .A(_1393_),
    .B(_175_),
    .C(_211_),
    .Y(_212_)
);

INVX1 _2440_ (
    .A(_212_),
    .Y(_1665_[1])
);

OAI21X1 _2441_ (
    .A(_193_),
    .B(_188_),
    .C(ABL[2]),
    .Y(_213_)
);

OAI21X1 _2442_ (
    .A(_838_),
    .B(_207_),
    .C(_213_),
    .Y(_214_)
);

AOI21X1 _2443_ (
    .A(_206_),
    .B(ADD[2]),
    .C(_214_),
    .Y(_215_)
);

OAI21X1 _2444_ (
    .A(_1325_),
    .B(_197_),
    .C(_215_),
    .Y(_216_)
);

AOI21X1 _2445_ (
    .A(_1401_),
    .B(_175_),
    .C(_216_),
    .Y(_217_)
);

INVX1 _2446_ (
    .A(_217_),
    .Y(_1665_[2])
);

INVX1 _2447_ (
    .A(ABL[3]),
    .Y(_218_)
);

OAI22X1 _2448_ (
    .A(_218_),
    .B(_200_),
    .C(_1327_),
    .D(_207_),
    .Y(_219_)
);

AOI21X1 _2449_ (
    .A(_206_),
    .B(ADD[3]),
    .C(_219_),
    .Y(_220_)
);

OAI21X1 _2450_ (
    .A(_1326_),
    .B(_197_),
    .C(_220_),
    .Y(_221_)
);

AOI21X1 _2451_ (
    .A(_1411_),
    .B(_175_),
    .C(_221_),
    .Y(_222_)
);

INVX1 _2452_ (
    .A(_222_),
    .Y(_1665_[3])
);

INVX1 _2453_ (
    .A(ABL[4]),
    .Y(_223_)
);

AOI22X1 _2454_ (
    .A(ADD[4]),
    .B(_1039_),
    .C(_191_),
    .D(DIMUX[4]),
    .Y(_224_)
);

OAI21X1 _2455_ (
    .A(_223_),
    .B(_200_),
    .C(_224_),
    .Y(_225_)
);

AOI21X1 _2456_ (
    .A(_198_),
    .B(ADD[4]),
    .C(_225_),
    .Y(_226_)
);

OAI21X1 _2457_ (
    .A(_1328_),
    .B(_197_),
    .C(_226_),
    .Y(_227_)
);

AOI21X1 _2458_ (
    .A(_1419_),
    .B(_175_),
    .C(_227_),
    .Y(_228_)
);

INVX1 _2459_ (
    .A(_228_),
    .Y(_1665_[4])
);

INVX1 _2460_ (
    .A(ABL[5]),
    .Y(_229_)
);

OAI22X1 _2461_ (
    .A(_229_),
    .B(_200_),
    .C(_844_),
    .D(_207_),
    .Y(_230_)
);

AOI21X1 _2462_ (
    .A(_206_),
    .B(ADD[5]),
    .C(_230_),
    .Y(_231_)
);

OAI21X1 _2463_ (
    .A(_1330_),
    .B(_197_),
    .C(_231_),
    .Y(_232_)
);

AOI21X1 _2464_ (
    .A(_1427_),
    .B(_175_),
    .C(_232_),
    .Y(_233_)
);

INVX1 _2465_ (
    .A(_233_),
    .Y(_1665_[5])
);

INVX1 _2466_ (
    .A(ABL[6]),
    .Y(_234_)
);

OAI22X1 _2467_ (
    .A(_846_),
    .B(_207_),
    .C(_234_),
    .D(_200_),
    .Y(_235_)
);

AOI21X1 _2468_ (
    .A(_206_),
    .B(ADD[6]),
    .C(_235_),
    .Y(_236_)
);

OAI21X1 _2469_ (
    .A(_1331_),
    .B(_197_),
    .C(_236_),
    .Y(_237_)
);

AOI21X1 _2470_ (
    .A(_1435_),
    .B(_175_),
    .C(_237_),
    .Y(_238_)
);

INVX1 _2471_ (
    .A(_238_),
    .Y(_1665_[6])
);

INVX1 _2472_ (
    .A(ABL[7]),
    .Y(_239_)
);

OAI22X1 _2473_ (
    .A(_239_),
    .B(_200_),
    .C(_847_),
    .D(_207_),
    .Y(_240_)
);

AOI21X1 _2474_ (
    .A(_206_),
    .B(\ALU.N ),
    .C(_240_),
    .Y(_241_)
);

OAI21X1 _2475_ (
    .A(_1332_),
    .B(_197_),
    .C(_241_),
    .Y(_242_)
);

AOI21X1 _2476_ (
    .A(_1445_),
    .B(_175_),
    .C(_242_),
    .Y(_243_)
);

INVX1 _2477_ (
    .A(_243_),
    .Y(_1665_[7])
);

OAI21X1 _2478_ (
    .A(_1386_),
    .B(_189_),
    .C(_174_),
    .Y(_244_)
);

AOI22X1 _2479_ (
    .A(ABH[0]),
    .B(_1039_),
    .C(_193_),
    .D(ADD[0]),
    .Y(_245_)
);

OAI21X1 _2480_ (
    .A(_1304_),
    .B(_186_),
    .C(_245_),
    .Y(_246_)
);

NOR3X1 _2481_ (
    .A(_244_),
    .B(_246_),
    .C(_178_),
    .Y(_247_)
);

OAI21X1 _2482_ (
    .A(_123_),
    .B(_197_),
    .C(_247_),
    .Y(_1665_[8])
);

OAI21X1 _2483_ (
    .A(_185_),
    .B(_183_),
    .C(DIMUX[1]),
    .Y(_248_)
);

INVX1 _2484_ (
    .A(_248_),
    .Y(_249_)
);

INVX1 _2485_ (
    .A(ABH[1]),
    .Y(_250_)
);

AOI22X1 _2486_ (
    .A(ABH[1]),
    .B(_1039_),
    .C(_193_),
    .D(ADD[1]),
    .Y(_251_)
);

OAI21X1 _2487_ (
    .A(_250_),
    .B(_189_),
    .C(_251_),
    .Y(_252_)
);

NOR2X1 _2488_ (
    .A(_252_),
    .B(_249_),
    .Y(_253_)
);

OAI21X1 _2489_ (
    .A(_134_),
    .B(_197_),
    .C(_253_),
    .Y(_1665_[9])
);

OAI21X1 _2490_ (
    .A(_185_),
    .B(_183_),
    .C(DIMUX[2]),
    .Y(_254_)
);

INVX1 _2491_ (
    .A(_254_),
    .Y(_255_)
);

AOI21X1 _2492_ (
    .A(_193_),
    .B(ADD[2]),
    .C(_1404_),
    .Y(_256_)
);

OAI21X1 _2493_ (
    .A(_1403_),
    .B(_189_),
    .C(_256_),
    .Y(_257_)
);

NOR2X1 _2494_ (
    .A(_257_),
    .B(_255_),
    .Y(_258_)
);

OAI21X1 _2495_ (
    .A(_140_),
    .B(_197_),
    .C(_258_),
    .Y(_1665_[10])
);

OAI21X1 _2496_ (
    .A(_185_),
    .B(_183_),
    .C(DIMUX[3]),
    .Y(_259_)
);

INVX1 _2497_ (
    .A(_259_),
    .Y(_260_)
);

INVX1 _2498_ (
    .A(ABH[3]),
    .Y(_261_)
);

AOI22X1 _2499_ (
    .A(ABH[3]),
    .B(_1039_),
    .C(_193_),
    .D(ADD[3]),
    .Y(_262_)
);

OAI21X1 _2500_ (
    .A(_261_),
    .B(_189_),
    .C(_262_),
    .Y(_263_)
);

NOR2X1 _2501_ (
    .A(_263_),
    .B(_260_),
    .Y(_264_)
);

OAI21X1 _2502_ (
    .A(_146_),
    .B(_197_),
    .C(_264_),
    .Y(_1665_[11])
);

INVX1 _2503_ (
    .A(ABH[4]),
    .Y(_265_)
);

NAND2X1 _2504_ (
    .A(ADD[4]),
    .B(_193_),
    .Y(_266_)
);

OAI21X1 _2505_ (
    .A(_265_),
    .B(_189_),
    .C(_266_),
    .Y(_267_)
);

OAI21X1 _2506_ (
    .A(_185_),
    .B(_183_),
    .C(DIMUX[4]),
    .Y(_268_)
);

OAI21X1 _2507_ (
    .A(_265_),
    .B(_1162_),
    .C(_268_),
    .Y(_269_)
);

NOR2X1 _2508_ (
    .A(_267_),
    .B(_269_),
    .Y(_270_)
);

OAI21X1 _2509_ (
    .A(_152_),
    .B(_197_),
    .C(_270_),
    .Y(_1665_[12])
);

INVX1 _2510_ (
    .A(PC[13]),
    .Y(_271_)
);

OAI21X1 _2511_ (
    .A(_185_),
    .B(_183_),
    .C(DIMUX[5]),
    .Y(_272_)
);

INVX1 _2512_ (
    .A(_272_),
    .Y(_273_)
);

INVX1 _2513_ (
    .A(ABH[5]),
    .Y(_274_)
);

AOI22X1 _2514_ (
    .A(ABH[5]),
    .B(_1039_),
    .C(_193_),
    .D(ADD[5]),
    .Y(_275_)
);

OAI21X1 _2515_ (
    .A(_274_),
    .B(_189_),
    .C(_275_),
    .Y(_276_)
);

NOR2X1 _2516_ (
    .A(_276_),
    .B(_273_),
    .Y(_277_)
);

OAI21X1 _2517_ (
    .A(_271_),
    .B(_197_),
    .C(_277_),
    .Y(_1665_[13])
);

OAI21X1 _2518_ (
    .A(_185_),
    .B(_183_),
    .C(DIMUX[6]),
    .Y(_278_)
);

INVX1 _2519_ (
    .A(_278_),
    .Y(_279_)
);

AOI21X1 _2520_ (
    .A(_193_),
    .B(ADD[6]),
    .C(_1438_),
    .Y(_280_)
);

OAI21X1 _2521_ (
    .A(_1437_),
    .B(_189_),
    .C(_280_),
    .Y(_281_)
);

NOR2X1 _2522_ (
    .A(_281_),
    .B(_279_),
    .Y(_282_)
);

OAI21X1 _2523_ (
    .A(_161_),
    .B(_197_),
    .C(_282_),
    .Y(_1665_[14])
);

OAI21X1 _2524_ (
    .A(_185_),
    .B(_183_),
    .C(DIMUX[7]),
    .Y(_283_)
);

INVX1 _2525_ (
    .A(_283_),
    .Y(_284_)
);

AOI21X1 _2526_ (
    .A(_193_),
    .B(\ALU.N ),
    .C(_1448_),
    .Y(_285_)
);

OAI21X1 _2527_ (
    .A(_1447_),
    .B(_189_),
    .C(_285_),
    .Y(_286_)
);

NOR2X1 _2528_ (
    .A(_286_),
    .B(_284_),
    .Y(_287_)
);

OAI21X1 _2529_ (
    .A(_167_),
    .B(_197_),
    .C(_287_),
    .Y(_1665_[15])
);

AND2X2 _2530_ (
    .A(adc_sbc),
    .B(D),
    .Y(_0_)
);

AND2X2 _2531_ (
    .A(_955_),
    .B(adc_bcd),
    .Y(\ALU.BCD )
);

INVX1 _2532_ (
    .A(shift_right),
    .Y(_288_)
);

NOR2X1 _2533_ (
    .A(_288_),
    .B(_1454_),
    .Y(\ALU.right )
);

INVX8 _2534_ (
    .A(reset),
    .Y(_1_)
);

OAI21X1 _2535_ (
    .A(_923__bF$buf1),
    .B(_1047_),
    .C(_184_),
    .Y(_289_)
);

NOR2X1 _2536_ (
    .A(_874_),
    .B(_859__bF$buf3),
    .Y(_290_)
);

NAND2X1 _2537_ (
    .A(_853_),
    .B(_1157_),
    .Y(_291_)
);

OAI21X1 _2538_ (
    .A(state[4]),
    .B(_954_),
    .C(_291_),
    .Y(_292_)
);

NOR3X1 _2539_ (
    .A(_290_),
    .B(_292_),
    .C(_289_),
    .Y(_293_)
);

NAND3X1 _2540_ (
    .A(_1075_),
    .B(_986_),
    .C(_1231_),
    .Y(_294_)
);

NOR2X1 _2541_ (
    .A(_1163_),
    .B(_294_),
    .Y(_295_)
);

NAND2X1 _2542_ (
    .A(_295_),
    .B(_293_),
    .Y(_296_)
);

NAND2X1 _2543_ (
    .A(_900_),
    .B(_1157_),
    .Y(_297_)
);

OAI22X1 _2544_ (
    .A(_854__bF$buf3),
    .B(_900_),
    .C(_938_),
    .D(_996_),
    .Y(_298_)
);

NAND3X1 _2545_ (
    .A(_297_),
    .B(_1162_),
    .C(_298_),
    .Y(_299_)
);

NAND3X1 _2546_ (
    .A(_859__bF$buf2),
    .B(_192_),
    .C(_1074__bF$buf3),
    .Y(_300_)
);

NAND3X1 _2547_ (
    .A(_856__bF$buf0),
    .B(_950_),
    .C(_868_),
    .Y(_301_)
);

OAI21X1 _2548_ (
    .A(_923__bF$buf0),
    .B(_1035_),
    .C(_301_),
    .Y(_302_)
);

INVX1 _2549_ (
    .A(_302_),
    .Y(_303_)
);

OAI21X1 _2550_ (
    .A(_300_),
    .B(_299_),
    .C(_303_),
    .Y(_304_)
);

INVX2 _2551_ (
    .A(_304_),
    .Y(_305_)
);

NOR2X1 _2552_ (
    .A(_859__bF$buf1),
    .B(_868_),
    .Y(_306_)
);

AOI22X1 _2553_ (
    .A(ABL[0]),
    .B(_306_),
    .C(_299_),
    .D(ADD[0]),
    .Y(_307_)
);

OAI21X1 _2554_ (
    .A(_1303_),
    .B(_305_),
    .C(_307_),
    .Y(_308_)
);

NOR2X1 _2555_ (
    .A(_296_),
    .B(_308_),
    .Y(_309_)
);

NAND2X1 _2556_ (
    .A(PC[0]),
    .B(_304_),
    .Y(_310_)
);

AOI22X1 _2557_ (
    .A(_293_),
    .B(_295_),
    .C(_310_),
    .D(_307_),
    .Y(_311_)
);

INVX1 _2558_ (
    .A(_311_),
    .Y(_312_)
);

NAND2X1 _2559_ (
    .A(RDY_bF$buf7),
    .B(_312_),
    .Y(_313_)
);

OAI22X1 _2560_ (
    .A(RDY_bF$buf6),
    .B(_1303_),
    .C(_309_),
    .D(_313_),
    .Y(_2_)
);

OAI21X1 _2561_ (
    .A(_899__bF$buf1),
    .B(_1035_),
    .C(_298_),
    .Y(_314_)
);

OAI21X1 _2562_ (
    .A(_1039_),
    .B(_314_),
    .C(ADD[1]),
    .Y(_315_)
);

INVX1 _2563_ (
    .A(res),
    .Y(_316_)
);

AOI22X1 _2564_ (
    .A(ABL[1]),
    .B(_306_),
    .C(_1144_),
    .D(_316_),
    .Y(_317_)
);

AND2X2 _2565_ (
    .A(_315_),
    .B(_317_),
    .Y(_318_)
);

OAI21X1 _2566_ (
    .A(_1323_),
    .B(_305_),
    .C(_318_),
    .Y(_319_)
);

NOR2X1 _2567_ (
    .A(_311_),
    .B(_319_),
    .Y(_320_)
);

NAND2X1 _2568_ (
    .A(_311_),
    .B(_319_),
    .Y(_321_)
);

NAND2X1 _2569_ (
    .A(RDY_bF$buf5),
    .B(_321_),
    .Y(_322_)
);

OAI22X1 _2570_ (
    .A(RDY_bF$buf4),
    .B(_1323_),
    .C(_320_),
    .D(_322_),
    .Y(_3_)
);

NAND2X1 _2571_ (
    .A(PC[2]),
    .B(_836__bF$buf1),
    .Y(_323_)
);

NOR2X1 _2572_ (
    .A(res),
    .B(_866_),
    .Y(_324_)
);

NAND2X1 _2573_ (
    .A(ABL[2]),
    .B(_306_),
    .Y(_325_)
);

OAI21X1 _2574_ (
    .A(_1074__bF$buf2),
    .B(_324_),
    .C(_325_),
    .Y(_326_)
);

AOI21X1 _2575_ (
    .A(ADD[2]),
    .B(_299_),
    .C(_326_),
    .Y(_327_)
);

OAI21X1 _2576_ (
    .A(_1325_),
    .B(_305_),
    .C(_327_),
    .Y(_328_)
);

XOR2X1 _2577_ (
    .A(_321_),
    .B(_328_),
    .Y(_329_)
);

OAI21X1 _2578_ (
    .A(_836__bF$buf0),
    .B(_329_),
    .C(_323_),
    .Y(_4_)
);

INVX1 _2579_ (
    .A(_321_),
    .Y(_330_)
);

INVX2 _2580_ (
    .A(_306_),
    .Y(_331_)
);

OAI21X1 _2581_ (
    .A(_218_),
    .B(_331_),
    .C(_1074__bF$buf1),
    .Y(_332_)
);

AOI21X1 _2582_ (
    .A(ADD[3]),
    .B(_299_),
    .C(_332_),
    .Y(_333_)
);

OAI21X1 _2583_ (
    .A(_1326_),
    .B(_305_),
    .C(_333_),
    .Y(_334_)
);

AOI21X1 _2584_ (
    .A(_330_),
    .B(_328_),
    .C(_334_),
    .Y(_335_)
);

NAND2X1 _2585_ (
    .A(PC[2]),
    .B(_304_),
    .Y(_336_)
);

NAND2X1 _2586_ (
    .A(PC[3]),
    .B(_304_),
    .Y(_337_)
);

AOI22X1 _2587_ (
    .A(_336_),
    .B(_327_),
    .C(_337_),
    .D(_333_),
    .Y(_338_)
);

NAND3X1 _2588_ (
    .A(_311_),
    .B(_319_),
    .C(_338_),
    .Y(_339_)
);

NAND2X1 _2589_ (
    .A(RDY_bF$buf3),
    .B(_339_),
    .Y(_340_)
);

OAI22X1 _2590_ (
    .A(RDY_bF$buf2),
    .B(_1326_),
    .C(_340_),
    .D(_335_),
    .Y(_5_)
);

NAND2X1 _2591_ (
    .A(PC[4]),
    .B(_836__bF$buf7),
    .Y(_341_)
);

OAI21X1 _2592_ (
    .A(_223_),
    .B(_331_),
    .C(_1074__bF$buf0),
    .Y(_342_)
);

AOI21X1 _2593_ (
    .A(ADD[4]),
    .B(_299_),
    .C(_342_),
    .Y(_343_)
);

OAI21X1 _2594_ (
    .A(_1328_),
    .B(_305_),
    .C(_343_),
    .Y(_344_)
);

XOR2X1 _2595_ (
    .A(_339_),
    .B(_344_),
    .Y(_345_)
);

OAI21X1 _2596_ (
    .A(_836__bF$buf6),
    .B(_345_),
    .C(_341_),
    .Y(_6_)
);

INVX1 _2597_ (
    .A(_339_),
    .Y(_346_)
);

OAI21X1 _2598_ (
    .A(_229_),
    .B(_331_),
    .C(_1074__bF$buf3),
    .Y(_347_)
);

AOI21X1 _2599_ (
    .A(ADD[5]),
    .B(_299_),
    .C(_347_),
    .Y(_348_)
);

OAI21X1 _2600_ (
    .A(_1330_),
    .B(_305_),
    .C(_348_),
    .Y(_349_)
);

AOI21X1 _2601_ (
    .A(_346_),
    .B(_344_),
    .C(_349_),
    .Y(_350_)
);

NAND2X1 _2602_ (
    .A(PC[4]),
    .B(_304_),
    .Y(_351_)
);

NAND2X1 _2603_ (
    .A(PC[5]),
    .B(_304_),
    .Y(_352_)
);

AOI22X1 _2604_ (
    .A(_351_),
    .B(_343_),
    .C(_352_),
    .D(_348_),
    .Y(_353_)
);

INVX1 _2605_ (
    .A(_353_),
    .Y(_354_)
);

OAI21X1 _2606_ (
    .A(_354_),
    .B(_339_),
    .C(RDY_bF$buf1),
    .Y(_355_)
);

OAI22X1 _2607_ (
    .A(RDY_bF$buf0),
    .B(_1330_),
    .C(_355_),
    .D(_350_),
    .Y(_7_)
);

OAI21X1 _2608_ (
    .A(_234_),
    .B(_331_),
    .C(_1074__bF$buf2),
    .Y(_356_)
);

AOI21X1 _2609_ (
    .A(ADD[6]),
    .B(_299_),
    .C(_356_),
    .Y(_357_)
);

OAI21X1 _2610_ (
    .A(_1331_),
    .B(_305_),
    .C(_357_),
    .Y(_358_)
);

AOI21X1 _2611_ (
    .A(_346_),
    .B(_353_),
    .C(_358_),
    .Y(_359_)
);

NAND3X1 _2612_ (
    .A(_353_),
    .B(_358_),
    .C(_346_),
    .Y(_360_)
);

NAND2X1 _2613_ (
    .A(RDY_bF$buf8),
    .B(_360_),
    .Y(_361_)
);

OAI22X1 _2614_ (
    .A(RDY_bF$buf7),
    .B(_1331_),
    .C(_359_),
    .D(_361_),
    .Y(_8_)
);

NAND2X1 _2615_ (
    .A(PC[7]),
    .B(_836__bF$buf5),
    .Y(_362_)
);

OAI21X1 _2616_ (
    .A(_239_),
    .B(_331_),
    .C(_1074__bF$buf1),
    .Y(_363_)
);

AOI21X1 _2617_ (
    .A(\ALU.N ),
    .B(_299_),
    .C(_363_),
    .Y(_364_)
);

OAI21X1 _2618_ (
    .A(_1332_),
    .B(_305_),
    .C(_364_),
    .Y(_365_)
);

XOR2X1 _2619_ (
    .A(_360_),
    .B(_365_),
    .Y(_366_)
);

OAI21X1 _2620_ (
    .A(_836__bF$buf4),
    .B(_366_),
    .C(_362_),
    .Y(_9_)
);

AOI21X1 _2621_ (
    .A(_298_),
    .B(_297_),
    .C(_1304_),
    .Y(_367_)
);

OAI22X1 _2622_ (
    .A(_1386_),
    .B(_1162_),
    .C(_123_),
    .D(_301_),
    .Y(_368_)
);

NAND3X1 _2623_ (
    .A(ADD[0]),
    .B(_856__bF$buf3),
    .C(_1157_),
    .Y(_369_)
);

NAND3X1 _2624_ (
    .A(ABH[0]),
    .B(_874_),
    .C(_1343_),
    .Y(_370_)
);

NAND3X1 _2625_ (
    .A(_1074__bF$buf0),
    .B(_369_),
    .C(_370_),
    .Y(_371_)
);

NOR3X1 _2626_ (
    .A(_368_),
    .B(_371_),
    .C(_367_),
    .Y(_372_)
);

AOI22X1 _2627_ (
    .A(_917__bF$buf3),
    .B(_899__bF$buf0),
    .C(_992_),
    .D(_954_),
    .Y(_373_)
);

NOR3X1 _2628_ (
    .A(_1031_),
    .B(_1039_),
    .C(_373_),
    .Y(_374_)
);

INVX1 _2629_ (
    .A(_300_),
    .Y(_375_)
);

NAND3X1 _2630_ (
    .A(PC[8]),
    .B(_375_),
    .C(_374_),
    .Y(_376_)
);

AND2X2 _2631_ (
    .A(_372_),
    .B(_376_),
    .Y(_377_)
);

NAND2X1 _2632_ (
    .A(PC[6]),
    .B(_304_),
    .Y(_378_)
);

NAND2X1 _2633_ (
    .A(PC[7]),
    .B(_304_),
    .Y(_379_)
);

AOI22X1 _2634_ (
    .A(_378_),
    .B(_357_),
    .C(_379_),
    .D(_364_),
    .Y(_380_)
);

NAND2X1 _2635_ (
    .A(_353_),
    .B(_380_),
    .Y(_381_)
);

NOR2X1 _2636_ (
    .A(_381_),
    .B(_339_),
    .Y(_382_)
);

AND2X2 _2637_ (
    .A(_382_),
    .B(_377_),
    .Y(_383_)
);

NOR2X1 _2638_ (
    .A(_377_),
    .B(_382_),
    .Y(_384_)
);

OAI21X1 _2639_ (
    .A(_384_),
    .B(_383_),
    .C(RDY_bF$buf6),
    .Y(_385_)
);

OAI21X1 _2640_ (
    .A(RDY_bF$buf5),
    .B(_123_),
    .C(_385_),
    .Y(_10_)
);

INVX1 _2641_ (
    .A(_377_),
    .Y(_386_)
);

AOI21X1 _2642_ (
    .A(_374_),
    .B(_375_),
    .C(_290_),
    .Y(_387_)
);

AOI22X1 _2643_ (
    .A(ADD[1]),
    .B(_1038_),
    .C(_306_),
    .D(ABH[1]),
    .Y(_388_)
);

NAND3X1 _2644_ (
    .A(_1074__bF$buf3),
    .B(_1395_),
    .C(_388_),
    .Y(_389_)
);

AOI21X1 _2645_ (
    .A(DIMUX[1]),
    .B(_314_),
    .C(_389_),
    .Y(_390_)
);

OAI21X1 _2646_ (
    .A(_134_),
    .B(_387_),
    .C(_390_),
    .Y(_391_)
);

INVX1 _2647_ (
    .A(_391_),
    .Y(_392_)
);

AOI21X1 _2648_ (
    .A(_382_),
    .B(_386_),
    .C(_392_),
    .Y(_393_)
);

NAND2X1 _2649_ (
    .A(_386_),
    .B(_382_),
    .Y(_394_)
);

NOR2X1 _2650_ (
    .A(_391_),
    .B(_394_),
    .Y(_395_)
);

OAI21X1 _2651_ (
    .A(_393_),
    .B(_395_),
    .C(RDY_bF$buf4),
    .Y(_396_)
);

OAI21X1 _2652_ (
    .A(RDY_bF$buf3),
    .B(_134_),
    .C(_396_),
    .Y(_11_)
);

NOR2X1 _2653_ (
    .A(_377_),
    .B(_392_),
    .Y(_397_)
);

NAND2X1 _2654_ (
    .A(_397_),
    .B(_382_),
    .Y(_398_)
);

INVX1 _2655_ (
    .A(_398_),
    .Y(_399_)
);

AOI21X1 _2656_ (
    .A(_298_),
    .B(_297_),
    .C(_838_),
    .Y(_400_)
);

OAI22X1 _2657_ (
    .A(_1403_),
    .B(_1162_),
    .C(_140_),
    .D(_301_),
    .Y(_401_)
);

NAND3X1 _2658_ (
    .A(ADD[2]),
    .B(_856__bF$buf2),
    .C(_1157_),
    .Y(_402_)
);

NAND3X1 _2659_ (
    .A(ABH[2]),
    .B(_874_),
    .C(_1343_),
    .Y(_403_)
);

NAND3X1 _2660_ (
    .A(_1074__bF$buf2),
    .B(_402_),
    .C(_403_),
    .Y(_404_)
);

NOR3X1 _2661_ (
    .A(_401_),
    .B(_404_),
    .C(_400_),
    .Y(_405_)
);

NAND3X1 _2662_ (
    .A(PC[10]),
    .B(_375_),
    .C(_374_),
    .Y(_406_)
);

AND2X2 _2663_ (
    .A(_405_),
    .B(_406_),
    .Y(_407_)
);

INVX1 _2664_ (
    .A(_407_),
    .Y(_408_)
);

NOR2X1 _2665_ (
    .A(_408_),
    .B(_399_),
    .Y(_409_)
);

OAI21X1 _2666_ (
    .A(_407_),
    .B(_398_),
    .C(RDY_bF$buf2),
    .Y(_410_)
);

OAI22X1 _2667_ (
    .A(RDY_bF$buf1),
    .B(_140_),
    .C(_410_),
    .D(_409_),
    .Y(_12_)
);

AOI22X1 _2668_ (
    .A(ADD[3]),
    .B(_1038_),
    .C(_306_),
    .D(ABH[3]),
    .Y(_411_)
);

NAND3X1 _2669_ (
    .A(_1074__bF$buf1),
    .B(_1413_),
    .C(_411_),
    .Y(_412_)
);

AOI21X1 _2670_ (
    .A(DIMUX[3]),
    .B(_314_),
    .C(_412_),
    .Y(_413_)
);

OAI21X1 _2671_ (
    .A(_146_),
    .B(_387_),
    .C(_413_),
    .Y(_414_)
);

INVX1 _2672_ (
    .A(_414_),
    .Y(_415_)
);

OAI21X1 _2673_ (
    .A(_407_),
    .B(_398_),
    .C(_415_),
    .Y(_416_)
);

NAND3X1 _2674_ (
    .A(_408_),
    .B(_414_),
    .C(_399_),
    .Y(_417_)
);

NAND3X1 _2675_ (
    .A(RDY_bF$buf0),
    .B(_416_),
    .C(_417_),
    .Y(_418_)
);

OAI21X1 _2676_ (
    .A(RDY_bF$buf8),
    .B(_146_),
    .C(_418_),
    .Y(_13_)
);

AOI22X1 _2677_ (
    .A(ADD[4]),
    .B(_1038_),
    .C(_306_),
    .D(ABH[4]),
    .Y(_419_)
);

NAND3X1 _2678_ (
    .A(_1074__bF$buf0),
    .B(_1421_),
    .C(_419_),
    .Y(_420_)
);

AOI21X1 _2679_ (
    .A(DIMUX[4]),
    .B(_314_),
    .C(_420_),
    .Y(_421_)
);

OAI21X1 _2680_ (
    .A(_152_),
    .B(_387_),
    .C(_421_),
    .Y(_422_)
);

NOR2X1 _2681_ (
    .A(_407_),
    .B(_415_),
    .Y(_423_)
);

NAND3X1 _2682_ (
    .A(_397_),
    .B(_423_),
    .C(_382_),
    .Y(_424_)
);

NOR2X1 _2683_ (
    .A(_422_),
    .B(_424_),
    .Y(_425_)
);

INVX1 _2684_ (
    .A(_422_),
    .Y(_426_)
);

AOI22X1 _2685_ (
    .A(_372_),
    .B(_376_),
    .C(_405_),
    .D(_406_),
    .Y(_427_)
);

NAND3X1 _2686_ (
    .A(_391_),
    .B(_414_),
    .C(_427_),
    .Y(_428_)
);

NOR3X1 _2687_ (
    .A(_428_),
    .B(_381_),
    .C(_339_),
    .Y(_429_)
);

NOR2X1 _2688_ (
    .A(_426_),
    .B(_429_),
    .Y(_430_)
);

OAI21X1 _2689_ (
    .A(_430_),
    .B(_425_),
    .C(RDY_bF$buf7),
    .Y(_431_)
);

OAI21X1 _2690_ (
    .A(RDY_bF$buf6),
    .B(_152_),
    .C(_431_),
    .Y(_14_)
);

AOI22X1 _2691_ (
    .A(ADD[5]),
    .B(_1038_),
    .C(_306_),
    .D(ABH[5]),
    .Y(_432_)
);

NAND3X1 _2692_ (
    .A(_1074__bF$buf3),
    .B(_1429_),
    .C(_432_),
    .Y(_433_)
);

AOI21X1 _2693_ (
    .A(DIMUX[5]),
    .B(_314_),
    .C(_433_),
    .Y(_434_)
);

OAI21X1 _2694_ (
    .A(_271_),
    .B(_387_),
    .C(_434_),
    .Y(_435_)
);

OAI21X1 _2695_ (
    .A(_426_),
    .B(_424_),
    .C(_435_),
    .Y(_436_)
);

INVX1 _2696_ (
    .A(_435_),
    .Y(_437_)
);

NAND3X1 _2697_ (
    .A(_422_),
    .B(_437_),
    .C(_429_),
    .Y(_438_)
);

NAND3X1 _2698_ (
    .A(RDY_bF$buf5),
    .B(_438_),
    .C(_436_),
    .Y(_439_)
);

NAND2X1 _2699_ (
    .A(_836__bF$buf3),
    .B(_271_),
    .Y(_440_)
);

AND2X2 _2700_ (
    .A(_439_),
    .B(_440_),
    .Y(_15_)
);

NAND2X1 _2701_ (
    .A(PC[14]),
    .B(_836__bF$buf2),
    .Y(_441_)
);

AOI22X1 _2702_ (
    .A(ADD[6]),
    .B(_1038_),
    .C(_306_),
    .D(ABH[6]),
    .Y(_442_)
);

NAND3X1 _2703_ (
    .A(_1074__bF$buf2),
    .B(_442_),
    .C(_1439_),
    .Y(_443_)
);

AOI21X1 _2704_ (
    .A(DIMUX[6]),
    .B(_314_),
    .C(_443_),
    .Y(_444_)
);

OAI21X1 _2705_ (
    .A(_161_),
    .B(_387_),
    .C(_444_),
    .Y(_445_)
);

NOR2X1 _2706_ (
    .A(_426_),
    .B(_437_),
    .Y(_446_)
);

NAND2X1 _2707_ (
    .A(_446_),
    .B(_429_),
    .Y(_447_)
);

XOR2X1 _2708_ (
    .A(_447_),
    .B(_445_),
    .Y(_448_)
);

OAI21X1 _2709_ (
    .A(_836__bF$buf1),
    .B(_448_),
    .C(_441_),
    .Y(_16_)
);

NAND2X1 _2710_ (
    .A(PC[15]),
    .B(_836__bF$buf0),
    .Y(_449_)
);

AOI22X1 _2711_ (
    .A(\ALU.N ),
    .B(_1038_),
    .C(_306_),
    .D(ABH[7]),
    .Y(_450_)
);

NAND3X1 _2712_ (
    .A(_1074__bF$buf1),
    .B(_450_),
    .C(_1449_),
    .Y(_451_)
);

AOI21X1 _2713_ (
    .A(DIMUX[7]),
    .B(_314_),
    .C(_451_),
    .Y(_452_)
);

OAI21X1 _2714_ (
    .A(_167_),
    .B(_387_),
    .C(_452_),
    .Y(_453_)
);

NAND3X1 _2715_ (
    .A(_446_),
    .B(_445_),
    .C(_429_),
    .Y(_454_)
);

XOR2X1 _2716_ (
    .A(_454_),
    .B(_453_),
    .Y(_455_)
);

OAI21X1 _2717_ (
    .A(_836__bF$buf7),
    .B(_455_),
    .C(_449_),
    .Y(_17_)
);

INVX1 _2718_ (
    .A(NMI_1),
    .Y(_456_)
);

NAND3X1 _2719_ (
    .A(NMI),
    .B(_456_),
    .C(_866_),
    .Y(_457_)
);

OAI21X1 _2720_ (
    .A(_866_),
    .B(_1076_),
    .C(_457_),
    .Y(_18_)
);

INVX1 _2721_ (
    .A(cond_code[0]),
    .Y(_458_)
);

INVX2 _2722_ (
    .A(_886_),
    .Y(_459_)
);

NAND2X1 _2723_ (
    .A(RDY_bF$buf4),
    .B(_459_),
    .Y(_460_)
);

OAI21X1 _2724_ (
    .A(RDY_bF$buf3),
    .B(_458_),
    .C(_460_),
    .Y(_19_)
);

NAND2X1 _2725_ (
    .A(cond_code[1]),
    .B(_836__bF$buf6),
    .Y(_461_)
);

OAI21X1 _2726_ (
    .A(_836__bF$buf5),
    .B(_1091_),
    .C(_461_),
    .Y(_20_)
);

NAND2X1 _2727_ (
    .A(cond_code[2]),
    .B(_836__bF$buf4),
    .Y(_462_)
);

OAI21X1 _2728_ (
    .A(_836__bF$buf3),
    .B(_890_),
    .C(_462_),
    .Y(_21_)
);

INVX2 _2729_ (
    .A(plp),
    .Y(_463_)
);

OAI22X1 _2730_ (
    .A(_463_),
    .B(_860__bF$buf1),
    .C(_893_),
    .D(_1105_),
    .Y(_22_)
);

INVX1 _2731_ (
    .A(_983_),
    .Y(_464_)
);

NOR2X1 _2732_ (
    .A(_861__bF$buf0),
    .B(_464_),
    .Y(_465_)
);

NAND2X1 _2733_ (
    .A(_1191_),
    .B(_465_),
    .Y(_466_)
);

OAI21X1 _2734_ (
    .A(_127_),
    .B(_860__bF$buf0),
    .C(_466_),
    .Y(_23_)
);

OAI21X1 _2735_ (
    .A(_836__bF$buf2),
    .B(_859__bF$buf0),
    .C(clc),
    .Y(_467_)
);

NAND2X1 _2736_ (
    .A(_886_),
    .B(_1143_),
    .Y(_468_)
);

OR2X2 _2737_ (
    .A(_464_),
    .B(_1190_),
    .Y(_469_)
);

OAI21X1 _2738_ (
    .A(_468_),
    .B(_469_),
    .C(_467_),
    .Y(_24_)
);

INVX1 _2739_ (
    .A(sec),
    .Y(_470_)
);

NOR2X1 _2740_ (
    .A(_859__bF$buf3),
    .B(_460_),
    .Y(_471_)
);

NAND2X1 _2741_ (
    .A(_965_),
    .B(_471_),
    .Y(_472_)
);

OAI22X1 _2742_ (
    .A(_470_),
    .B(_860__bF$buf4),
    .C(_472_),
    .D(_469_),
    .Y(_25_)
);

OAI21X1 _2743_ (
    .A(_836__bF$buf1),
    .B(_859__bF$buf2),
    .C(cld),
    .Y(_473_)
);

NOR2X1 _2744_ (
    .A(_890_),
    .B(_1091_),
    .Y(_474_)
);

NAND2X1 _2745_ (
    .A(_474_),
    .B(_983_),
    .Y(_475_)
);

OAI21X1 _2746_ (
    .A(_468_),
    .B(_475_),
    .C(_473_),
    .Y(_26_)
);

INVX1 _2747_ (
    .A(sed),
    .Y(_476_)
);

OAI22X1 _2748_ (
    .A(_476_),
    .B(_860__bF$buf3),
    .C(_475_),
    .D(_472_),
    .Y(_27_)
);

OAI21X1 _2749_ (
    .A(_836__bF$buf0),
    .B(_859__bF$buf1),
    .C(cli),
    .Y(_477_)
);

NAND2X1 _2750_ (
    .A(_1098_),
    .B(_983_),
    .Y(_478_)
);

OAI21X1 _2751_ (
    .A(_468_),
    .B(_478_),
    .C(_477_),
    .Y(_28_)
);

INVX1 _2752_ (
    .A(sei),
    .Y(_479_)
);

OAI22X1 _2753_ (
    .A(_479_),
    .B(_860__bF$buf2),
    .C(_478_),
    .D(_472_),
    .Y(_29_)
);

INVX1 _2754_ (
    .A(clv),
    .Y(_480_)
);

NOR2X1 _2755_ (
    .A(_890_),
    .B(_893_),
    .Y(_481_)
);

NAND2X1 _2756_ (
    .A(_459_),
    .B(_481_),
    .Y(_482_)
);

NOR2X1 _2757_ (
    .A(_883_),
    .B(_482_),
    .Y(_483_)
);

NAND2X1 _2758_ (
    .A(_483_),
    .B(_465_),
    .Y(_484_)
);

OAI21X1 _2759_ (
    .A(_480_),
    .B(_860__bF$buf1),
    .C(_484_),
    .Y(_30_)
);

NOR2X1 _2760_ (
    .A(_886_),
    .B(_893_),
    .Y(_485_)
);

NAND3X1 _2761_ (
    .A(_1119_),
    .B(_1186_),
    .C(_485_),
    .Y(_486_)
);

OR2X2 _2762_ (
    .A(_486_),
    .B(_1092_),
    .Y(_487_)
);

OAI21X1 _2763_ (
    .A(_836__bF$buf7),
    .B(_859__bF$buf0),
    .C(bit_ins),
    .Y(_488_)
);

OAI21X1 _2764_ (
    .A(_861__bF$buf3),
    .B(_487_),
    .C(_488_),
    .Y(_31_)
);

NOR2X1 _2765_ (
    .A(_974_),
    .B(_1178_),
    .Y(_489_)
);

NOR2X1 _2766_ (
    .A(_974_),
    .B(_971_),
    .Y(_490_)
);

OAI21X1 _2767_ (
    .A(_886_),
    .B(_1091_),
    .C(_490_),
    .Y(_491_)
);

OAI21X1 _2768_ (
    .A(_886_),
    .B(_491_),
    .C(_487_),
    .Y(_492_)
);

NOR2X1 _2769_ (
    .A(_489_),
    .B(_492_),
    .Y(_493_)
);

OAI21X1 _2770_ (
    .A(_1092_),
    .B(_486_),
    .C(_491_),
    .Y(_494_)
);

OAI21X1 _2771_ (
    .A(_489_),
    .B(_494_),
    .C(_860__bF$buf0),
    .Y(_495_)
);

INVX1 _2772_ (
    .A(_495_),
    .Y(_496_)
);

AOI22X1 _2773_ (
    .A(_1452_),
    .B(_861__bF$buf2),
    .C(_493_),
    .D(_496_),
    .Y(_32_)
);

NOR2X1 _2774_ (
    .A(_489_),
    .B(_494_),
    .Y(_497_)
);

INVX1 _2775_ (
    .A(_474_),
    .Y(_498_)
);

INVX1 _2776_ (
    .A(_1179_),
    .Y(_499_)
);

NAND2X1 _2777_ (
    .A(_474_),
    .B(_982_),
    .Y(_500_)
);

OR2X2 _2778_ (
    .A(_499_),
    .B(_500_),
    .Y(_501_)
);

NOR2X1 _2779_ (
    .A(_872_),
    .B(_1178_),
    .Y(_502_)
);

AOI21X1 _2780_ (
    .A(_502_),
    .B(_886_),
    .C(_972_),
    .Y(_503_)
);

OAI21X1 _2781_ (
    .A(_498_),
    .B(_503_),
    .C(_501_),
    .Y(_504_)
);

NAND2X1 _2782_ (
    .A(_883_),
    .B(_474_),
    .Y(_505_)
);

NAND3X1 _2783_ (
    .A(_1187_),
    .B(_883_),
    .C(_1186_),
    .Y(_506_)
);

OAI22X1 _2784_ (
    .A(_498_),
    .B(_506_),
    .C(_505_),
    .D(_1189_),
    .Y(_507_)
);

INVX1 _2785_ (
    .A(_507_),
    .Y(_508_)
);

NAND2X1 _2786_ (
    .A(_481_),
    .B(_982_),
    .Y(_509_)
);

OAI21X1 _2787_ (
    .A(_464_),
    .B(_509_),
    .C(_508_),
    .Y(_510_)
);

NOR2X1 _2788_ (
    .A(_510_),
    .B(_504_),
    .Y(_511_)
);

INVX1 _2789_ (
    .A(_1178_),
    .Y(_512_)
);

NAND2X1 _2790_ (
    .A(_886_),
    .B(_893_),
    .Y(_513_)
);

NOR2X1 _2791_ (
    .A(_971_),
    .B(_513_),
    .Y(_514_)
);

OAI21X1 _2792_ (
    .A(_512_),
    .B(_514_),
    .C(_890_),
    .Y(_515_)
);

NAND2X1 _2793_ (
    .A(_515_),
    .B(_511_),
    .Y(_516_)
);

OAI21X1 _2794_ (
    .A(_497_),
    .B(_516_),
    .C(_860__bF$buf4),
    .Y(_517_)
);

OAI21X1 _2795_ (
    .A(_1456_),
    .B(_860__bF$buf3),
    .C(_517_),
    .Y(_33_)
);

INVX1 _2796_ (
    .A(op[2]),
    .Y(_518_)
);

OAI21X1 _2797_ (
    .A(_1178_),
    .B(_894_),
    .C(_860__bF$buf2),
    .Y(_519_)
);

NOR2X1 _2798_ (
    .A(_519_),
    .B(_494_),
    .Y(_520_)
);

AOI22X1 _2799_ (
    .A(_518_),
    .B(_861__bF$buf1),
    .C(_511_),
    .D(_520_),
    .Y(_34_)
);

OAI21X1 _2800_ (
    .A(_117_),
    .B(_860__bF$buf1),
    .C(_495_),
    .Y(_35_)
);

INVX1 _2801_ (
    .A(_489_),
    .Y(_521_)
);

OAI21X1 _2802_ (
    .A(_967_),
    .B(_1119_),
    .C(_471_),
    .Y(_522_)
);

OAI22X1 _2803_ (
    .A(_1293_),
    .B(_860__bF$buf0),
    .C(_521_),
    .D(_522_),
    .Y(_36_)
);

OAI21X1 _2804_ (
    .A(_836__bF$buf6),
    .B(_859__bF$buf3),
    .C(_288_),
    .Y(_523_)
);

AND2X2 _2805_ (
    .A(_519_),
    .B(_523_),
    .Y(_37_)
);

NOR2X1 _2806_ (
    .A(_890_),
    .B(_861__bF$buf0),
    .Y(_524_)
);

AOI22X1 _2807_ (
    .A(compare),
    .B(_861__bF$buf3),
    .C(_514_),
    .D(_524_),
    .Y(_525_)
);

OAI21X1 _2808_ (
    .A(_861__bF$buf2),
    .B(_508_),
    .C(_525_),
    .Y(_38_)
);

NAND2X1 _2809_ (
    .A(_860__bF$buf4),
    .B(_489_),
    .Y(_526_)
);

OAI22X1 _2810_ (
    .A(_1295_),
    .B(_860__bF$buf3),
    .C(_1109_),
    .D(_526_),
    .Y(_39_)
);

OAI21X1 _2811_ (
    .A(_1343_),
    .B(_1001_),
    .C(RDY_bF$buf2),
    .Y(_527_)
);

NAND2X1 _2812_ (
    .A(adc_bcd),
    .B(_527_),
    .Y(_528_)
);

NOR2X1 _2813_ (
    .A(_886_),
    .B(_1091_),
    .Y(_529_)
);

INVX1 _2814_ (
    .A(_527_),
    .Y(_530_)
);

NAND3X1 _2815_ (
    .A(_529_),
    .B(_530_),
    .C(_972_),
    .Y(_531_)
);

NAND2X1 _2816_ (
    .A(D),
    .B(_890_),
    .Y(_532_)
);

OAI21X1 _2817_ (
    .A(_532_),
    .B(_531_),
    .C(_528_),
    .Y(_40_)
);

INVX1 _2818_ (
    .A(adc_sbc),
    .Y(_533_)
);

OAI21X1 _2819_ (
    .A(_533_),
    .B(_530_),
    .C(_531_),
    .Y(_41_)
);

INVX1 _2820_ (
    .A(_505_),
    .Y(_534_)
);

AOI22X1 _2821_ (
    .A(inc),
    .B(_861__bF$buf1),
    .C(_465_),
    .D(_534_),
    .Y(_535_)
);

NAND3X1 _2822_ (
    .A(_459_),
    .B(_474_),
    .C(_502_),
    .Y(_536_)
);

OAI21X1 _2823_ (
    .A(_861__bF$buf0),
    .B(_536_),
    .C(_535_),
    .Y(_42_)
);

OAI21X1 _2824_ (
    .A(_836__bF$buf5),
    .B(_859__bF$buf2),
    .C(load_only),
    .Y(_537_)
);

OAI21X1 _2825_ (
    .A(_861__bF$buf3),
    .B(_482_),
    .C(_537_),
    .Y(_43_)
);

INVX1 _2826_ (
    .A(_481_),
    .Y(_538_)
);

NAND3X1 _2827_ (
    .A(_860__bF$buf2),
    .B(_538_),
    .C(_502_),
    .Y(_539_)
);

OAI21X1 _2828_ (
    .A(_1064_),
    .B(_860__bF$buf1),
    .C(_539_),
    .Y(_44_)
);

INVX1 _2829_ (
    .A(_524_),
    .Y(_540_)
);

OAI21X1 _2830_ (
    .A(_836__bF$buf4),
    .B(_859__bF$buf1),
    .C(store),
    .Y(_541_)
);

OAI21X1 _2831_ (
    .A(_885_),
    .B(_892_),
    .C(_868_),
    .Y(_542_)
);

NOR2X1 _2832_ (
    .A(_970_),
    .B(_872_),
    .Y(_543_)
);

OAI21X1 _2833_ (
    .A(_543_),
    .B(_972_),
    .C(_542_),
    .Y(_544_)
);

OAI21X1 _2834_ (
    .A(_540_),
    .B(_544_),
    .C(_541_),
    .Y(_45_)
);

NOR2X1 _2835_ (
    .A(_883_),
    .B(_538_),
    .Y(_545_)
);

OAI21X1 _2836_ (
    .A(_883_),
    .B(_1110_),
    .C(_973_),
    .Y(_546_)
);

AOI21X1 _2837_ (
    .A(_545_),
    .B(_502_),
    .C(_546_),
    .Y(_547_)
);

OAI21X1 _2838_ (
    .A(_836__bF$buf3),
    .B(_859__bF$buf0),
    .C(index_y),
    .Y(_548_)
);

OAI21X1 _2839_ (
    .A(_861__bF$buf2),
    .B(_547_),
    .C(_548_),
    .Y(_46_)
);

NAND2X1 _2840_ (
    .A(_886_),
    .B(_974_),
    .Y(_549_)
);

NAND2X1 _2841_ (
    .A(_1091_),
    .B(_1119_),
    .Y(_550_)
);

OAI21X1 _2842_ (
    .A(_549_),
    .B(_550_),
    .C(_500_),
    .Y(_551_)
);

NAND2X1 _2843_ (
    .A(_1186_),
    .B(_551_),
    .Y(_552_)
);

NOR2X1 _2844_ (
    .A(_890_),
    .B(_887_),
    .Y(_553_)
);

AND2X2 _2845_ (
    .A(_545_),
    .B(_886_),
    .Y(_554_)
);

OAI21X1 _2846_ (
    .A(_553_),
    .B(_554_),
    .C(_983_),
    .Y(_555_)
);

NAND2X1 _2847_ (
    .A(_552_),
    .B(_555_),
    .Y(_556_)
);

NAND2X1 _2848_ (
    .A(_1179_),
    .B(_483_),
    .Y(_557_)
);

INVX1 _2849_ (
    .A(_557_),
    .Y(_558_)
);

OAI21X1 _2850_ (
    .A(_558_),
    .B(_556_),
    .C(_860__bF$buf0),
    .Y(_559_)
);

OAI21X1 _2851_ (
    .A(_1359_),
    .B(_860__bF$buf4),
    .C(_559_),
    .Y(_47_)
);

NAND2X1 _2852_ (
    .A(_474_),
    .B(_1099_),
    .Y(_560_)
);

NOR2X1 _2853_ (
    .A(_879_),
    .B(_560_),
    .Y(_561_)
);

INVX1 _2854_ (
    .A(_561_),
    .Y(_562_)
);

NOR2X1 _2855_ (
    .A(_459_),
    .B(_1109_),
    .Y(_563_)
);

NAND3X1 _2856_ (
    .A(_512_),
    .B(_481_),
    .C(_563_),
    .Y(_564_)
);

NAND3X1 _2857_ (
    .A(_562_),
    .B(_564_),
    .C(_501_),
    .Y(_565_)
);

OAI21X1 _2858_ (
    .A(_565_),
    .B(_556_),
    .C(_860__bF$buf3),
    .Y(_566_)
);

OAI21X1 _2859_ (
    .A(_1333_),
    .B(_860__bF$buf2),
    .C(_566_),
    .Y(_48_)
);

INVX1 _2860_ (
    .A(dst_reg[0]),
    .Y(_567_)
);

NAND2X1 _2861_ (
    .A(_883_),
    .B(_983_),
    .Y(_568_)
);

OAI21X1 _2862_ (
    .A(_1119_),
    .B(_883_),
    .C(_1186_),
    .Y(_569_)
);

OAI22X1 _2863_ (
    .A(_482_),
    .B(_569_),
    .C(_549_),
    .D(_568_),
    .Y(_570_)
);

NAND2X1 _2864_ (
    .A(_886_),
    .B(_545_),
    .Y(_571_)
);

OAI21X1 _2865_ (
    .A(_499_),
    .B(_571_),
    .C(_984_),
    .Y(_572_)
);

OAI21X1 _2866_ (
    .A(_572_),
    .B(_570_),
    .C(_860__bF$buf1),
    .Y(_573_)
);

OAI21X1 _2867_ (
    .A(_567_),
    .B(_860__bF$buf0),
    .C(_573_),
    .Y(_49_)
);

INVX1 _2868_ (
    .A(_570_),
    .Y(_574_)
);

INVX1 _2869_ (
    .A(_482_),
    .Y(_575_)
);

AOI22X1 _2870_ (
    .A(_512_),
    .B(_575_),
    .C(_561_),
    .D(_969_),
    .Y(_576_)
);

NAND3X1 _2871_ (
    .A(_501_),
    .B(_576_),
    .C(_574_),
    .Y(_577_)
);

INVX1 _2872_ (
    .A(_577_),
    .Y(_578_)
);

OAI21X1 _2873_ (
    .A(_836__bF$buf2),
    .B(_859__bF$buf3),
    .C(dst_reg[1]),
    .Y(_579_)
);

OAI21X1 _2874_ (
    .A(_861__bF$buf1),
    .B(_578_),
    .C(_579_),
    .Y(_50_)
);

INVX1 _2875_ (
    .A(load_reg),
    .Y(_580_)
);

NAND2X1 _2876_ (
    .A(_543_),
    .B(_483_),
    .Y(_581_)
);

OAI21X1 _2877_ (
    .A(_459_),
    .B(_890_),
    .C(_972_),
    .Y(_582_)
);

NOR2X1 _2878_ (
    .A(_970_),
    .B(_459_),
    .Y(_583_)
);

NAND3X1 _2879_ (
    .A(_969_),
    .B(_481_),
    .C(_583_),
    .Y(_584_)
);

NAND3X1 _2880_ (
    .A(_582_),
    .B(_584_),
    .C(_581_),
    .Y(_585_)
);

OAI21X1 _2881_ (
    .A(_1092_),
    .B(_499_),
    .C(_568_),
    .Y(_586_)
);

NOR2X1 _2882_ (
    .A(_970_),
    .B(_965_),
    .Y(_587_)
);

NAND2X1 _2883_ (
    .A(_587_),
    .B(_575_),
    .Y(_588_)
);

NAND3X1 _2884_ (
    .A(_588_),
    .B(_557_),
    .C(_501_),
    .Y(_589_)
);

OR2X2 _2885_ (
    .A(_589_),
    .B(_586_),
    .Y(_590_)
);

OAI21X1 _2886_ (
    .A(_585_),
    .B(_590_),
    .C(_860__bF$buf4),
    .Y(_591_)
);

OAI21X1 _2887_ (
    .A(_580_),
    .B(_860__bF$buf3),
    .C(_591_),
    .Y(_51_)
);

NOR2X1 _2888_ (
    .A(_316_),
    .B(_1343_),
    .Y(_52_)
);

OAI21X1 _2889_ (
    .A(_980_),
    .B(_1058_),
    .C(RDY_bF$buf1),
    .Y(_592_)
);

NOR2X1 _2890_ (
    .A(reset),
    .B(_592_),
    .Y(_593_)
);

INVX2 _2891_ (
    .A(_593_),
    .Y(_594_)
);

OAI21X1 _2892_ (
    .A(reset),
    .B(_592_),
    .C(IRHOLD[0]),
    .Y(_595_)
);

OAI21X1 _2893_ (
    .A(_1304_),
    .B(_594_),
    .C(_595_),
    .Y(_53_)
);

OAI21X1 _2894_ (
    .A(reset),
    .B(_592_),
    .C(IRHOLD[1]),
    .Y(_596_)
);

OAI21X1 _2895_ (
    .A(_1324_),
    .B(_594_),
    .C(_596_),
    .Y(_54_)
);

OAI21X1 _2896_ (
    .A(reset),
    .B(_592_),
    .C(IRHOLD[2]),
    .Y(_597_)
);

OAI21X1 _2897_ (
    .A(_838_),
    .B(_594_),
    .C(_597_),
    .Y(_55_)
);

OAI21X1 _2898_ (
    .A(reset),
    .B(_592_),
    .C(IRHOLD[3]),
    .Y(_598_)
);

OAI21X1 _2899_ (
    .A(_1327_),
    .B(_594_),
    .C(_598_),
    .Y(_56_)
);

OAI21X1 _2900_ (
    .A(reset),
    .B(_592_),
    .C(IRHOLD[4]),
    .Y(_599_)
);

OAI21X1 _2901_ (
    .A(_1329_),
    .B(_594_),
    .C(_599_),
    .Y(_57_)
);

OAI21X1 _2902_ (
    .A(reset),
    .B(_592_),
    .C(IRHOLD[5]),
    .Y(_600_)
);

OAI21X1 _2903_ (
    .A(_844_),
    .B(_594_),
    .C(_600_),
    .Y(_58_)
);

OAI21X1 _2904_ (
    .A(reset),
    .B(_592_),
    .C(IRHOLD[6]),
    .Y(_601_)
);

OAI21X1 _2905_ (
    .A(_846_),
    .B(_594_),
    .C(_601_),
    .Y(_59_)
);

OAI21X1 _2906_ (
    .A(reset),
    .B(_592_),
    .C(IRHOLD[7]),
    .Y(_602_)
);

OAI21X1 _2907_ (
    .A(_847_),
    .B(_594_),
    .C(_602_),
    .Y(_60_)
);

OAI21X1 _2908_ (
    .A(_863_),
    .B(_860__bF$buf2),
    .C(_592_),
    .Y(_61_)
);

OAI21X1 _2909_ (
    .A(_917__bF$buf2),
    .B(_1035_),
    .C(_859__bF$buf2),
    .Y(_603_)
);

AOI21X1 _2910_ (
    .A(_955_),
    .B(bit_ins),
    .C(_603_),
    .Y(_604_)
);

NOR2X1 _2911_ (
    .A(plp),
    .B(_859__bF$buf1),
    .Y(_605_)
);

NOR2X1 _2912_ (
    .A(adc_sbc),
    .B(clv),
    .Y(_606_)
);

AOI21X1 _2913_ (
    .A(_605_),
    .B(_606_),
    .C(_604_),
    .Y(_607_)
);

INVX1 _2914_ (
    .A(ADD[6]),
    .Y(_608_)
);

NAND3X1 _2915_ (
    .A(\ALU.V ),
    .B(_463_),
    .C(_480_),
    .Y(_609_)
);

OAI21X1 _2916_ (
    .A(_463_),
    .B(_608_),
    .C(_609_),
    .Y(_610_)
);

NAND2X1 _2917_ (
    .A(_610_),
    .B(_1343_),
    .Y(_611_)
);

OAI21X1 _2918_ (
    .A(_846_),
    .B(_1343_),
    .C(_611_),
    .Y(_612_)
);

NAND2X1 _2919_ (
    .A(_612_),
    .B(_607_),
    .Y(_613_)
);

OAI21X1 _2920_ (
    .A(_1127_),
    .B(_607_),
    .C(_613_),
    .Y(_62_)
);

NOR2X1 _2921_ (
    .A(cld),
    .B(plp),
    .Y(_614_)
);

NAND2X1 _2922_ (
    .A(_476_),
    .B(_614_),
    .Y(_615_)
);

OAI21X1 _2923_ (
    .A(_859__bF$buf0),
    .B(_615_),
    .C(_603_),
    .Y(_616_)
);

NAND2X1 _2924_ (
    .A(D),
    .B(_616_),
    .Y(_617_)
);

INVX1 _2925_ (
    .A(ADD[3]),
    .Y(_618_)
);

INVX1 _2926_ (
    .A(_614_),
    .Y(_619_)
);

OAI21X1 _2927_ (
    .A(_463_),
    .B(_618_),
    .C(_619_),
    .Y(_620_)
);

MUX2X1 _2928_ (
    .A(_620_),
    .B(DIMUX[3]),
    .S(_1381_),
    .Y(_621_)
);

OAI21X1 _2929_ (
    .A(_616_),
    .B(_621_),
    .C(_617_),
    .Y(_63_)
);

NOR2X1 _2930_ (
    .A(cli),
    .B(_1205_),
    .Y(_622_)
);

NAND2X1 _2931_ (
    .A(_479_),
    .B(_622_),
    .Y(_623_)
);

INVX1 _2932_ (
    .A(_603_),
    .Y(_624_)
);

AOI21X1 _2933_ (
    .A(_624_),
    .B(_1075_),
    .C(_605_),
    .Y(_625_)
);

OAI21X1 _2934_ (
    .A(_1204_),
    .B(_625_),
    .C(_623_),
    .Y(_626_)
);

INVX1 _2935_ (
    .A(ADD[2]),
    .Y(_627_)
);

NOR2X1 _2936_ (
    .A(_627_),
    .B(_1204_),
    .Y(_628_)
);

OAI21X1 _2937_ (
    .A(_628_),
    .B(_622_),
    .C(_1381_),
    .Y(_629_)
);

OAI21X1 _2938_ (
    .A(_838_),
    .B(_1381_),
    .C(_629_),
    .Y(_630_)
);

NOR2X1 _2939_ (
    .A(_1076_),
    .B(_630_),
    .Y(_631_)
);

NAND2X1 _2940_ (
    .A(I),
    .B(_626_),
    .Y(_632_)
);

OAI21X1 _2941_ (
    .A(_626_),
    .B(_631_),
    .C(_632_),
    .Y(_64_)
);

OAI21X1 _2942_ (
    .A(_1350_),
    .B(_1356_),
    .C(load_reg),
    .Y(_633_)
);

INVX1 _2943_ (
    .A(_605_),
    .Y(_634_)
);

NOR2X1 _2944_ (
    .A(compare),
    .B(_634_),
    .Y(_635_)
);

AOI22X1 _2945_ (
    .A(_935_),
    .B(_604_),
    .C(_633_),
    .D(_635_),
    .Y(_636_)
);

NOR2X1 _2946_ (
    .A(N),
    .B(_636_),
    .Y(_637_)
);

OAI21X1 _2947_ (
    .A(_463_),
    .B(\ALU.N ),
    .C(_1343_),
    .Y(_638_)
);

OAI21X1 _2948_ (
    .A(_847_),
    .B(_1343_),
    .C(_638_),
    .Y(_639_)
);

INVX1 _2949_ (
    .A(\ALU.N ),
    .Y(_640_)
);

OAI21X1 _2950_ (
    .A(_605_),
    .B(_934_),
    .C(_640_),
    .Y(_641_)
);

OAI21X1 _2951_ (
    .A(_934_),
    .B(_639_),
    .C(_641_),
    .Y(_642_)
);

AOI21X1 _2952_ (
    .A(_636_),
    .B(_642_),
    .C(_637_),
    .Y(_65_)
);

INVX1 _2953_ (
    .A(Z),
    .Y(_643_)
);

INVX1 _2954_ (
    .A(bit_ins),
    .Y(_644_)
);

AND2X2 _2955_ (
    .A(_633_),
    .B(_635_),
    .Y(_645_)
);

AOI22X1 _2956_ (
    .A(_935_),
    .B(_624_),
    .C(_645_),
    .D(_644_),
    .Y(_646_)
);

OAI21X1 _2957_ (
    .A(_917__bF$buf1),
    .B(_933_),
    .C(_624_),
    .Y(_647_)
);

NAND2X1 _2958_ (
    .A(_644_),
    .B(_645_),
    .Y(_648_)
);

INVX1 _2959_ (
    .A(\ALU.Z ),
    .Y(_649_)
);

MUX2X1 _2960_ (
    .A(ADD[1]),
    .B(\ALU.Z ),
    .S(plp),
    .Y(_650_)
);

AOI21X1 _2961_ (
    .A(_1381_),
    .B(_650_),
    .C(_934_),
    .Y(_651_)
);

OAI21X1 _2962_ (
    .A(DIMUX[1]),
    .B(_1381_),
    .C(_651_),
    .Y(_652_)
);

OAI21X1 _2963_ (
    .A(_649_),
    .B(_935_),
    .C(_652_),
    .Y(_653_)
);

NAND3X1 _2964_ (
    .A(_647_),
    .B(_653_),
    .C(_648_),
    .Y(_654_)
);

OAI21X1 _2965_ (
    .A(_643_),
    .B(_646_),
    .C(_654_),
    .Y(_66_)
);

NOR2X1 _2966_ (
    .A(write_back),
    .B(_859__bF$buf3),
    .Y(_655_)
);

NAND3X1 _2967_ (
    .A(_1295_),
    .B(_533_),
    .C(_1297_),
    .Y(_656_)
);

NOR2X1 _2968_ (
    .A(plp),
    .B(clc),
    .Y(_657_)
);

NAND2X1 _2969_ (
    .A(_470_),
    .B(_657_),
    .Y(_658_)
);

OR2X2 _2970_ (
    .A(_658_),
    .B(_656_),
    .Y(_659_)
);

OAI21X1 _2971_ (
    .A(_1295_),
    .B(_935_),
    .C(_1381_),
    .Y(_660_)
);

AOI21X1 _2972_ (
    .A(_655_),
    .B(_659_),
    .C(_660_),
    .Y(_661_)
);

NAND2X1 _2973_ (
    .A(C),
    .B(_661_),
    .Y(_662_)
);

AOI21X1 _2974_ (
    .A(plp),
    .B(ADD[0]),
    .C(_657_),
    .Y(_663_)
);

NAND2X1 _2975_ (
    .A(\ALU.CO ),
    .B(_656_),
    .Y(_664_)
);

OAI21X1 _2976_ (
    .A(_656_),
    .B(_663_),
    .C(_664_),
    .Y(_665_)
);

MUX2X1 _2977_ (
    .A(_665_),
    .B(DIMUX[0]),
    .S(_1381_),
    .Y(_666_)
);

OAI21X1 _2978_ (
    .A(_661_),
    .B(_666_),
    .C(_662_),
    .Y(_67_)
);

INVX1 _2979_ (
    .A(backwards),
    .Y(_667_)
);

NAND2X1 _2980_ (
    .A(RDY_bF$buf0),
    .B(DI[7]),
    .Y(_668_)
);

OAI21X1 _2981_ (
    .A(RDY_bF$buf8),
    .B(_667_),
    .C(_668_),
    .Y(_68_)
);

NAND2X1 _2982_ (
    .A(_1351_),
    .B(_1356_),
    .Y(_669_)
);

OAI21X1 _2983_ (
    .A(_923__bF$buf3),
    .B(_1082_),
    .C(_1232_),
    .Y(_670_)
);

OAI21X1 _2984_ (
    .A(_957_),
    .B(_899__bF$buf4),
    .C(_1080_),
    .Y(_671_)
);

OR2X2 _2985_ (
    .A(_671_),
    .B(_670_),
    .Y(_672_)
);

OAI21X1 _2986_ (
    .A(_580_),
    .B(_634_),
    .C(_176_),
    .Y(_673_)
);

OAI21X1 _2987_ (
    .A(_673_),
    .B(_672_),
    .C(RDY_bF$buf7),
    .Y(_674_)
);

NOR2X1 _2988_ (
    .A(_674_),
    .B(_669_),
    .Y(_675_)
);

OAI21X1 _2989_ (
    .A(_899__bF$buf3),
    .B(_1313_),
    .C(ADD[0]),
    .Y(_676_)
);

OAI21X1 _2990_ (
    .A(_1304_),
    .B(_1080_),
    .C(_676_),
    .Y(_677_)
);

INVX1 _2991_ (
    .A(_677_),
    .Y(_678_)
);

NOR2X1 _2992_ (
    .A(\AXYS[0] [0]),
    .B(_675_),
    .Y(_679_)
);

AOI21X1 _2993_ (
    .A(_675_),
    .B(_678_),
    .C(_679_),
    .Y(_69_)
);

NOR2X1 _2994_ (
    .A(\AXYS[0] [1]),
    .B(_675_),
    .Y(_680_)
);

NAND3X1 _2995_ (
    .A(adj_bcd),
    .B(adc_bcd),
    .C(\ALU.HC ),
    .Y(_681_)
);

NOR2X1 _2996_ (
    .A(adc_bcd),
    .B(\ALU.HC ),
    .Y(_682_)
);

NAND2X1 _2997_ (
    .A(adj_bcd),
    .B(_682_),
    .Y(_683_)
);

NAND2X1 _2998_ (
    .A(_681_),
    .B(_683_),
    .Y(_684_)
);

NAND2X1 _2999_ (
    .A(ADD[1]),
    .B(_684_),
    .Y(_685_)
);

INVX1 _3000_ (
    .A(_685_),
    .Y(_686_)
);

NOR2X1 _3001_ (
    .A(_1081_),
    .B(_686_),
    .Y(_687_)
);

OAI21X1 _3002_ (
    .A(ADD[1]),
    .B(_684_),
    .C(_687_),
    .Y(_688_)
);

OAI21X1 _3003_ (
    .A(_1324_),
    .B(_1080_),
    .C(_688_),
    .Y(_689_)
);

INVX1 _3004_ (
    .A(_689_),
    .Y(_690_)
);

AOI21X1 _3005_ (
    .A(_675_),
    .B(_690_),
    .C(_680_),
    .Y(_70_)
);

NOR2X1 _3006_ (
    .A(\AXYS[0] [2]),
    .B(_675_),
    .Y(_691_)
);

XNOR2X1 _3007_ (
    .A(_681_),
    .B(ADD[2]),
    .Y(_692_)
);

NAND2X1 _3008_ (
    .A(_692_),
    .B(_686_),
    .Y(_693_)
);

OAI21X1 _3009_ (
    .A(_899__bF$buf2),
    .B(_1313_),
    .C(_693_),
    .Y(_694_)
);

INVX1 _3010_ (
    .A(_694_),
    .Y(_695_)
);

OAI21X1 _3011_ (
    .A(_686_),
    .B(_692_),
    .C(_695_),
    .Y(_696_)
);

OAI21X1 _3012_ (
    .A(_838_),
    .B(_1080_),
    .C(_696_),
    .Y(_697_)
);

INVX1 _3013_ (
    .A(_697_),
    .Y(_698_)
);

AOI21X1 _3014_ (
    .A(_675_),
    .B(_698_),
    .C(_691_),
    .Y(_71_)
);

OAI21X1 _3015_ (
    .A(_627_),
    .B(_681_),
    .C(_693_),
    .Y(_699_)
);

XOR2X1 _3016_ (
    .A(_683_),
    .B(_618_),
    .Y(_700_)
);

XOR2X1 _3017_ (
    .A(_699_),
    .B(_700_),
    .Y(_701_)
);

OAI21X1 _3018_ (
    .A(_899__bF$buf1),
    .B(_1313_),
    .C(_701_),
    .Y(_702_)
);

OAI21X1 _3019_ (
    .A(_1327_),
    .B(_1080_),
    .C(_702_),
    .Y(_703_)
);

INVX1 _3020_ (
    .A(_703_),
    .Y(_704_)
);

NOR2X1 _3021_ (
    .A(\AXYS[0] [3]),
    .B(_675_),
    .Y(_705_)
);

AOI21X1 _3022_ (
    .A(_675_),
    .B(_704_),
    .C(_705_),
    .Y(_72_)
);

OAI21X1 _3023_ (
    .A(_899__bF$buf0),
    .B(_1313_),
    .C(ADD[4]),
    .Y(_706_)
);

OAI21X1 _3024_ (
    .A(_1329_),
    .B(_1080_),
    .C(_706_),
    .Y(_707_)
);

INVX1 _3025_ (
    .A(_707_),
    .Y(_708_)
);

NOR2X1 _3026_ (
    .A(\AXYS[0] [4]),
    .B(_675_),
    .Y(_709_)
);

AOI21X1 _3027_ (
    .A(_675_),
    .B(_708_),
    .C(_709_),
    .Y(_73_)
);

NOR2X1 _3028_ (
    .A(\AXYS[0] [5]),
    .B(_675_),
    .Y(_710_)
);

NAND3X1 _3029_ (
    .A(adj_bcd),
    .B(adc_bcd),
    .C(\ALU.CO ),
    .Y(_711_)
);

NOR2X1 _3030_ (
    .A(adc_bcd),
    .B(\ALU.CO ),
    .Y(_712_)
);

NAND2X1 _3031_ (
    .A(adj_bcd),
    .B(_712_),
    .Y(_713_)
);

NAND2X1 _3032_ (
    .A(_711_),
    .B(_713_),
    .Y(_714_)
);

INVX1 _3033_ (
    .A(ADD[5]),
    .Y(_715_)
);

INVX1 _3034_ (
    .A(_714_),
    .Y(_716_)
);

OAI21X1 _3035_ (
    .A(_715_),
    .B(_716_),
    .C(_1080_),
    .Y(_717_)
);

INVX1 _3036_ (
    .A(_717_),
    .Y(_718_)
);

OAI21X1 _3037_ (
    .A(ADD[5]),
    .B(_714_),
    .C(_718_),
    .Y(_719_)
);

OAI21X1 _3038_ (
    .A(_844_),
    .B(_1080_),
    .C(_719_),
    .Y(_720_)
);

INVX1 _3039_ (
    .A(_720_),
    .Y(_721_)
);

AOI21X1 _3040_ (
    .A(_675_),
    .B(_721_),
    .C(_710_),
    .Y(_74_)
);

NOR2X1 _3041_ (
    .A(\AXYS[0] [6]),
    .B(_675_),
    .Y(_722_)
);

NOR2X1 _3042_ (
    .A(_715_),
    .B(_716_),
    .Y(_723_)
);

XNOR2X1 _3043_ (
    .A(_711_),
    .B(ADD[6]),
    .Y(_724_)
);

AOI21X1 _3044_ (
    .A(_723_),
    .B(_724_),
    .C(_1081_),
    .Y(_725_)
);

OAI21X1 _3045_ (
    .A(_723_),
    .B(_724_),
    .C(_725_),
    .Y(_726_)
);

OAI21X1 _3046_ (
    .A(_846_),
    .B(_1080_),
    .C(_726_),
    .Y(_727_)
);

INVX1 _3047_ (
    .A(_727_),
    .Y(_728_)
);

AOI21X1 _3048_ (
    .A(_675_),
    .B(_728_),
    .C(_722_),
    .Y(_75_)
);

NAND2X1 _3049_ (
    .A(_724_),
    .B(_723_),
    .Y(_729_)
);

OAI21X1 _3050_ (
    .A(_608_),
    .B(_711_),
    .C(_729_),
    .Y(_730_)
);

XNOR2X1 _3051_ (
    .A(_713_),
    .B(\ALU.N ),
    .Y(_731_)
);

XOR2X1 _3052_ (
    .A(_730_),
    .B(_731_),
    .Y(_732_)
);

OAI21X1 _3053_ (
    .A(_899__bF$buf4),
    .B(_1313_),
    .C(_732_),
    .Y(_733_)
);

OAI21X1 _3054_ (
    .A(_847_),
    .B(_1080_),
    .C(_733_),
    .Y(_734_)
);

INVX1 _3055_ (
    .A(_734_),
    .Y(_735_)
);

NOR2X1 _3056_ (
    .A(\AXYS[0] [7]),
    .B(_675_),
    .Y(_736_)
);

AOI21X1 _3057_ (
    .A(_675_),
    .B(_735_),
    .C(_736_),
    .Y(_76_)
);

INVX2 _3058_ (
    .A(_1361_),
    .Y(_737_)
);

OR2X2 _3059_ (
    .A(_737_),
    .B(_674_),
    .Y(_738_)
);

OAI21X1 _3060_ (
    .A(_674_),
    .B(_737_),
    .C(\AXYS[1] [0]),
    .Y(_739_)
);

OAI21X1 _3061_ (
    .A(_678_),
    .B(_738_),
    .C(_739_),
    .Y(_77_)
);

OAI21X1 _3062_ (
    .A(_674_),
    .B(_737_),
    .C(\AXYS[1] [1]),
    .Y(_740_)
);

OAI21X1 _3063_ (
    .A(_690_),
    .B(_738_),
    .C(_740_),
    .Y(_78_)
);

OAI21X1 _3064_ (
    .A(_674_),
    .B(_737_),
    .C(\AXYS[1] [2]),
    .Y(_741_)
);

OAI21X1 _3065_ (
    .A(_698_),
    .B(_738_),
    .C(_741_),
    .Y(_79_)
);

OAI21X1 _3066_ (
    .A(_674_),
    .B(_737_),
    .C(\AXYS[1] [3]),
    .Y(_742_)
);

OAI21X1 _3067_ (
    .A(_704_),
    .B(_738_),
    .C(_742_),
    .Y(_80_)
);

OAI21X1 _3068_ (
    .A(_674_),
    .B(_737_),
    .C(\AXYS[1] [4]),
    .Y(_743_)
);

OAI21X1 _3069_ (
    .A(_708_),
    .B(_738_),
    .C(_743_),
    .Y(_81_)
);

OAI21X1 _3070_ (
    .A(_674_),
    .B(_737_),
    .C(\AXYS[1] [5]),
    .Y(_744_)
);

OAI21X1 _3071_ (
    .A(_721_),
    .B(_738_),
    .C(_744_),
    .Y(_82_)
);

OAI21X1 _3072_ (
    .A(_674_),
    .B(_737_),
    .C(\AXYS[1] [6]),
    .Y(_745_)
);

OAI21X1 _3073_ (
    .A(_728_),
    .B(_738_),
    .C(_745_),
    .Y(_83_)
);

OAI21X1 _3074_ (
    .A(_674_),
    .B(_737_),
    .C(\AXYS[1] [7]),
    .Y(_746_)
);

OAI21X1 _3075_ (
    .A(_735_),
    .B(_738_),
    .C(_746_),
    .Y(_84_)
);

INVX1 _3076_ (
    .A(_1365_),
    .Y(_747_)
);

NOR2X1 _3077_ (
    .A(_674_),
    .B(_747_),
    .Y(_748_)
);

NOR2X1 _3078_ (
    .A(\AXYS[2] [0]),
    .B(_748_),
    .Y(_749_)
);

AOI21X1 _3079_ (
    .A(_678_),
    .B(_748_),
    .C(_749_),
    .Y(_85_)
);

NOR2X1 _3080_ (
    .A(\AXYS[2] [1]),
    .B(_748_),
    .Y(_750_)
);

AOI21X1 _3081_ (
    .A(_690_),
    .B(_748_),
    .C(_750_),
    .Y(_86_)
);

NOR2X1 _3082_ (
    .A(\AXYS[2] [2]),
    .B(_748_),
    .Y(_751_)
);

AOI21X1 _3083_ (
    .A(_698_),
    .B(_748_),
    .C(_751_),
    .Y(_87_)
);

NOR2X1 _3084_ (
    .A(\AXYS[2] [3]),
    .B(_748_),
    .Y(_752_)
);

AOI21X1 _3085_ (
    .A(_704_),
    .B(_748_),
    .C(_752_),
    .Y(_88_)
);

NOR2X1 _3086_ (
    .A(\AXYS[2] [4]),
    .B(_748_),
    .Y(_753_)
);

AOI21X1 _3087_ (
    .A(_708_),
    .B(_748_),
    .C(_753_),
    .Y(_89_)
);

NOR2X1 _3088_ (
    .A(\AXYS[2] [5]),
    .B(_748_),
    .Y(_754_)
);

AOI21X1 _3089_ (
    .A(_721_),
    .B(_748_),
    .C(_754_),
    .Y(_90_)
);

NOR2X1 _3090_ (
    .A(\AXYS[2] [6]),
    .B(_748_),
    .Y(_755_)
);

AOI21X1 _3091_ (
    .A(_728_),
    .B(_748_),
    .C(_755_),
    .Y(_91_)
);

NOR2X1 _3092_ (
    .A(\AXYS[2] [7]),
    .B(_748_),
    .Y(_756_)
);

AOI21X1 _3093_ (
    .A(_735_),
    .B(_748_),
    .C(_756_),
    .Y(_92_)
);

INVX1 _3094_ (
    .A(_1366_),
    .Y(_757_)
);

NOR2X1 _3095_ (
    .A(_674_),
    .B(_757_),
    .Y(_758_)
);

NOR2X1 _3096_ (
    .A(\AXYS[3] [0]),
    .B(_758_),
    .Y(_759_)
);

AOI21X1 _3097_ (
    .A(_678_),
    .B(_758_),
    .C(_759_),
    .Y(_93_)
);

NOR2X1 _3098_ (
    .A(\AXYS[3] [1]),
    .B(_758_),
    .Y(_760_)
);

AOI21X1 _3099_ (
    .A(_690_),
    .B(_758_),
    .C(_760_),
    .Y(_94_)
);

NOR2X1 _3100_ (
    .A(\AXYS[3] [2]),
    .B(_758_),
    .Y(_761_)
);

AOI21X1 _3101_ (
    .A(_698_),
    .B(_758_),
    .C(_761_),
    .Y(_95_)
);

NOR2X1 _3102_ (
    .A(\AXYS[3] [3]),
    .B(_758_),
    .Y(_762_)
);

AOI21X1 _3103_ (
    .A(_704_),
    .B(_758_),
    .C(_762_),
    .Y(_96_)
);

NOR2X1 _3104_ (
    .A(\AXYS[3] [4]),
    .B(_758_),
    .Y(_763_)
);

AOI21X1 _3105_ (
    .A(_708_),
    .B(_758_),
    .C(_763_),
    .Y(_97_)
);

NOR2X1 _3106_ (
    .A(\AXYS[3] [5]),
    .B(_758_),
    .Y(_764_)
);

AOI21X1 _3107_ (
    .A(_721_),
    .B(_758_),
    .C(_764_),
    .Y(_98_)
);

NOR2X1 _3108_ (
    .A(\AXYS[3] [6]),
    .B(_758_),
    .Y(_765_)
);

AOI21X1 _3109_ (
    .A(_728_),
    .B(_758_),
    .C(_765_),
    .Y(_99_)
);

NOR2X1 _3110_ (
    .A(\AXYS[3] [7]),
    .B(_758_),
    .Y(_766_)
);

AOI21X1 _3111_ (
    .A(_735_),
    .B(_758_),
    .C(_766_),
    .Y(_100_)
);

OAI21X1 _3112_ (
    .A(_851_),
    .B(_931_),
    .C(_1106_),
    .Y(_767_)
);

OAI21X1 _3113_ (
    .A(_853_),
    .B(_914_),
    .C(_767_),
    .Y(_768_)
);

NAND2X1 _3114_ (
    .A(_1373_),
    .B(_768_),
    .Y(_769_)
);

OAI21X1 _3115_ (
    .A(_899__bF$buf3),
    .B(_905_),
    .C(_859__bF$buf2),
    .Y(_770_)
);

NOR2X1 _3116_ (
    .A(_770_),
    .B(_1204_),
    .Y(_771_)
);

NOR2X1 _3117_ (
    .A(_1210_),
    .B(_991_),
    .Y(_772_)
);

AOI21X1 _3118_ (
    .A(_1339_),
    .B(_914_),
    .C(_1007_),
    .Y(_773_)
);

AND2X2 _3119_ (
    .A(_772_),
    .B(_773_),
    .Y(_774_)
);

NAND3X1 _3120_ (
    .A(_1334_),
    .B(_771_),
    .C(_774_),
    .Y(_775_)
);

NOR2X1 _3121_ (
    .A(_769_),
    .B(_775_),
    .Y(_776_)
);

OAI21X1 _3122_ (
    .A(_1051_),
    .B(_1144_),
    .C(_916_),
    .Y(_777_)
);

OAI21X1 _3123_ (
    .A(_853_),
    .B(state[4]),
    .C(_1009_),
    .Y(_778_)
);

AND2X2 _3124_ (
    .A(_777_),
    .B(_778_),
    .Y(_779_)
);

NAND3X1 _3125_ (
    .A(_1052_),
    .B(_771_),
    .C(_774_),
    .Y(_780_)
);

OAI21X1 _3126_ (
    .A(_917__bF$buf0),
    .B(_990_),
    .C(_772_),
    .Y(_781_)
);

OR2X2 _3127_ (
    .A(_781_),
    .B(_770_),
    .Y(_782_)
);

AOI22X1 _3128_ (
    .A(_856__bF$buf1),
    .B(_1007_),
    .C(_1051_),
    .D(_914_),
    .Y(_783_)
);

NOR2X1 _3129_ (
    .A(_1227_),
    .B(_1204_),
    .Y(_784_)
);

NAND3X1 _3130_ (
    .A(_1374_),
    .B(_784_),
    .C(_783_),
    .Y(_785_)
);

OAI21X1 _3131_ (
    .A(_785_),
    .B(_782_),
    .C(_780_),
    .Y(_786_)
);

INVX1 _3132_ (
    .A(_769_),
    .Y(_787_)
);

OAI21X1 _3133_ (
    .A(_923__bF$buf2),
    .B(_1313_),
    .C(_1334_),
    .Y(_788_)
);

NAND3X1 _3134_ (
    .A(_913_),
    .B(_1057_),
    .C(_1286_),
    .Y(_789_)
);

NOR2X1 _3135_ (
    .A(_788_),
    .B(_789_),
    .Y(_790_)
);

AND2X2 _3136_ (
    .A(_790_),
    .B(_787_),
    .Y(_791_)
);

AOI22X1 _3137_ (
    .A(_779_),
    .B(_776_),
    .C(_786_),
    .D(_791_),
    .Y(_792_)
);

AOI21X1 _3138_ (
    .A(_900_),
    .B(_938_),
    .C(_670_),
    .Y(_793_)
);

OAI21X1 _3139_ (
    .A(_917__bF$buf4),
    .B(_921_),
    .C(_1045_),
    .Y(_794_)
);

NOR2X1 _3140_ (
    .A(_292_),
    .B(_794_),
    .Y(_795_)
);

AND2X2 _3141_ (
    .A(_795_),
    .B(_793_),
    .Y(_796_)
);

INVX1 _3142_ (
    .A(_184_),
    .Y(_797_)
);

NOR2X1 _3143_ (
    .A(_797_),
    .B(_1308_),
    .Y(_798_)
);

OAI21X1 _3144_ (
    .A(_854__bF$buf2),
    .B(_900_),
    .C(_852_),
    .Y(_799_)
);

OAI21X1 _3145_ (
    .A(state[4]),
    .B(_1062_),
    .C(_799_),
    .Y(_800_)
);

INVX1 _3146_ (
    .A(_800_),
    .Y(_801_)
);

AND2X2 _3147_ (
    .A(_801_),
    .B(_1319_),
    .Y(_802_)
);

NAND3X1 _3148_ (
    .A(_798_),
    .B(_802_),
    .C(_796_),
    .Y(_803_)
);

OAI21X1 _3149_ (
    .A(_923__bF$buf1),
    .B(_1082_),
    .C(_291_),
    .Y(_804_)
);

OAI21X1 _3150_ (
    .A(_856__bF$buf0),
    .B(_913_),
    .C(_1057_),
    .Y(_805_)
);

NOR2X1 _3151_ (
    .A(_804_),
    .B(_805_),
    .Y(_806_)
);

AND2X2 _3152_ (
    .A(_806_),
    .B(_1319_),
    .Y(_807_)
);

NAND3X1 _3153_ (
    .A(_798_),
    .B(_801_),
    .C(_807_),
    .Y(_808_)
);

OAI21X1 _3154_ (
    .A(_938_),
    .B(_1009_),
    .C(_856__bF$buf3),
    .Y(_809_)
);

INVX1 _3155_ (
    .A(_939_),
    .Y(_810_)
);

NOR2X1 _3156_ (
    .A(_810_),
    .B(_794_),
    .Y(_811_)
);

NAND3X1 _3157_ (
    .A(_777_),
    .B(_809_),
    .C(_811_),
    .Y(_812_)
);

NOR2X1 _3158_ (
    .A(_812_),
    .B(_808_),
    .Y(_813_)
);

AOI21X1 _3159_ (
    .A(_813_),
    .B(_776_),
    .C(_836__bF$buf1),
    .Y(_814_)
);

OAI21X1 _3160_ (
    .A(_792_),
    .B(_803_),
    .C(_814_),
    .Y(_815_)
);

NAND2X1 _3161_ (
    .A(ABL[0]),
    .B(_815__bF$buf4),
    .Y(_816_)
);

OAI21X1 _3162_ (
    .A(_815__bF$buf3),
    .B(_205_),
    .C(_816_),
    .Y(_101_)
);

NAND2X1 _3163_ (
    .A(ABL[1]),
    .B(_815__bF$buf2),
    .Y(_817_)
);

OAI21X1 _3164_ (
    .A(_815__bF$buf1),
    .B(_212_),
    .C(_817_),
    .Y(_102_)
);

NAND2X1 _3165_ (
    .A(ABL[2]),
    .B(_815__bF$buf0),
    .Y(_818_)
);

OAI21X1 _3166_ (
    .A(_815__bF$buf4),
    .B(_217_),
    .C(_818_),
    .Y(_103_)
);

NAND2X1 _3167_ (
    .A(ABL[3]),
    .B(_815__bF$buf3),
    .Y(_819_)
);

OAI21X1 _3168_ (
    .A(_815__bF$buf2),
    .B(_222_),
    .C(_819_),
    .Y(_104_)
);

NAND2X1 _3169_ (
    .A(ABL[4]),
    .B(_815__bF$buf1),
    .Y(_820_)
);

OAI21X1 _3170_ (
    .A(_815__bF$buf0),
    .B(_228_),
    .C(_820_),
    .Y(_105_)
);

NAND2X1 _3171_ (
    .A(ABL[5]),
    .B(_815__bF$buf4),
    .Y(_821_)
);

OAI21X1 _3172_ (
    .A(_815__bF$buf3),
    .B(_233_),
    .C(_821_),
    .Y(_106_)
);

NAND2X1 _3173_ (
    .A(ABL[6]),
    .B(_815__bF$buf2),
    .Y(_822_)
);

OAI21X1 _3174_ (
    .A(_815__bF$buf1),
    .B(_238_),
    .C(_822_),
    .Y(_107_)
);

NAND2X1 _3175_ (
    .A(ABL[7]),
    .B(_815__bF$buf0),
    .Y(_823_)
);

OAI21X1 _3176_ (
    .A(_815__bF$buf4),
    .B(_243_),
    .C(_823_),
    .Y(_108_)
);

NOR2X1 _3177_ (
    .A(_815__bF$buf3),
    .B(_1665_[8]),
    .Y(_824_)
);

AOI21X1 _3178_ (
    .A(_1386_),
    .B(_815__bF$buf2),
    .C(_824_),
    .Y(_109_)
);

NOR2X1 _3179_ (
    .A(_815__bF$buf1),
    .B(_1665_[9]),
    .Y(_825_)
);

AOI21X1 _3180_ (
    .A(_250_),
    .B(_815__bF$buf0),
    .C(_825_),
    .Y(_110_)
);

NOR2X1 _3181_ (
    .A(_815__bF$buf4),
    .B(_1665_[10]),
    .Y(_826_)
);

AOI21X1 _3182_ (
    .A(_1403_),
    .B(_815__bF$buf3),
    .C(_826_),
    .Y(_111_)
);

NOR2X1 _3183_ (
    .A(_815__bF$buf2),
    .B(_1665_[11]),
    .Y(_827_)
);

AOI21X1 _3184_ (
    .A(_261_),
    .B(_815__bF$buf1),
    .C(_827_),
    .Y(_112_)
);

NOR2X1 _3185_ (
    .A(_815__bF$buf0),
    .B(_1665_[12]),
    .Y(_828_)
);

AOI21X1 _3186_ (
    .A(_265_),
    .B(_815__bF$buf4),
    .C(_828_),
    .Y(_113_)
);

NOR2X1 _3187_ (
    .A(_815__bF$buf3),
    .B(_1665_[13]),
    .Y(_829_)
);

AOI21X1 _3188_ (
    .A(_274_),
    .B(_815__bF$buf2),
    .C(_829_),
    .Y(_114_)
);

NOR2X1 _3189_ (
    .A(_815__bF$buf1),
    .B(_1665_[14]),
    .Y(_830_)
);

AOI21X1 _3190_ (
    .A(_1437_),
    .B(_815__bF$buf0),
    .C(_830_),
    .Y(_115_)
);

NOR2X1 _3191_ (
    .A(_815__bF$buf4),
    .B(_1665_[15]),
    .Y(_831_)
);

AOI21X1 _3192_ (
    .A(_1447_),
    .B(_815__bF$buf3),
    .C(_831_),
    .Y(_116_)
);

DFFSR _3193_ (
    .CLK(clk_bF$buf10),
    .D(_1463_[0]),
    .Q(state[0]),
    .R(_1__bF$buf10),
    .S(vdd)
);

DFFSR _3194_ (
    .CLK(clk_bF$buf9),
    .D(_1463_[1]),
    .Q(state[1]),
    .R(_1__bF$buf9),
    .S(vdd)
);

DFFSR _3195_ (
    .CLK(clk_bF$buf8),
    .D(_1463_[2]),
    .Q(state[2]),
    .R(_1__bF$buf8),
    .S(vdd)
);

DFFSR _3196_ (
    .CLK(clk_bF$buf7),
    .D(_1463_[3]),
    .Q(state[3]),
    .R(vdd),
    .S(_1__bF$buf7)
);

DFFSR _3197_ (
    .CLK(clk_bF$buf6),
    .D(_1463_[4]),
    .Q(state[4]),
    .R(_1__bF$buf6),
    .S(vdd)
);

DFFSR _3198_ (
    .CLK(clk_bF$buf5),
    .D(_1463_[5]),
    .Q(state[5]),
    .R(_1__bF$buf5),
    .S(vdd)
);

DFFSR _3199_ (
    .CLK(clk_bF$buf4),
    .D(_2_),
    .Q(PC[0]),
    .R(_1__bF$buf4),
    .S(vdd)
);

DFFSR _3200_ (
    .CLK(clk_bF$buf3),
    .D(_3_),
    .Q(PC[1]),
    .R(_1__bF$buf3),
    .S(vdd)
);

DFFSR _3201_ (
    .CLK(clk_bF$buf2),
    .D(_4_),
    .Q(PC[2]),
    .R(_1__bF$buf2),
    .S(vdd)
);

DFFSR _3202_ (
    .CLK(clk_bF$buf1),
    .D(_5_),
    .Q(PC[3]),
    .R(_1__bF$buf1),
    .S(vdd)
);

DFFSR _3203_ (
    .CLK(clk_bF$buf0),
    .D(_6_),
    .Q(PC[4]),
    .R(_1__bF$buf0),
    .S(vdd)
);

DFFSR _3204_ (
    .CLK(clk_bF$buf10),
    .D(_7_),
    .Q(PC[5]),
    .R(_1__bF$buf10),
    .S(vdd)
);

DFFSR _3205_ (
    .CLK(clk_bF$buf9),
    .D(_8_),
    .Q(PC[6]),
    .R(_1__bF$buf9),
    .S(vdd)
);

DFFSR _3206_ (
    .CLK(clk_bF$buf8),
    .D(_9_),
    .Q(PC[7]),
    .R(_1__bF$buf8),
    .S(vdd)
);

DFFSR _3207_ (
    .CLK(clk_bF$buf7),
    .D(_10_),
    .Q(PC[8]),
    .R(_1__bF$buf7),
    .S(vdd)
);

DFFSR _3208_ (
    .CLK(clk_bF$buf6),
    .D(_11_),
    .Q(PC[9]),
    .R(_1__bF$buf6),
    .S(vdd)
);

DFFSR _3209_ (
    .CLK(clk_bF$buf5),
    .D(_12_),
    .Q(PC[10]),
    .R(_1__bF$buf5),
    .S(vdd)
);

DFFSR _3210_ (
    .CLK(clk_bF$buf4),
    .D(_13_),
    .Q(PC[11]),
    .R(_1__bF$buf4),
    .S(vdd)
);

DFFSR _3211_ (
    .CLK(clk_bF$buf3),
    .D(_14_),
    .Q(PC[12]),
    .R(_1__bF$buf3),
    .S(vdd)
);

DFFSR _3212_ (
    .CLK(clk_bF$buf2),
    .D(_15_),
    .Q(PC[13]),
    .R(_1__bF$buf2),
    .S(vdd)
);

DFFSR _3213_ (
    .CLK(clk_bF$buf1),
    .D(_16_),
    .Q(PC[14]),
    .R(_1__bF$buf1),
    .S(vdd)
);

DFFSR _3214_ (
    .CLK(clk_bF$buf0),
    .D(_17_),
    .Q(PC[15]),
    .R(_1__bF$buf0),
    .S(vdd)
);

DFFSR _3215_ (
    .CLK(clk_bF$buf10),
    .D(NMI),
    .Q(NMI_1),
    .R(_1__bF$buf10),
    .S(vdd)
);

DFFSR _3216_ (
    .CLK(clk_bF$buf9),
    .D(_18_),
    .Q(NMI_edge),
    .R(_1__bF$buf9),
    .S(vdd)
);

DFFSR _3217_ (
    .CLK(clk_bF$buf8),
    .D(_19_),
    .Q(cond_code[0]),
    .R(_1__bF$buf8),
    .S(vdd)
);

DFFSR _3218_ (
    .CLK(clk_bF$buf7),
    .D(_20_),
    .Q(cond_code[1]),
    .R(_1__bF$buf7),
    .S(vdd)
);

DFFSR _3219_ (
    .CLK(clk_bF$buf6),
    .D(_21_),
    .Q(cond_code[2]),
    .R(_1__bF$buf6),
    .S(vdd)
);

DFFSR _3220_ (
    .CLK(clk_bF$buf5),
    .D(_22_),
    .Q(plp),
    .R(_1__bF$buf5),
    .S(vdd)
);

DFFSR _3221_ (
    .CLK(clk_bF$buf4),
    .D(_23_),
    .Q(php),
    .R(_1__bF$buf4),
    .S(vdd)
);

DFFSR _3222_ (
    .CLK(clk_bF$buf3),
    .D(_24_),
    .Q(clc),
    .R(_1__bF$buf3),
    .S(vdd)
);

DFFSR _3223_ (
    .CLK(clk_bF$buf2),
    .D(_25_),
    .Q(sec),
    .R(_1__bF$buf2),
    .S(vdd)
);

DFFSR _3224_ (
    .CLK(clk_bF$buf1),
    .D(_26_),
    .Q(cld),
    .R(_1__bF$buf1),
    .S(vdd)
);

DFFSR _3225_ (
    .CLK(clk_bF$buf0),
    .D(_27_),
    .Q(sed),
    .R(_1__bF$buf0),
    .S(vdd)
);

DFFSR _3226_ (
    .CLK(clk_bF$buf10),
    .D(_28_),
    .Q(cli),
    .R(_1__bF$buf10),
    .S(vdd)
);

DFFSR _3227_ (
    .CLK(clk_bF$buf9),
    .D(_29_),
    .Q(sei),
    .R(_1__bF$buf9),
    .S(vdd)
);

DFFSR _3228_ (
    .CLK(clk_bF$buf8),
    .D(_30_),
    .Q(clv),
    .R(_1__bF$buf8),
    .S(vdd)
);

DFFSR _3229_ (
    .CLK(clk_bF$buf7),
    .D(_31_),
    .Q(bit_ins),
    .R(_1__bF$buf7),
    .S(vdd)
);

DFFSR _3230_ (
    .CLK(clk_bF$buf6),
    .D(_32_),
    .Q(op[0]),
    .R(_1__bF$buf6),
    .S(vdd)
);

DFFSR _3231_ (
    .CLK(clk_bF$buf5),
    .D(_33_),
    .Q(op[1]),
    .R(_1__bF$buf5),
    .S(vdd)
);

DFFSR _3232_ (
    .CLK(clk_bF$buf4),
    .D(_34_),
    .Q(op[2]),
    .R(_1__bF$buf4),
    .S(vdd)
);

DFFSR _3233_ (
    .CLK(clk_bF$buf3),
    .D(_35_),
    .Q(op[3]),
    .R(_1__bF$buf3),
    .S(vdd)
);

DFFSR _3234_ (
    .CLK(clk_bF$buf2),
    .D(_36_),
    .Q(rotate),
    .R(_1__bF$buf2),
    .S(vdd)
);

DFFSR _3235_ (
    .CLK(clk_bF$buf1),
    .D(_37_),
    .Q(shift_right),
    .R(_1__bF$buf1),
    .S(vdd)
);

DFFSR _3236_ (
    .CLK(clk_bF$buf0),
    .D(_38_),
    .Q(compare),
    .R(_1__bF$buf0),
    .S(vdd)
);

DFFSR _3237_ (
    .CLK(clk_bF$buf10),
    .D(_39_),
    .Q(shift),
    .R(_1__bF$buf10),
    .S(vdd)
);

DFFSR _3238_ (
    .CLK(clk_bF$buf9),
    .D(_40_),
    .Q(adc_bcd),
    .R(_1__bF$buf9),
    .S(vdd)
);

DFFSR _3239_ (
    .CLK(clk_bF$buf8),
    .D(_41_),
    .Q(adc_sbc),
    .R(_1__bF$buf8),
    .S(vdd)
);

DFFSR _3240_ (
    .CLK(clk_bF$buf7),
    .D(_42_),
    .Q(inc),
    .R(_1__bF$buf7),
    .S(vdd)
);

DFFSR _3241_ (
    .CLK(clk_bF$buf6),
    .D(_43_),
    .Q(load_only),
    .R(_1__bF$buf6),
    .S(vdd)
);

DFFSR _3242_ (
    .CLK(clk_bF$buf5),
    .D(_44_),
    .Q(write_back),
    .R(_1__bF$buf5),
    .S(vdd)
);

DFFSR _3243_ (
    .CLK(clk_bF$buf4),
    .D(_45_),
    .Q(store),
    .R(_1__bF$buf4),
    .S(vdd)
);

DFFSR _3244_ (
    .CLK(clk_bF$buf3),
    .D(_46_),
    .Q(index_y),
    .R(_1__bF$buf3),
    .S(vdd)
);

DFFSR _3245_ (
    .CLK(clk_bF$buf2),
    .D(_47_),
    .Q(src_reg[0]),
    .R(_1__bF$buf2),
    .S(vdd)
);

DFFSR _3246_ (
    .CLK(clk_bF$buf1),
    .D(_48_),
    .Q(src_reg[1]),
    .R(_1__bF$buf1),
    .S(vdd)
);

DFFSR _3247_ (
    .CLK(clk_bF$buf0),
    .D(_49_),
    .Q(dst_reg[0]),
    .R(_1__bF$buf0),
    .S(vdd)
);

DFFSR _3248_ (
    .CLK(clk_bF$buf10),
    .D(_50_),
    .Q(dst_reg[1]),
    .R(_1__bF$buf10),
    .S(vdd)
);

DFFSR _3249_ (
    .CLK(clk_bF$buf9),
    .D(_51_),
    .Q(load_reg),
    .R(_1__bF$buf9),
    .S(vdd)
);

DFFSR _3250_ (
    .CLK(clk_bF$buf8),
    .D(DIMUX[0]),
    .Q(DIHOLD[0]),
    .R(_1__bF$buf8),
    .S(vdd)
);

DFFSR _3251_ (
    .CLK(clk_bF$buf7),
    .D(DIMUX[1]),
    .Q(DIHOLD[1]),
    .R(_1__bF$buf7),
    .S(vdd)
);

DFFSR _3252_ (
    .CLK(clk_bF$buf6),
    .D(DIMUX[2]),
    .Q(DIHOLD[2]),
    .R(_1__bF$buf6),
    .S(vdd)
);

DFFSR _3253_ (
    .CLK(clk_bF$buf5),
    .D(DIMUX[3]),
    .Q(DIHOLD[3]),
    .R(_1__bF$buf5),
    .S(vdd)
);

DFFSR _3254_ (
    .CLK(clk_bF$buf4),
    .D(DIMUX[4]),
    .Q(DIHOLD[4]),
    .R(_1__bF$buf4),
    .S(vdd)
);

DFFSR _3255_ (
    .CLK(clk_bF$buf3),
    .D(DIMUX[5]),
    .Q(DIHOLD[5]),
    .R(_1__bF$buf3),
    .S(vdd)
);

DFFSR _3256_ (
    .CLK(clk_bF$buf2),
    .D(DIMUX[6]),
    .Q(DIHOLD[6]),
    .R(_1__bF$buf2),
    .S(vdd)
);

DFFSR _3257_ (
    .CLK(clk_bF$buf1),
    .D(DIMUX[7]),
    .Q(DIHOLD[7]),
    .R(_1__bF$buf1),
    .S(vdd)
);

DFFSR _3258_ (
    .CLK(clk_bF$buf0),
    .D(_52_),
    .Q(res),
    .R(vdd),
    .S(_1__bF$buf0)
);

DFFPOSX1 _3259_ (
    .CLK(clk_bF$buf10),
    .D(_53_),
    .Q(IRHOLD[0])
);

DFFPOSX1 _3260_ (
    .CLK(clk_bF$buf9),
    .D(_54_),
    .Q(IRHOLD[1])
);

DFFPOSX1 _3261_ (
    .CLK(clk_bF$buf8),
    .D(_55_),
    .Q(IRHOLD[2])
);

DFFPOSX1 _3262_ (
    .CLK(clk_bF$buf7),
    .D(_56_),
    .Q(IRHOLD[3])
);

DFFPOSX1 _3263_ (
    .CLK(clk_bF$buf6),
    .D(_57_),
    .Q(IRHOLD[4])
);

DFFPOSX1 _3264_ (
    .CLK(clk_bF$buf5),
    .D(_58_),
    .Q(IRHOLD[5])
);

DFFPOSX1 _3265_ (
    .CLK(clk_bF$buf4),
    .D(_59_),
    .Q(IRHOLD[6])
);

DFFPOSX1 _3266_ (
    .CLK(clk_bF$buf3),
    .D(_60_),
    .Q(IRHOLD[7])
);

DFFSR _3267_ (
    .CLK(clk_bF$buf2),
    .D(_61_),
    .Q(IRHOLD_valid),
    .R(_1__bF$buf10),
    .S(vdd)
);

DFFSR _3268_ (
    .CLK(clk_bF$buf1),
    .D(_62_),
    .Q(V),
    .R(_1__bF$buf9),
    .S(vdd)
);

DFFSR _3269_ (
    .CLK(clk_bF$buf0),
    .D(_63_),
    .Q(D),
    .R(_1__bF$buf8),
    .S(vdd)
);

DFFSR _3270_ (
    .CLK(clk_bF$buf10),
    .D(_64_),
    .Q(I),
    .R(_1__bF$buf7),
    .S(vdd)
);

DFFSR _3271_ (
    .CLK(clk_bF$buf9),
    .D(_65_),
    .Q(N),
    .R(_1__bF$buf6),
    .S(vdd)
);

DFFSR _3272_ (
    .CLK(clk_bF$buf8),
    .D(_66_),
    .Q(Z),
    .R(_1__bF$buf5),
    .S(vdd)
);

DFFSR _3273_ (
    .CLK(clk_bF$buf7),
    .D(_67_),
    .Q(C),
    .R(_1__bF$buf4),
    .S(vdd)
);

DFFSR _3274_ (
    .CLK(clk_bF$buf6),
    .D(_68_),
    .Q(backwards),
    .R(_1__bF$buf3),
    .S(vdd)
);

DFFSR _3275_ (
    .CLK(clk_bF$buf5),
    .D(_69_),
    .Q(\AXYS[0] [0]),
    .R(_1__bF$buf2),
    .S(vdd)
);

DFFSR _3276_ (
    .CLK(clk_bF$buf4),
    .D(_70_),
    .Q(\AXYS[0] [1]),
    .R(_1__bF$buf1),
    .S(vdd)
);

DFFSR _3277_ (
    .CLK(clk_bF$buf3),
    .D(_71_),
    .Q(\AXYS[0] [2]),
    .R(_1__bF$buf0),
    .S(vdd)
);

DFFSR _3278_ (
    .CLK(clk_bF$buf2),
    .D(_72_),
    .Q(\AXYS[0] [3]),
    .R(_1__bF$buf10),
    .S(vdd)
);

DFFSR _3279_ (
    .CLK(clk_bF$buf1),
    .D(_73_),
    .Q(\AXYS[0] [4]),
    .R(_1__bF$buf9),
    .S(vdd)
);

DFFSR _3280_ (
    .CLK(clk_bF$buf0),
    .D(_74_),
    .Q(\AXYS[0] [5]),
    .R(_1__bF$buf8),
    .S(vdd)
);

DFFSR _3281_ (
    .CLK(clk_bF$buf10),
    .D(_75_),
    .Q(\AXYS[0] [6]),
    .R(_1__bF$buf7),
    .S(vdd)
);

DFFSR _3282_ (
    .CLK(clk_bF$buf9),
    .D(_76_),
    .Q(\AXYS[0] [7]),
    .R(_1__bF$buf6),
    .S(vdd)
);

DFFSR _3283_ (
    .CLK(clk_bF$buf8),
    .D(_77_),
    .Q(\AXYS[1] [0]),
    .R(_1__bF$buf5),
    .S(vdd)
);

DFFSR _3284_ (
    .CLK(clk_bF$buf7),
    .D(_78_),
    .Q(\AXYS[1] [1]),
    .R(_1__bF$buf4),
    .S(vdd)
);

DFFSR _3285_ (
    .CLK(clk_bF$buf6),
    .D(_79_),
    .Q(\AXYS[1] [2]),
    .R(_1__bF$buf3),
    .S(vdd)
);

DFFSR _3286_ (
    .CLK(clk_bF$buf5),
    .D(_80_),
    .Q(\AXYS[1] [3]),
    .R(_1__bF$buf2),
    .S(vdd)
);

DFFSR _3287_ (
    .CLK(clk_bF$buf4),
    .D(_81_),
    .Q(\AXYS[1] [4]),
    .R(_1__bF$buf1),
    .S(vdd)
);

DFFSR _3288_ (
    .CLK(clk_bF$buf3),
    .D(_82_),
    .Q(\AXYS[1] [5]),
    .R(_1__bF$buf0),
    .S(vdd)
);

DFFSR _3289_ (
    .CLK(clk_bF$buf2),
    .D(_83_),
    .Q(\AXYS[1] [6]),
    .R(_1__bF$buf10),
    .S(vdd)
);

DFFSR _3290_ (
    .CLK(clk_bF$buf1),
    .D(_84_),
    .Q(\AXYS[1] [7]),
    .R(_1__bF$buf9),
    .S(vdd)
);

DFFSR _3291_ (
    .CLK(clk_bF$buf0),
    .D(_85_),
    .Q(\AXYS[2] [0]),
    .R(_1__bF$buf8),
    .S(vdd)
);

DFFSR _3292_ (
    .CLK(clk_bF$buf10),
    .D(_86_),
    .Q(\AXYS[2] [1]),
    .R(_1__bF$buf7),
    .S(vdd)
);

DFFSR _3293_ (
    .CLK(clk_bF$buf9),
    .D(_87_),
    .Q(\AXYS[2] [2]),
    .R(_1__bF$buf6),
    .S(vdd)
);

DFFSR _3294_ (
    .CLK(clk_bF$buf8),
    .D(_88_),
    .Q(\AXYS[2] [3]),
    .R(_1__bF$buf5),
    .S(vdd)
);

DFFSR _3295_ (
    .CLK(clk_bF$buf7),
    .D(_89_),
    .Q(\AXYS[2] [4]),
    .R(_1__bF$buf4),
    .S(vdd)
);

DFFSR _3296_ (
    .CLK(clk_bF$buf6),
    .D(_90_),
    .Q(\AXYS[2] [5]),
    .R(_1__bF$buf3),
    .S(vdd)
);

DFFSR _3297_ (
    .CLK(clk_bF$buf5),
    .D(_91_),
    .Q(\AXYS[2] [6]),
    .R(_1__bF$buf2),
    .S(vdd)
);

DFFSR _3298_ (
    .CLK(clk_bF$buf4),
    .D(_92_),
    .Q(\AXYS[2] [7]),
    .R(_1__bF$buf1),
    .S(vdd)
);

DFFSR _3299_ (
    .CLK(clk_bF$buf3),
    .D(_0_),
    .Q(adj_bcd),
    .R(_1__bF$buf0),
    .S(vdd)
);

DFFSR _3300_ (
    .CLK(clk_bF$buf2),
    .D(_93_),
    .Q(\AXYS[3] [0]),
    .R(_1__bF$buf10),
    .S(vdd)
);

DFFSR _3301_ (
    .CLK(clk_bF$buf1),
    .D(_94_),
    .Q(\AXYS[3] [1]),
    .R(_1__bF$buf9),
    .S(vdd)
);

DFFSR _3302_ (
    .CLK(clk_bF$buf0),
    .D(_95_),
    .Q(\AXYS[3] [2]),
    .R(_1__bF$buf8),
    .S(vdd)
);

DFFSR _3303_ (
    .CLK(clk_bF$buf10),
    .D(_96_),
    .Q(\AXYS[3] [3]),
    .R(_1__bF$buf7),
    .S(vdd)
);

DFFSR _3304_ (
    .CLK(clk_bF$buf9),
    .D(_97_),
    .Q(\AXYS[3] [4]),
    .R(_1__bF$buf6),
    .S(vdd)
);

DFFSR _3305_ (
    .CLK(clk_bF$buf8),
    .D(_98_),
    .Q(\AXYS[3] [5]),
    .R(_1__bF$buf5),
    .S(vdd)
);

DFFSR _3306_ (
    .CLK(clk_bF$buf7),
    .D(_99_),
    .Q(\AXYS[3] [6]),
    .R(_1__bF$buf4),
    .S(vdd)
);

DFFSR _3307_ (
    .CLK(clk_bF$buf6),
    .D(_100_),
    .Q(\AXYS[3] [7]),
    .R(_1__bF$buf3),
    .S(vdd)
);

DFFSR _3308_ (
    .CLK(clk_bF$buf5),
    .D(_101_),
    .Q(ABL[0]),
    .R(_1__bF$buf2),
    .S(vdd)
);

DFFSR _3309_ (
    .CLK(clk_bF$buf4),
    .D(_102_),
    .Q(ABL[1]),
    .R(_1__bF$buf1),
    .S(vdd)
);

DFFSR _3310_ (
    .CLK(clk_bF$buf3),
    .D(_103_),
    .Q(ABL[2]),
    .R(_1__bF$buf0),
    .S(vdd)
);

DFFSR _3311_ (
    .CLK(clk_bF$buf2),
    .D(_104_),
    .Q(ABL[3]),
    .R(_1__bF$buf10),
    .S(vdd)
);

DFFSR _3312_ (
    .CLK(clk_bF$buf1),
    .D(_105_),
    .Q(ABL[4]),
    .R(_1__bF$buf9),
    .S(vdd)
);

DFFSR _3313_ (
    .CLK(clk_bF$buf0),
    .D(_106_),
    .Q(ABL[5]),
    .R(_1__bF$buf8),
    .S(vdd)
);

DFFSR _3314_ (
    .CLK(clk_bF$buf10),
    .D(_107_),
    .Q(ABL[6]),
    .R(_1__bF$buf7),
    .S(vdd)
);

DFFSR _3315_ (
    .CLK(clk_bF$buf9),
    .D(_108_),
    .Q(ABL[7]),
    .R(_1__bF$buf6),
    .S(vdd)
);

DFFSR _3316_ (
    .CLK(clk_bF$buf8),
    .D(_109_),
    .Q(ABH[0]),
    .R(_1__bF$buf5),
    .S(vdd)
);

DFFSR _3317_ (
    .CLK(clk_bF$buf7),
    .D(_110_),
    .Q(ABH[1]),
    .R(_1__bF$buf4),
    .S(vdd)
);

DFFSR _3318_ (
    .CLK(clk_bF$buf6),
    .D(_111_),
    .Q(ABH[2]),
    .R(_1__bF$buf3),
    .S(vdd)
);

DFFSR _3319_ (
    .CLK(clk_bF$buf5),
    .D(_112_),
    .Q(ABH[3]),
    .R(_1__bF$buf2),
    .S(vdd)
);

DFFSR _3320_ (
    .CLK(clk_bF$buf4),
    .D(_113_),
    .Q(ABH[4]),
    .R(_1__bF$buf1),
    .S(vdd)
);

DFFSR _3321_ (
    .CLK(clk_bF$buf3),
    .D(_114_),
    .Q(ABH[5]),
    .R(_1__bF$buf0),
    .S(vdd)
);

DFFSR _3322_ (
    .CLK(clk_bF$buf2),
    .D(_115_),
    .Q(ABH[6]),
    .R(_1__bF$buf10),
    .S(vdd)
);

DFFSR _3323_ (
    .CLK(clk_bF$buf1),
    .D(_116_),
    .Q(ABH[7]),
    .R(_1__bF$buf9),
    .S(vdd)
);

OR2X2 _3324_ (
    .A(ADD[0]),
    .B(ADD[3]),
    .Y(_1622_)
);

NOR2X1 _3325_ (
    .A(ADD[5]),
    .B(ADD[4]),
    .Y(_1623_)
);

NOR2X1 _3326_ (
    .A(\ALU.N ),
    .B(ADD[6]),
    .Y(_1624_)
);

NOR2X1 _3327_ (
    .A(ADD[1]),
    .B(ADD[2]),
    .Y(_1625_)
);

NAND3X1 _3328_ (
    .A(_1623_),
    .B(_1624_),
    .C(_1625_),
    .Y(_1626_)
);

NOR2X1 _3329_ (
    .A(_1622_),
    .B(_1626_),
    .Y(\ALU.Z )
);

XOR2X1 _3330_ (
    .A(\ALU.AI7 ),
    .B(\ALU.CO ),
    .Y(_1627_)
);

XNOR2X1 _3331_ (
    .A(\ALU.N ),
    .B(\ALU.BI7 ),
    .Y(_1628_)
);

XNOR2X1 _3332_ (
    .A(_1627_),
    .B(_1628_),
    .Y(\ALU.V )
);

INVX4 _3333_ (
    .A(reset),
    .Y(_1464_)
);

INVX4 _3334_ (
    .A(RDY_bF$buf6),
    .Y(_1629_)
);

NAND2X1 _3335_ (
    .A(\ALU.right ),
    .B(\ALU.CI ),
    .Y(_1630_)
);

INVX2 _3336_ (
    .A(\ALU.op [1]),
    .Y(_1631_)
);

NAND2X1 _3337_ (
    .A(\ALU.op [0]),
    .B(_1631_),
    .Y(_1632_)
);

INVX2 _3338_ (
    .A(\ALU.op [0]),
    .Y(_1633_)
);

AND2X2 _3339_ (
    .A(_1633_),
    .B(\ALU.BI [7]),
    .Y(_1634_)
);

NAND2X1 _3340_ (
    .A(AI[7]),
    .B(_1634_),
    .Y(_1635_)
);

AOI22X1 _3341_ (
    .A(_1631_),
    .B(\ALU.BI [7]),
    .C(_1635_),
    .D(_1632_),
    .Y(_1636_)
);

INVX2 _3342_ (
    .A(\ALU.right ),
    .Y(_1637_)
);

OAI21X1 _3343_ (
    .A(AI[7]),
    .B(_1634_),
    .C(_1637_),
    .Y(_1638_)
);

OAI21X1 _3344_ (
    .A(_1638_),
    .B(_1636_),
    .C(_1630_),
    .Y(_1639_)
);

INVX4 _3345_ (
    .A(\ALU.op [3]),
    .Y(_1640_)
);

OAI21X1 _3346_ (
    .A(\ALU.op [2]),
    .B(\ALU.BI [7]),
    .C(_1640_),
    .Y(_1641_)
);

AOI21X1 _3347_ (
    .A(\ALU.op [2]),
    .B(\ALU.BI [7]),
    .C(_1641_),
    .Y(_1642_)
);

NOR2X1 _3348_ (
    .A(\ALU.op [2]),
    .B(_1640_),
    .Y(_1643_)
);

AOI21X1 _3349_ (
    .A(_1639_),
    .B(_1643_),
    .C(_1642_),
    .Y(_1644_)
);

NAND2X1 _3350_ (
    .A(\ALU.BI7 ),
    .B(_1629__bF$buf3),
    .Y(_1645_)
);

OAI21X1 _3351_ (
    .A(_1629__bF$buf2),
    .B(_1644_),
    .C(_1645_),
    .Y(_1465_)
);

INVX1 _3352_ (
    .A(\ALU.CO ),
    .Y(_1646_)
);

OAI21X1 _3353_ (
    .A(_1642_),
    .B(_1643_),
    .C(_1639_),
    .Y(_1647_)
);

NAND2X1 _3354_ (
    .A(\ALU.right ),
    .B(AI[7]),
    .Y(_1648_)
);

AND2X2 _3355_ (
    .A(_1633_),
    .B(\ALU.BI [6]),
    .Y(_1649_)
);

NAND2X1 _3356_ (
    .A(AI[6]),
    .B(_1649_),
    .Y(_1650_)
);

AOI22X1 _3357_ (
    .A(_1631_),
    .B(\ALU.BI [6]),
    .C(_1650_),
    .D(_1632_),
    .Y(_1651_)
);

OAI21X1 _3358_ (
    .A(AI[6]),
    .B(_1649_),
    .C(_1637_),
    .Y(_1652_)
);

OAI21X1 _3359_ (
    .A(_1652_),
    .B(_1651_),
    .C(_1648_),
    .Y(_1653_)
);

NAND2X1 _3360_ (
    .A(\ALU.op [2]),
    .B(_1640_),
    .Y(_1654_)
);

INVX2 _3361_ (
    .A(\ALU.op [2]),
    .Y(_1655_)
);

OAI21X1 _3362_ (
    .A(\ALU.op [3]),
    .B(\ALU.BI [6]),
    .C(_1655_),
    .Y(_1656_)
);

OAI21X1 _3363_ (
    .A(\ALU.BI [6]),
    .B(_1654_),
    .C(_1656_),
    .Y(_1657_)
);

NAND2X1 _3364_ (
    .A(\ALU.right ),
    .B(AI[6]),
    .Y(_1658_)
);

AND2X2 _3365_ (
    .A(_1633_),
    .B(\ALU.BI [5]),
    .Y(_1659_)
);

NAND2X1 _3366_ (
    .A(AI[5]),
    .B(_1659_),
    .Y(_1660_)
);

AOI22X1 _3367_ (
    .A(_1631_),
    .B(\ALU.BI [5]),
    .C(_1660_),
    .D(_1632_),
    .Y(_1661_)
);

OAI21X1 _3368_ (
    .A(AI[5]),
    .B(_1659_),
    .C(_1637_),
    .Y(_1662_)
);

OAI21X1 _3369_ (
    .A(_1662_),
    .B(_1661_),
    .C(_1658_),
    .Y(_1663_)
);

OAI21X1 _3370_ (
    .A(\ALU.op [3]),
    .B(\ALU.BI [5]),
    .C(_1655_),
    .Y(_1664_)
);

OAI21X1 _3371_ (
    .A(\ALU.BI [5]),
    .B(_1654_),
    .C(_1664_),
    .Y(_1477_)
);

NAND2X1 _3372_ (
    .A(_1477_),
    .B(_1663_),
    .Y(_1478_)
);

NAND2X1 _3373_ (
    .A(\ALU.right ),
    .B(AI[5]),
    .Y(_1479_)
);

AND2X2 _3374_ (
    .A(_1633_),
    .B(\ALU.BI [4]),
    .Y(_1480_)
);

NAND2X1 _3375_ (
    .A(AI[4]),
    .B(_1480_),
    .Y(_1481_)
);

AOI22X1 _3376_ (
    .A(_1631_),
    .B(\ALU.BI [4]),
    .C(_1481_),
    .D(_1632_),
    .Y(_1482_)
);

OAI21X1 _3377_ (
    .A(AI[4]),
    .B(_1480_),
    .C(_1637_),
    .Y(_1483_)
);

OAI21X1 _3378_ (
    .A(_1483_),
    .B(_1482_),
    .C(_1479_),
    .Y(_1484_)
);

OAI21X1 _3379_ (
    .A(\ALU.op [3]),
    .B(\ALU.BI [4]),
    .C(_1655_),
    .Y(_1485_)
);

OAI21X1 _3380_ (
    .A(\ALU.BI [4]),
    .B(_1654_),
    .C(_1485_),
    .Y(_1486_)
);

NAND2X1 _3381_ (
    .A(\ALU.right ),
    .B(AI[4]),
    .Y(_1487_)
);

AND2X2 _3382_ (
    .A(_1633_),
    .B(\ALU.BI [3]),
    .Y(_1488_)
);

NAND2X1 _3383_ (
    .A(AI[3]),
    .B(_1488_),
    .Y(_1489_)
);

AOI22X1 _3384_ (
    .A(_1631_),
    .B(\ALU.BI [3]),
    .C(_1489_),
    .D(_1632_),
    .Y(_1490_)
);

OAI21X1 _3385_ (
    .A(AI[3]),
    .B(_1488_),
    .C(_1637_),
    .Y(_1491_)
);

OAI21X1 _3386_ (
    .A(_1491_),
    .B(_1490_),
    .C(_1487_),
    .Y(_1492_)
);

OAI21X1 _3387_ (
    .A(\ALU.op [3]),
    .B(\ALU.BI [3]),
    .C(_1655_),
    .Y(_1493_)
);

OAI21X1 _3388_ (
    .A(\ALU.BI [3]),
    .B(_1654_),
    .C(_1493_),
    .Y(_1494_)
);

NAND2X1 _3389_ (
    .A(_1494_),
    .B(_1492_),
    .Y(_1495_)
);

INVX1 _3390_ (
    .A(_1643_),
    .Y(_1496_)
);

AND2X2 _3391_ (
    .A(_1494_),
    .B(_1496_),
    .Y(_1497_)
);

OAI21X1 _3392_ (
    .A(_1492_),
    .B(_1497_),
    .C(_1495_),
    .Y(_1498_)
);

INVX1 _3393_ (
    .A(_1498_),
    .Y(_1499_)
);

NAND2X1 _3394_ (
    .A(AI[3]),
    .B(\ALU.right ),
    .Y(_1500_)
);

NAND3X1 _3395_ (
    .A(\ALU.BI [2]),
    .B(AI[2]),
    .C(_1633_),
    .Y(_1501_)
);

AOI22X1 _3396_ (
    .A(\ALU.BI [2]),
    .B(_1631_),
    .C(_1501_),
    .D(_1632_),
    .Y(_1502_)
);

INVX1 _3397_ (
    .A(\ALU.BI [2]),
    .Y(_1503_)
);

INVX1 _3398_ (
    .A(AI[2]),
    .Y(_1504_)
);

OAI21X1 _3399_ (
    .A(\ALU.op [0]),
    .B(_1503_),
    .C(_1504_),
    .Y(_1505_)
);

NAND2X1 _3400_ (
    .A(_1637_),
    .B(_1505_),
    .Y(_1506_)
);

OAI21X1 _3401_ (
    .A(_1506_),
    .B(_1502_),
    .C(_1500_),
    .Y(_1507_)
);

NOR2X1 _3402_ (
    .A(\ALU.BI [2]),
    .B(\ALU.op [3]),
    .Y(_1508_)
);

XOR2X1 _3403_ (
    .A(_1508_),
    .B(_1655_),
    .Y(_1509_)
);

NAND3X1 _3404_ (
    .A(\ALU.BI [1]),
    .B(AI[1]),
    .C(_1633_),
    .Y(_1510_)
);

AOI22X1 _3405_ (
    .A(_1631_),
    .B(\ALU.BI [1]),
    .C(_1510_),
    .D(_1632_),
    .Y(_1511_)
);

INVX1 _3406_ (
    .A(\ALU.BI [1]),
    .Y(_1512_)
);

NOR2X1 _3407_ (
    .A(\ALU.op [0]),
    .B(_1512_),
    .Y(_1513_)
);

OAI21X1 _3408_ (
    .A(AI[1]),
    .B(_1513_),
    .C(_1637_),
    .Y(_1514_)
);

OAI22X1 _3409_ (
    .A(_1504_),
    .B(_1637_),
    .C(_1511_),
    .D(_1514_),
    .Y(_1515_)
);

OAI21X1 _3410_ (
    .A(\ALU.op [2]),
    .B(\ALU.BI [1]),
    .C(_1640_),
    .Y(_1516_)
);

AOI21X1 _3411_ (
    .A(\ALU.op [2]),
    .B(\ALU.BI [1]),
    .C(_1516_),
    .Y(_1517_)
);

OAI21X1 _3412_ (
    .A(_1643_),
    .B(_1517_),
    .C(_1515_),
    .Y(_1518_)
);

NAND2X1 _3413_ (
    .A(\ALU.BI [0]),
    .B(_1633_),
    .Y(_1519_)
);

NAND2X1 _3414_ (
    .A(\ALU.op [1]),
    .B(AI[0]),
    .Y(_1520_)
);

AOI22X1 _3415_ (
    .A(\ALU.BI [0]),
    .B(_1520_),
    .C(_1632_),
    .D(_1519_),
    .Y(_1521_)
);

INVX1 _3416_ (
    .A(\ALU.BI [0]),
    .Y(_1522_)
);

INVX1 _3417_ (
    .A(AI[0]),
    .Y(_1523_)
);

OAI21X1 _3418_ (
    .A(\ALU.op [0]),
    .B(_1522_),
    .C(_1523_),
    .Y(_1524_)
);

NAND2X1 _3419_ (
    .A(_1637_),
    .B(_1524_),
    .Y(_1525_)
);

NAND2X1 _3420_ (
    .A(\ALU.right ),
    .B(AI[1]),
    .Y(_1526_)
);

OAI21X1 _3421_ (
    .A(_1521_),
    .B(_1525_),
    .C(_1526_),
    .Y(_1527_)
);

OAI21X1 _3422_ (
    .A(\ALU.op [2]),
    .B(\ALU.BI [0]),
    .C(_1640_),
    .Y(_1528_)
);

INVX1 _3423_ (
    .A(_1528_),
    .Y(_1529_)
);

OAI21X1 _3424_ (
    .A(_1655_),
    .B(_1522_),
    .C(_1529_),
    .Y(_1530_)
);

OAI21X1 _3425_ (
    .A(_1640_),
    .B(\ALU.op [2]),
    .C(_1530_),
    .Y(_1531_)
);

OAI21X1 _3426_ (
    .A(_1640_),
    .B(_1655_),
    .C(\ALU.CI ),
    .Y(_1532_)
);

NOR2X1 _3427_ (
    .A(\ALU.right ),
    .B(_1532_),
    .Y(_1533_)
);

MUX2X1 _3428_ (
    .A(\ALU.op [1]),
    .B(_1522_),
    .S(\ALU.op [0]),
    .Y(_1534_)
);

NAND2X1 _3429_ (
    .A(\ALU.BI [0]),
    .B(_1520_),
    .Y(_1535_)
);

NAND2X1 _3430_ (
    .A(_1535_),
    .B(_1534_),
    .Y(_1536_)
);

AOI21X1 _3431_ (
    .A(_1519_),
    .B(_1523_),
    .C(\ALU.right ),
    .Y(_1537_)
);

NAND2X1 _3432_ (
    .A(_1537_),
    .B(_1536_),
    .Y(_1538_)
);

NAND3X1 _3433_ (
    .A(_1526_),
    .B(_1530_),
    .C(_1538_),
    .Y(_1539_)
);

AOI22X1 _3434_ (
    .A(_1527_),
    .B(_1531_),
    .C(_1539_),
    .D(_1533_),
    .Y(_1540_)
);

NOR2X1 _3435_ (
    .A(_1517_),
    .B(_1515_),
    .Y(_1541_)
);

OAI21X1 _3436_ (
    .A(_1541_),
    .B(_1540_),
    .C(_1518_),
    .Y(_1542_)
);

NAND2X1 _3437_ (
    .A(_1509_),
    .B(_1507_),
    .Y(_1543_)
);

NAND2X1 _3438_ (
    .A(_1640_),
    .B(_1509_),
    .Y(_1544_)
);

INVX1 _3439_ (
    .A(_1544_),
    .Y(_1545_)
);

OAI21X1 _3440_ (
    .A(_1507_),
    .B(_1545_),
    .C(_1543_),
    .Y(_1546_)
);

INVX1 _3441_ (
    .A(_1546_),
    .Y(_1547_)
);

AOI22X1 _3442_ (
    .A(_1507_),
    .B(_1509_),
    .C(_1542_),
    .D(_1547_),
    .Y(_1548_)
);

XOR2X1 _3443_ (
    .A(_1548_),
    .B(_1499_),
    .Y(_1549_)
);

AOI21X1 _3444_ (
    .A(\ALU.op [2]),
    .B(\ALU.BI [0]),
    .C(_1528_),
    .Y(_1550_)
);

OAI21X1 _3445_ (
    .A(_1643_),
    .B(_1550_),
    .C(_1527_),
    .Y(_1551_)
);

INVX1 _3446_ (
    .A(_1533_),
    .Y(_1552_)
);

NOR2X1 _3447_ (
    .A(_1550_),
    .B(_1527_),
    .Y(_1553_)
);

OAI21X1 _3448_ (
    .A(_1552_),
    .B(_1553_),
    .C(_1551_),
    .Y(_1554_)
);

INVX1 _3449_ (
    .A(_1517_),
    .Y(_1555_)
);

OAI21X1 _3450_ (
    .A(_1640_),
    .B(\ALU.op [2]),
    .C(_1555_),
    .Y(_1556_)
);

MUX2X1 _3451_ (
    .A(_1556_),
    .B(_1555_),
    .S(_1515_),
    .Y(_1557_)
);

NAND2X1 _3452_ (
    .A(_1557_),
    .B(_1554_),
    .Y(_1558_)
);

OAI21X1 _3453_ (
    .A(_1515_),
    .B(_1517_),
    .C(_1518_),
    .Y(_1559_)
);

NAND2X1 _3454_ (
    .A(_1540_),
    .B(_1559_),
    .Y(_1560_)
);

NAND2X1 _3455_ (
    .A(_1560_),
    .B(_1558_),
    .Y(_1561_)
);

NAND2X1 _3456_ (
    .A(_1546_),
    .B(_1542_),
    .Y(_1562_)
);

NAND3X1 _3457_ (
    .A(_1518_),
    .B(_1547_),
    .C(_1558_),
    .Y(_1563_)
);

NAND3X1 _3458_ (
    .A(_1562_),
    .B(_1561_),
    .C(_1563_),
    .Y(_1564_)
);

NAND2X1 _3459_ (
    .A(\ALU.BCD ),
    .B(_1564_),
    .Y(_1565_)
);

OAI21X1 _3460_ (
    .A(_1498_),
    .B(_1548_),
    .C(_1495_),
    .Y(_1566_)
);

INVX1 _3461_ (
    .A(_1566_),
    .Y(_1567_)
);

OAI21X1 _3462_ (
    .A(_1565_),
    .B(_1549_),
    .C(_1567_),
    .Y(_1568_)
);

NAND2X1 _3463_ (
    .A(_1486_),
    .B(_1484_),
    .Y(_1569_)
);

OAI21X1 _3464_ (
    .A(_1640_),
    .B(\ALU.op [2]),
    .C(_1486_),
    .Y(_1570_)
);

INVX1 _3465_ (
    .A(_1570_),
    .Y(_1571_)
);

OAI21X1 _3466_ (
    .A(_1484_),
    .B(_1571_),
    .C(_1569_),
    .Y(_1572_)
);

INVX1 _3467_ (
    .A(_1572_),
    .Y(_1573_)
);

AOI22X1 _3468_ (
    .A(_1484_),
    .B(_1486_),
    .C(_1568_),
    .D(_1573_),
    .Y(_1574_)
);

OAI21X1 _3469_ (
    .A(_1640_),
    .B(\ALU.op [2]),
    .C(_1477_),
    .Y(_1575_)
);

INVX1 _3470_ (
    .A(_1575_),
    .Y(_1576_)
);

OAI21X1 _3471_ (
    .A(_1663_),
    .B(_1576_),
    .C(_1478_),
    .Y(_1577_)
);

OAI21X1 _3472_ (
    .A(_1577_),
    .B(_1574_),
    .C(_1478_),
    .Y(_1578_)
);

NAND2X1 _3473_ (
    .A(_1657_),
    .B(_1653_),
    .Y(_1579_)
);

OAI21X1 _3474_ (
    .A(_1640_),
    .B(\ALU.op [2]),
    .C(_1657_),
    .Y(_1580_)
);

INVX1 _3475_ (
    .A(_1580_),
    .Y(_1581_)
);

OAI21X1 _3476_ (
    .A(_1653_),
    .B(_1581_),
    .C(_1579_),
    .Y(_1582_)
);

INVX1 _3477_ (
    .A(_1582_),
    .Y(_1583_)
);

AOI22X1 _3478_ (
    .A(_1653_),
    .B(_1657_),
    .C(_1578_),
    .D(_1583_),
    .Y(_1584_)
);

OAI21X1 _3479_ (
    .A(_1639_),
    .B(_1642_),
    .C(_1647_),
    .Y(_1585_)
);

OAI21X1 _3480_ (
    .A(_1585_),
    .B(_1584_),
    .C(_1647_),
    .Y(_1586_)
);

NAND2X1 _3481_ (
    .A(\ALU.right ),
    .B(AI[0]),
    .Y(_1587_)
);

XOR2X1 _3482_ (
    .A(_1586_),
    .B(_1587_),
    .Y(_1588_)
);

XOR2X1 _3483_ (
    .A(_1584_),
    .B(_1585_),
    .Y(_1589_)
);

INVX1 _3484_ (
    .A(\ALU.BCD ),
    .Y(_1590_)
);

XOR2X1 _3485_ (
    .A(_1548_),
    .B(_1498_),
    .Y(_1591_)
);

XOR2X1 _3486_ (
    .A(_1542_),
    .B(_1546_),
    .Y(_1592_)
);

AOI21X1 _3487_ (
    .A(_1592_),
    .B(_1561_),
    .C(_1590_),
    .Y(_1593_)
);

AOI21X1 _3488_ (
    .A(_1593_),
    .B(_1591_),
    .C(_1566_),
    .Y(_1594_)
);

OAI21X1 _3489_ (
    .A(_1572_),
    .B(_1594_),
    .C(_1569_),
    .Y(_1595_)
);

INVX1 _3490_ (
    .A(_1577_),
    .Y(_1596_)
);

NAND2X1 _3491_ (
    .A(_1596_),
    .B(_1595_),
    .Y(_1597_)
);

NAND2X1 _3492_ (
    .A(_1577_),
    .B(_1574_),
    .Y(_1598_)
);

NAND2X1 _3493_ (
    .A(_1598_),
    .B(_1597_),
    .Y(_1599_)
);

NAND2X1 _3494_ (
    .A(_1583_),
    .B(_1578_),
    .Y(_1600_)
);

NAND3X1 _3495_ (
    .A(_1478_),
    .B(_1582_),
    .C(_1597_),
    .Y(_1601_)
);

NAND2X1 _3496_ (
    .A(_1601_),
    .B(_1600_),
    .Y(_1602_)
);

AOI21X1 _3497_ (
    .A(_1602_),
    .B(_1599_),
    .C(_1590_),
    .Y(_1603_)
);

AOI21X1 _3498_ (
    .A(_1589_),
    .B(_1603_),
    .C(_1629__bF$buf1),
    .Y(_1604_)
);

AOI22X1 _3499_ (
    .A(_1646_),
    .B(_1629__bF$buf0),
    .C(_1604_),
    .D(_1588_),
    .Y(_1466_)
);

NAND2X1 _3500_ (
    .A(\ALU.HC ),
    .B(_1629__bF$buf3),
    .Y(_1605_)
);

OAI21X1 _3501_ (
    .A(_1629__bF$buf2),
    .B(_1594_),
    .C(_1605_),
    .Y(_1467_)
);

NAND2X1 _3502_ (
    .A(ADD[0]),
    .B(_1629__bF$buf1),
    .Y(_1606_)
);

AOI21X1 _3503_ (
    .A(_1551_),
    .B(_1539_),
    .C(_1533_),
    .Y(_1607_)
);

OAI21X1 _3504_ (
    .A(_1527_),
    .B(_1550_),
    .C(_1551_),
    .Y(_1608_)
);

OAI21X1 _3505_ (
    .A(_1552_),
    .B(_1608_),
    .C(RDY_bF$buf5),
    .Y(_1609_)
);

OAI21X1 _3506_ (
    .A(_1607_),
    .B(_1609_),
    .C(_1606_),
    .Y(_1468_)
);

NAND2X1 _3507_ (
    .A(ADD[1]),
    .B(_1629__bF$buf0),
    .Y(_1610_)
);

OAI21X1 _3508_ (
    .A(_1629__bF$buf3),
    .B(_1561_),
    .C(_1610_),
    .Y(_1469_)
);

NAND2X1 _3509_ (
    .A(ADD[2]),
    .B(_1629__bF$buf2),
    .Y(_1611_)
);

OAI21X1 _3510_ (
    .A(_1629__bF$buf1),
    .B(_1592_),
    .C(_1611_),
    .Y(_1470_)
);

NAND2X1 _3511_ (
    .A(ADD[3]),
    .B(_1629__bF$buf0),
    .Y(_1612_)
);

OAI21X1 _3512_ (
    .A(_1629__bF$buf3),
    .B(_1549_),
    .C(_1612_),
    .Y(_1471_)
);

NAND2X1 _3513_ (
    .A(ADD[4]),
    .B(_1629__bF$buf2),
    .Y(_1613_)
);

NOR2X1 _3514_ (
    .A(_1573_),
    .B(_1568_),
    .Y(_1614_)
);

OAI21X1 _3515_ (
    .A(_1572_),
    .B(_1594_),
    .C(RDY_bF$buf4),
    .Y(_1615_)
);

OAI21X1 _3516_ (
    .A(_1614_),
    .B(_1615_),
    .C(_1613_),
    .Y(_1472_)
);

NAND2X1 _3517_ (
    .A(ADD[5]),
    .B(_1629__bF$buf1),
    .Y(_1616_)
);

OAI21X1 _3518_ (
    .A(_1629__bF$buf0),
    .B(_1599_),
    .C(_1616_),
    .Y(_1473_)
);

NAND2X1 _3519_ (
    .A(ADD[6]),
    .B(_1629__bF$buf3),
    .Y(_1617_)
);

OAI21X1 _3520_ (
    .A(_1629__bF$buf2),
    .B(_1602_),
    .C(_1617_),
    .Y(_1474_)
);

INVX1 _3521_ (
    .A(\ALU.N ),
    .Y(_1618_)
);

NAND2X1 _3522_ (
    .A(RDY_bF$buf3),
    .B(_1589_),
    .Y(_1619_)
);

OAI21X1 _3523_ (
    .A(_1618_),
    .B(RDY_bF$buf2),
    .C(_1619_),
    .Y(_1475_)
);

INVX1 _3524_ (
    .A(\ALU.AI7 ),
    .Y(_1620_)
);

NAND2X1 _3525_ (
    .A(AI[7]),
    .B(RDY_bF$buf1),
    .Y(_1621_)
);

OAI21X1 _3526_ (
    .A(RDY_bF$buf0),
    .B(_1620_),
    .C(_1621_),
    .Y(_1476_)
);

DFFSR _3527_ (
    .CLK(clk_bF$buf0),
    .D(_1465_),
    .Q(\ALU.BI7 ),
    .R(_1464_),
    .S(vdd)
);

DFFSR _3528_ (
    .CLK(clk_bF$buf10),
    .D(_1466_),
    .Q(\ALU.CO ),
    .R(_1464_),
    .S(vdd)
);

DFFSR _3529_ (
    .CLK(clk_bF$buf9),
    .D(_1467_),
    .Q(\ALU.HC ),
    .R(_1464_),
    .S(vdd)
);

DFFSR _3530_ (
    .CLK(clk_bF$buf8),
    .D(_1468_),
    .Q(ADD[0]),
    .R(_1464_),
    .S(vdd)
);

DFFSR _3531_ (
    .CLK(clk_bF$buf7),
    .D(_1469_),
    .Q(ADD[1]),
    .R(_1464_),
    .S(vdd)
);

DFFSR _3532_ (
    .CLK(clk_bF$buf6),
    .D(_1470_),
    .Q(ADD[2]),
    .R(_1464_),
    .S(vdd)
);

DFFSR _3533_ (
    .CLK(clk_bF$buf5),
    .D(_1471_),
    .Q(ADD[3]),
    .R(_1464_),
    .S(vdd)
);

DFFSR _3534_ (
    .CLK(clk_bF$buf4),
    .D(_1472_),
    .Q(ADD[4]),
    .R(_1464_),
    .S(vdd)
);

DFFSR _3535_ (
    .CLK(clk_bF$buf3),
    .D(_1473_),
    .Q(ADD[5]),
    .R(_1464_),
    .S(vdd)
);

DFFSR _3536_ (
    .CLK(clk_bF$buf2),
    .D(_1474_),
    .Q(ADD[6]),
    .R(_1464_),
    .S(vdd)
);

DFFSR _3537_ (
    .CLK(clk_bF$buf1),
    .D(_1475_),
    .Q(\ALU.N ),
    .R(_1464_),
    .S(vdd)
);

DFFSR _3538_ (
    .CLK(clk_bF$buf0),
    .D(_1476_),
    .Q(\ALU.AI7 ),
    .R(_1464_),
    .S(vdd)
);

BUFX2 _3539_ (
    .A(_1665_[0]),
    .Y(AB[0])
);

BUFX2 _3540_ (
    .A(_1665_[1]),
    .Y(AB[1])
);

BUFX2 _3541_ (
    .A(_1665_[10]),
    .Y(AB[10])
);

BUFX2 _3542_ (
    .A(_1665_[11]),
    .Y(AB[11])
);

BUFX2 _3543_ (
    .A(_1665_[12]),
    .Y(AB[12])
);

BUFX2 _3544_ (
    .A(_1665_[13]),
    .Y(AB[13])
);

BUFX2 _3545_ (
    .A(_1665_[14]),
    .Y(AB[14])
);

BUFX2 _3546_ (
    .A(_1665_[15]),
    .Y(AB[15])
);

BUFX2 _3547_ (
    .A(_1665_[2]),
    .Y(AB[2])
);

BUFX2 _3548_ (
    .A(_1665_[3]),
    .Y(AB[3])
);

BUFX2 _3549_ (
    .A(_1665_[4]),
    .Y(AB[4])
);

BUFX2 _3550_ (
    .A(_1665_[5]),
    .Y(AB[5])
);

BUFX2 _3551_ (
    .A(_1665_[6]),
    .Y(AB[6])
);

BUFX2 _3552_ (
    .A(_1665_[7]),
    .Y(AB[7])
);

BUFX2 _3553_ (
    .A(_1665_[8]),
    .Y(AB[8])
);

BUFX2 _3554_ (
    .A(_1665_[9]),
    .Y(AB[9])
);

BUFX2 _3555_ (
    .A(_1666_[0]),
    .Y(DO[0])
);

BUFX2 _3556_ (
    .A(_1666_[1]),
    .Y(DO[1])
);

BUFX2 _3557_ (
    .A(_1666_[2]),
    .Y(DO[2])
);

BUFX2 _3558_ (
    .A(_1666_[3]),
    .Y(DO[3])
);

BUFX2 _3559_ (
    .A(_1666_[4]),
    .Y(DO[4])
);

BUFX2 _3560_ (
    .A(_1666_[5]),
    .Y(DO[5])
);

BUFX2 _3561_ (
    .A(_1666_[6]),
    .Y(DO[6])
);

BUFX2 _3562_ (
    .A(_1666_[7]),
    .Y(DO[7])
);

BUFX2 _3563_ (
    .A(_1667_),
    .Y(WE)
);

endmodule

magic
tech scmos
magscale 1 30
timestamp 1715930203
<< checkpaint >>
rect -600 -600 380600 380600
<< metal1 >>
rect 106550 280415 113150 280550
rect 106550 280325 106655 280415
rect 106745 280325 106835 280415
rect 106925 280325 107015 280415
rect 107105 280325 107195 280415
rect 107285 280325 107375 280415
rect 107465 280325 107555 280415
rect 107645 280325 107735 280415
rect 107825 280325 107915 280415
rect 108005 280325 108095 280415
rect 108185 280325 108275 280415
rect 108365 280325 108455 280415
rect 108545 280325 108635 280415
rect 108725 280325 108815 280415
rect 108905 280325 108995 280415
rect 109085 280325 109175 280415
rect 109265 280325 109355 280415
rect 109445 280325 109535 280415
rect 109625 280325 109715 280415
rect 109805 280325 109895 280415
rect 109985 280325 110075 280415
rect 110165 280325 110255 280415
rect 110345 280325 110435 280415
rect 110525 280325 110615 280415
rect 110705 280325 110795 280415
rect 110885 280325 110975 280415
rect 111065 280325 111155 280415
rect 111245 280325 111335 280415
rect 111425 280325 111515 280415
rect 111605 280325 111695 280415
rect 111785 280325 111875 280415
rect 111965 280325 112055 280415
rect 112145 280325 112235 280415
rect 112325 280325 112415 280415
rect 112505 280325 112595 280415
rect 112685 280325 112775 280415
rect 112865 280325 112955 280415
rect 113045 280325 113150 280415
rect 106550 280235 113150 280325
rect 106550 280145 106655 280235
rect 106745 280145 106835 280235
rect 106925 280145 107015 280235
rect 107105 280145 107195 280235
rect 107285 280145 107375 280235
rect 107465 280145 107555 280235
rect 107645 280145 107735 280235
rect 107825 280145 107915 280235
rect 108005 280145 108095 280235
rect 108185 280145 108275 280235
rect 108365 280145 108455 280235
rect 108545 280145 108635 280235
rect 108725 280145 108815 280235
rect 108905 280145 108995 280235
rect 109085 280145 109175 280235
rect 109265 280145 109355 280235
rect 109445 280145 109535 280235
rect 109625 280145 109715 280235
rect 109805 280145 109895 280235
rect 109985 280145 110075 280235
rect 110165 280145 110255 280235
rect 110345 280145 110435 280235
rect 110525 280145 110615 280235
rect 110705 280145 110795 280235
rect 110885 280145 110975 280235
rect 111065 280145 111155 280235
rect 111245 280145 111335 280235
rect 111425 280145 111515 280235
rect 111605 280145 111695 280235
rect 111785 280145 111875 280235
rect 111965 280145 112055 280235
rect 112145 280145 112235 280235
rect 112325 280145 112415 280235
rect 112505 280145 112595 280235
rect 112685 280145 112775 280235
rect 112865 280145 112955 280235
rect 113045 280145 113150 280235
rect 106550 280055 113150 280145
rect 106550 279965 106655 280055
rect 106745 279965 106835 280055
rect 106925 279965 107015 280055
rect 107105 279965 107195 280055
rect 107285 279965 107375 280055
rect 107465 279965 107555 280055
rect 107645 279965 107735 280055
rect 107825 279965 107915 280055
rect 108005 279965 108095 280055
rect 108185 279965 108275 280055
rect 108365 279965 108455 280055
rect 108545 279965 108635 280055
rect 108725 279965 108815 280055
rect 108905 279965 108995 280055
rect 109085 279965 109175 280055
rect 109265 279965 109355 280055
rect 109445 279965 109535 280055
rect 109625 279965 109715 280055
rect 109805 279965 109895 280055
rect 109985 279965 110075 280055
rect 110165 279965 110255 280055
rect 110345 279965 110435 280055
rect 110525 279965 110615 280055
rect 110705 279965 110795 280055
rect 110885 279965 110975 280055
rect 111065 279965 111155 280055
rect 111245 279965 111335 280055
rect 111425 279965 111515 280055
rect 111605 279965 111695 280055
rect 111785 279965 111875 280055
rect 111965 279965 112055 280055
rect 112145 279965 112235 280055
rect 112325 279965 112415 280055
rect 112505 279965 112595 280055
rect 112685 279965 112775 280055
rect 112865 279965 112955 280055
rect 113045 279965 113150 280055
rect 106550 279875 113150 279965
rect 106550 279785 106655 279875
rect 106745 279785 106835 279875
rect 106925 279785 107015 279875
rect 107105 279785 107195 279875
rect 107285 279785 107375 279875
rect 107465 279785 107555 279875
rect 107645 279785 107735 279875
rect 107825 279785 107915 279875
rect 108005 279785 108095 279875
rect 108185 279785 108275 279875
rect 108365 279785 108455 279875
rect 108545 279785 108635 279875
rect 108725 279785 108815 279875
rect 108905 279785 108995 279875
rect 109085 279785 109175 279875
rect 109265 279785 109355 279875
rect 109445 279785 109535 279875
rect 109625 279785 109715 279875
rect 109805 279785 109895 279875
rect 109985 279785 110075 279875
rect 110165 279785 110255 279875
rect 110345 279785 110435 279875
rect 110525 279785 110615 279875
rect 110705 279785 110795 279875
rect 110885 279785 110975 279875
rect 111065 279785 111155 279875
rect 111245 279785 111335 279875
rect 111425 279785 111515 279875
rect 111605 279785 111695 279875
rect 111785 279785 111875 279875
rect 111965 279785 112055 279875
rect 112145 279785 112235 279875
rect 112325 279785 112415 279875
rect 112505 279785 112595 279875
rect 112685 279785 112775 279875
rect 112865 279785 112955 279875
rect 113045 279785 113150 279875
rect 106550 279650 113150 279785
rect 104300 278850 113150 279650
rect 265350 280445 274450 280550
rect 265350 280355 265445 280445
rect 265535 280355 265625 280445
rect 265715 280355 265805 280445
rect 265895 280355 265985 280445
rect 266075 280355 266165 280445
rect 266255 280355 266345 280445
rect 266435 280355 266525 280445
rect 266615 280355 266705 280445
rect 266795 280355 266885 280445
rect 266975 280355 267065 280445
rect 267155 280355 267245 280445
rect 267335 280355 267425 280445
rect 267515 280355 267605 280445
rect 267695 280355 267785 280445
rect 267875 280355 267965 280445
rect 268055 280355 268145 280445
rect 268235 280355 268325 280445
rect 268415 280355 268505 280445
rect 268595 280355 268685 280445
rect 268775 280355 268865 280445
rect 268955 280355 269045 280445
rect 269135 280355 269225 280445
rect 269315 280355 269405 280445
rect 269495 280355 269585 280445
rect 269675 280355 269765 280445
rect 269855 280355 269945 280445
rect 270035 280355 270125 280445
rect 270215 280355 270305 280445
rect 270395 280355 270485 280445
rect 270575 280355 270665 280445
rect 270755 280355 270845 280445
rect 270935 280355 271025 280445
rect 271115 280355 271205 280445
rect 271295 280355 271385 280445
rect 271475 280355 271565 280445
rect 271655 280355 271745 280445
rect 271835 280355 271925 280445
rect 272015 280355 272105 280445
rect 272195 280355 272285 280445
rect 272375 280355 272465 280445
rect 272555 280355 272645 280445
rect 272735 280355 272825 280445
rect 272915 280355 273005 280445
rect 273095 280355 273185 280445
rect 273275 280355 273365 280445
rect 273455 280355 273545 280445
rect 273635 280355 273725 280445
rect 273815 280355 273905 280445
rect 273995 280355 274085 280445
rect 274175 280355 274265 280445
rect 274355 280355 274450 280445
rect 265350 280265 274450 280355
rect 265350 280175 265445 280265
rect 265535 280175 265625 280265
rect 265715 280175 265805 280265
rect 265895 280175 265985 280265
rect 266075 280175 266165 280265
rect 266255 280175 266345 280265
rect 266435 280175 266525 280265
rect 266615 280175 266705 280265
rect 266795 280175 266885 280265
rect 266975 280175 267065 280265
rect 267155 280175 267245 280265
rect 267335 280175 267425 280265
rect 267515 280175 267605 280265
rect 267695 280175 267785 280265
rect 267875 280175 267965 280265
rect 268055 280175 268145 280265
rect 268235 280175 268325 280265
rect 268415 280175 268505 280265
rect 268595 280175 268685 280265
rect 268775 280175 268865 280265
rect 268955 280175 269045 280265
rect 269135 280175 269225 280265
rect 269315 280175 269405 280265
rect 269495 280175 269585 280265
rect 269675 280175 269765 280265
rect 269855 280175 269945 280265
rect 270035 280175 270125 280265
rect 270215 280175 270305 280265
rect 270395 280175 270485 280265
rect 270575 280175 270665 280265
rect 270755 280175 270845 280265
rect 270935 280175 271025 280265
rect 271115 280175 271205 280265
rect 271295 280175 271385 280265
rect 271475 280175 271565 280265
rect 271655 280175 271745 280265
rect 271835 280175 271925 280265
rect 272015 280175 272105 280265
rect 272195 280175 272285 280265
rect 272375 280175 272465 280265
rect 272555 280175 272645 280265
rect 272735 280175 272825 280265
rect 272915 280175 273005 280265
rect 273095 280175 273185 280265
rect 273275 280175 273365 280265
rect 273455 280175 273545 280265
rect 273635 280175 273725 280265
rect 273815 280175 273905 280265
rect 273995 280175 274085 280265
rect 274175 280175 274265 280265
rect 274355 280175 274450 280265
rect 265350 280085 274450 280175
rect 265350 279995 265445 280085
rect 265535 279995 265625 280085
rect 265715 279995 265805 280085
rect 265895 279995 265985 280085
rect 266075 279995 266165 280085
rect 266255 279995 266345 280085
rect 266435 279995 266525 280085
rect 266615 279995 266705 280085
rect 266795 279995 266885 280085
rect 266975 279995 267065 280085
rect 267155 279995 267245 280085
rect 267335 279995 267425 280085
rect 267515 279995 267605 280085
rect 267695 279995 267785 280085
rect 267875 279995 267965 280085
rect 268055 279995 268145 280085
rect 268235 279995 268325 280085
rect 268415 279995 268505 280085
rect 268595 279995 268685 280085
rect 268775 279995 268865 280085
rect 268955 279995 269045 280085
rect 269135 279995 269225 280085
rect 269315 279995 269405 280085
rect 269495 279995 269585 280085
rect 269675 279995 269765 280085
rect 269855 279995 269945 280085
rect 270035 279995 270125 280085
rect 270215 279995 270305 280085
rect 270395 279995 270485 280085
rect 270575 279995 270665 280085
rect 270755 279995 270845 280085
rect 270935 279995 271025 280085
rect 271115 279995 271205 280085
rect 271295 279995 271385 280085
rect 271475 279995 271565 280085
rect 271655 279995 271745 280085
rect 271835 279995 271925 280085
rect 272015 279995 272105 280085
rect 272195 279995 272285 280085
rect 272375 279995 272465 280085
rect 272555 279995 272645 280085
rect 272735 279995 272825 280085
rect 272915 279995 273005 280085
rect 273095 279995 273185 280085
rect 273275 279995 273365 280085
rect 273455 279995 273545 280085
rect 273635 279995 273725 280085
rect 273815 279995 273905 280085
rect 273995 279995 274085 280085
rect 274175 279995 274265 280085
rect 274355 279995 274450 280085
rect 265350 279905 274450 279995
rect 265350 279815 265445 279905
rect 265535 279815 265625 279905
rect 265715 279815 265805 279905
rect 265895 279815 265985 279905
rect 266075 279815 266165 279905
rect 266255 279815 266345 279905
rect 266435 279815 266525 279905
rect 266615 279815 266705 279905
rect 266795 279815 266885 279905
rect 266975 279815 267065 279905
rect 267155 279815 267245 279905
rect 267335 279815 267425 279905
rect 267515 279815 267605 279905
rect 267695 279815 267785 279905
rect 267875 279815 267965 279905
rect 268055 279815 268145 279905
rect 268235 279815 268325 279905
rect 268415 279815 268505 279905
rect 268595 279815 268685 279905
rect 268775 279815 268865 279905
rect 268955 279815 269045 279905
rect 269135 279815 269225 279905
rect 269315 279815 269405 279905
rect 269495 279815 269585 279905
rect 269675 279815 269765 279905
rect 269855 279815 269945 279905
rect 270035 279815 270125 279905
rect 270215 279815 270305 279905
rect 270395 279815 270485 279905
rect 270575 279815 270665 279905
rect 270755 279815 270845 279905
rect 270935 279815 271025 279905
rect 271115 279815 271205 279905
rect 271295 279815 271385 279905
rect 271475 279815 271565 279905
rect 271655 279815 271745 279905
rect 271835 279815 271925 279905
rect 272015 279815 272105 279905
rect 272195 279815 272285 279905
rect 272375 279815 272465 279905
rect 272555 279815 272645 279905
rect 272735 279815 272825 279905
rect 272915 279815 273005 279905
rect 273095 279815 273185 279905
rect 273275 279815 273365 279905
rect 273455 279815 273545 279905
rect 273635 279815 273725 279905
rect 273815 279815 273905 279905
rect 273995 279815 274085 279905
rect 274175 279815 274265 279905
rect 274355 279815 274450 279905
rect 265350 279725 274450 279815
rect 265350 279635 265445 279725
rect 265535 279635 265625 279725
rect 265715 279635 265805 279725
rect 265895 279635 265985 279725
rect 266075 279635 266165 279725
rect 266255 279635 266345 279725
rect 266435 279635 266525 279725
rect 266615 279635 266705 279725
rect 266795 279635 266885 279725
rect 266975 279635 267065 279725
rect 267155 279635 267245 279725
rect 267335 279635 267425 279725
rect 267515 279635 267605 279725
rect 267695 279635 267785 279725
rect 267875 279635 267965 279725
rect 268055 279635 268145 279725
rect 268235 279635 268325 279725
rect 268415 279635 268505 279725
rect 268595 279635 268685 279725
rect 268775 279635 268865 279725
rect 268955 279635 269045 279725
rect 269135 279635 269225 279725
rect 269315 279635 269405 279725
rect 269495 279635 269585 279725
rect 269675 279635 269765 279725
rect 269855 279635 269945 279725
rect 270035 279635 270125 279725
rect 270215 279635 270305 279725
rect 270395 279635 270485 279725
rect 270575 279635 270665 279725
rect 270755 279635 270845 279725
rect 270935 279635 271025 279725
rect 271115 279635 271205 279725
rect 271295 279635 271385 279725
rect 271475 279635 271565 279725
rect 271655 279635 271745 279725
rect 271835 279635 271925 279725
rect 272015 279635 272105 279725
rect 272195 279635 272285 279725
rect 272375 279635 272465 279725
rect 272555 279635 272645 279725
rect 272735 279635 272825 279725
rect 272915 279635 273005 279725
rect 273095 279635 273185 279725
rect 273275 279635 273365 279725
rect 273455 279635 273545 279725
rect 273635 279635 273725 279725
rect 273815 279635 273905 279725
rect 273995 279635 274085 279725
rect 274175 279635 274265 279725
rect 274355 279635 274450 279725
rect 265350 279545 274450 279635
rect 265350 279455 265445 279545
rect 265535 279455 265625 279545
rect 265715 279455 265805 279545
rect 265895 279455 265985 279545
rect 266075 279455 266165 279545
rect 266255 279455 266345 279545
rect 266435 279455 266525 279545
rect 266615 279455 266705 279545
rect 266795 279455 266885 279545
rect 266975 279455 267065 279545
rect 267155 279455 267245 279545
rect 267335 279455 267425 279545
rect 267515 279455 267605 279545
rect 267695 279455 267785 279545
rect 267875 279455 267965 279545
rect 268055 279455 268145 279545
rect 268235 279455 268325 279545
rect 268415 279455 268505 279545
rect 268595 279455 268685 279545
rect 268775 279455 268865 279545
rect 268955 279455 269045 279545
rect 269135 279455 269225 279545
rect 269315 279455 269405 279545
rect 269495 279455 269585 279545
rect 269675 279455 269765 279545
rect 269855 279455 269945 279545
rect 270035 279455 270125 279545
rect 270215 279455 270305 279545
rect 270395 279455 270485 279545
rect 270575 279455 270665 279545
rect 270755 279455 270845 279545
rect 270935 279455 271025 279545
rect 271115 279455 271205 279545
rect 271295 279455 271385 279545
rect 271475 279455 271565 279545
rect 271655 279455 271745 279545
rect 271835 279455 271925 279545
rect 272015 279455 272105 279545
rect 272195 279455 272285 279545
rect 272375 279455 272465 279545
rect 272555 279455 272645 279545
rect 272735 279455 272825 279545
rect 272915 279455 273005 279545
rect 273095 279455 273185 279545
rect 273275 279455 273365 279545
rect 273455 279455 273545 279545
rect 273635 279455 273725 279545
rect 273815 279455 273905 279545
rect 273995 279455 274085 279545
rect 274175 279455 274265 279545
rect 274355 279455 274450 279545
rect 265350 279350 274450 279455
rect 104300 269630 105200 278850
rect 265350 278150 276290 279350
rect 275390 269030 276290 278150
rect 104250 189850 104650 190650
rect 104300 100950 105200 103550
rect 275390 101450 276290 103619
rect 104298 100355 113150 100950
rect 104298 100350 106655 100355
rect 106550 100265 106655 100350
rect 106745 100265 106835 100355
rect 106925 100265 107015 100355
rect 107105 100265 107195 100355
rect 107285 100265 107375 100355
rect 107465 100265 107555 100355
rect 107645 100265 107735 100355
rect 107825 100265 107915 100355
rect 108005 100265 108095 100355
rect 108185 100265 108275 100355
rect 108365 100265 108455 100355
rect 108545 100265 108635 100355
rect 108725 100265 108815 100355
rect 108905 100265 108995 100355
rect 109085 100265 109175 100355
rect 109265 100265 109355 100355
rect 109445 100265 109535 100355
rect 109625 100265 109715 100355
rect 109805 100265 109895 100355
rect 109985 100265 110075 100355
rect 110165 100265 110255 100355
rect 110345 100265 110435 100355
rect 110525 100265 110615 100355
rect 110705 100265 110795 100355
rect 110885 100265 110975 100355
rect 111065 100265 111155 100355
rect 111245 100265 111335 100355
rect 111425 100265 111515 100355
rect 111605 100265 111695 100355
rect 111785 100265 111875 100355
rect 111965 100265 112055 100355
rect 112145 100265 112235 100355
rect 112325 100265 112415 100355
rect 112505 100265 112595 100355
rect 112685 100265 112775 100355
rect 112865 100265 112955 100355
rect 113045 100265 113150 100355
rect 106550 100175 113150 100265
rect 106550 100085 106655 100175
rect 106745 100085 106835 100175
rect 106925 100085 107015 100175
rect 107105 100085 107195 100175
rect 107285 100085 107375 100175
rect 107465 100085 107555 100175
rect 107645 100085 107735 100175
rect 107825 100085 107915 100175
rect 108005 100085 108095 100175
rect 108185 100085 108275 100175
rect 108365 100085 108455 100175
rect 108545 100085 108635 100175
rect 108725 100085 108815 100175
rect 108905 100085 108995 100175
rect 109085 100085 109175 100175
rect 109265 100085 109355 100175
rect 109445 100085 109535 100175
rect 109625 100085 109715 100175
rect 109805 100085 109895 100175
rect 109985 100085 110075 100175
rect 110165 100085 110255 100175
rect 110345 100085 110435 100175
rect 110525 100085 110615 100175
rect 110705 100085 110795 100175
rect 110885 100085 110975 100175
rect 111065 100085 111155 100175
rect 111245 100085 111335 100175
rect 111425 100085 111515 100175
rect 111605 100085 111695 100175
rect 111785 100085 111875 100175
rect 111965 100085 112055 100175
rect 112145 100085 112235 100175
rect 112325 100085 112415 100175
rect 112505 100085 112595 100175
rect 112685 100085 112775 100175
rect 112865 100085 112955 100175
rect 113045 100085 113150 100175
rect 106550 99995 113150 100085
rect 106550 99905 106655 99995
rect 106745 99905 106835 99995
rect 106925 99905 107015 99995
rect 107105 99905 107195 99995
rect 107285 99905 107375 99995
rect 107465 99905 107555 99995
rect 107645 99905 107735 99995
rect 107825 99905 107915 99995
rect 108005 99905 108095 99995
rect 108185 99905 108275 99995
rect 108365 99905 108455 99995
rect 108545 99905 108635 99995
rect 108725 99905 108815 99995
rect 108905 99905 108995 99995
rect 109085 99905 109175 99995
rect 109265 99905 109355 99995
rect 109445 99905 109535 99995
rect 109625 99905 109715 99995
rect 109805 99905 109895 99995
rect 109985 99905 110075 99995
rect 110165 99905 110255 99995
rect 110345 99905 110435 99995
rect 110525 99905 110615 99995
rect 110705 99905 110795 99995
rect 110885 99905 110975 99995
rect 111065 99905 111155 99995
rect 111245 99905 111335 99995
rect 111425 99905 111515 99995
rect 111605 99905 111695 99995
rect 111785 99905 111875 99995
rect 111965 99905 112055 99995
rect 112145 99905 112235 99995
rect 112325 99905 112415 99995
rect 112505 99905 112595 99995
rect 112685 99905 112775 99995
rect 112865 99905 112955 99995
rect 113045 99905 113150 99995
rect 106550 99815 113150 99905
rect 106550 99725 106655 99815
rect 106745 99725 106835 99815
rect 106925 99725 107015 99815
rect 107105 99725 107195 99815
rect 107285 99725 107375 99815
rect 107465 99725 107555 99815
rect 107645 99725 107735 99815
rect 107825 99725 107915 99815
rect 108005 99725 108095 99815
rect 108185 99725 108275 99815
rect 108365 99725 108455 99815
rect 108545 99725 108635 99815
rect 108725 99725 108815 99815
rect 108905 99725 108995 99815
rect 109085 99725 109175 99815
rect 109265 99725 109355 99815
rect 109445 99725 109535 99815
rect 109625 99725 109715 99815
rect 109805 99725 109895 99815
rect 109985 99725 110075 99815
rect 110165 99725 110255 99815
rect 110345 99725 110435 99815
rect 110525 99725 110615 99815
rect 110705 99725 110795 99815
rect 110885 99725 110975 99815
rect 111065 99725 111155 99815
rect 111245 99725 111335 99815
rect 111425 99725 111515 99815
rect 111605 99725 111695 99815
rect 111785 99725 111875 99815
rect 111965 99725 112055 99815
rect 112145 99725 112235 99815
rect 112325 99725 112415 99815
rect 112505 99725 112595 99815
rect 112685 99725 112775 99815
rect 112865 99725 112955 99815
rect 113045 99725 113150 99815
rect 106550 99635 113150 99725
rect 106550 99545 106655 99635
rect 106745 99545 106835 99635
rect 106925 99545 107015 99635
rect 107105 99545 107195 99635
rect 107285 99545 107375 99635
rect 107465 99545 107555 99635
rect 107645 99545 107735 99635
rect 107825 99545 107915 99635
rect 108005 99545 108095 99635
rect 108185 99545 108275 99635
rect 108365 99545 108455 99635
rect 108545 99545 108635 99635
rect 108725 99545 108815 99635
rect 108905 99545 108995 99635
rect 109085 99545 109175 99635
rect 109265 99545 109355 99635
rect 109445 99545 109535 99635
rect 109625 99545 109715 99635
rect 109805 99545 109895 99635
rect 109985 99545 110075 99635
rect 110165 99545 110255 99635
rect 110345 99545 110435 99635
rect 110525 99545 110615 99635
rect 110705 99545 110795 99635
rect 110885 99545 110975 99635
rect 111065 99545 111155 99635
rect 111245 99545 111335 99635
rect 111425 99545 111515 99635
rect 111605 99545 111695 99635
rect 111785 99545 111875 99635
rect 111965 99545 112055 99635
rect 112145 99545 112235 99635
rect 112325 99545 112415 99635
rect 112505 99545 112595 99635
rect 112685 99545 112775 99635
rect 112865 99545 112955 99635
rect 113045 99545 113150 99635
rect 106550 99441 113150 99545
rect 265350 100450 276290 101450
rect 265350 100305 274450 100450
rect 265350 100215 265445 100305
rect 265535 100215 265625 100305
rect 265715 100215 265805 100305
rect 265895 100215 265985 100305
rect 266075 100215 266165 100305
rect 266255 100215 266345 100305
rect 266435 100215 266525 100305
rect 266615 100215 266705 100305
rect 266795 100215 266885 100305
rect 266975 100215 267065 100305
rect 267155 100215 267245 100305
rect 267335 100215 267425 100305
rect 267515 100215 267605 100305
rect 267695 100215 267785 100305
rect 267875 100215 267965 100305
rect 268055 100215 268145 100305
rect 268235 100215 268325 100305
rect 268415 100215 268505 100305
rect 268595 100215 268685 100305
rect 268775 100215 268865 100305
rect 268955 100215 269045 100305
rect 269135 100215 269225 100305
rect 269315 100215 269405 100305
rect 269495 100215 269585 100305
rect 269675 100215 269765 100305
rect 269855 100215 269945 100305
rect 270035 100215 270125 100305
rect 270215 100215 270305 100305
rect 270395 100215 270485 100305
rect 270575 100215 270665 100305
rect 270755 100215 270845 100305
rect 270935 100215 271025 100305
rect 271115 100215 271205 100305
rect 271295 100215 271385 100305
rect 271475 100215 271565 100305
rect 271655 100215 271745 100305
rect 271835 100215 271925 100305
rect 272015 100215 272105 100305
rect 272195 100215 272285 100305
rect 272375 100215 272465 100305
rect 272555 100215 272645 100305
rect 272735 100215 272825 100305
rect 272915 100215 273005 100305
rect 273095 100215 273185 100305
rect 273275 100215 273365 100305
rect 273455 100215 273545 100305
rect 273635 100215 273725 100305
rect 273815 100215 273905 100305
rect 273995 100215 274085 100305
rect 274175 100215 274265 100305
rect 274355 100215 274450 100305
rect 265350 100125 274450 100215
rect 265350 100035 265445 100125
rect 265535 100035 265625 100125
rect 265715 100035 265805 100125
rect 265895 100035 265985 100125
rect 266075 100035 266165 100125
rect 266255 100035 266345 100125
rect 266435 100035 266525 100125
rect 266615 100035 266705 100125
rect 266795 100035 266885 100125
rect 266975 100035 267065 100125
rect 267155 100035 267245 100125
rect 267335 100035 267425 100125
rect 267515 100035 267605 100125
rect 267695 100035 267785 100125
rect 267875 100035 267965 100125
rect 268055 100035 268145 100125
rect 268235 100035 268325 100125
rect 268415 100035 268505 100125
rect 268595 100035 268685 100125
rect 268775 100035 268865 100125
rect 268955 100035 269045 100125
rect 269135 100035 269225 100125
rect 269315 100035 269405 100125
rect 269495 100035 269585 100125
rect 269675 100035 269765 100125
rect 269855 100035 269945 100125
rect 270035 100035 270125 100125
rect 270215 100035 270305 100125
rect 270395 100035 270485 100125
rect 270575 100035 270665 100125
rect 270755 100035 270845 100125
rect 270935 100035 271025 100125
rect 271115 100035 271205 100125
rect 271295 100035 271385 100125
rect 271475 100035 271565 100125
rect 271655 100035 271745 100125
rect 271835 100035 271925 100125
rect 272015 100035 272105 100125
rect 272195 100035 272285 100125
rect 272375 100035 272465 100125
rect 272555 100035 272645 100125
rect 272735 100035 272825 100125
rect 272915 100035 273005 100125
rect 273095 100035 273185 100125
rect 273275 100035 273365 100125
rect 273455 100035 273545 100125
rect 273635 100035 273725 100125
rect 273815 100035 273905 100125
rect 273995 100035 274085 100125
rect 274175 100035 274265 100125
rect 274355 100035 274450 100125
rect 265350 99945 274450 100035
rect 265350 99855 265445 99945
rect 265535 99855 265625 99945
rect 265715 99855 265805 99945
rect 265895 99855 265985 99945
rect 266075 99855 266165 99945
rect 266255 99855 266345 99945
rect 266435 99855 266525 99945
rect 266615 99855 266705 99945
rect 266795 99855 266885 99945
rect 266975 99855 267065 99945
rect 267155 99855 267245 99945
rect 267335 99855 267425 99945
rect 267515 99855 267605 99945
rect 267695 99855 267785 99945
rect 267875 99855 267965 99945
rect 268055 99855 268145 99945
rect 268235 99855 268325 99945
rect 268415 99855 268505 99945
rect 268595 99855 268685 99945
rect 268775 99855 268865 99945
rect 268955 99855 269045 99945
rect 269135 99855 269225 99945
rect 269315 99855 269405 99945
rect 269495 99855 269585 99945
rect 269675 99855 269765 99945
rect 269855 99855 269945 99945
rect 270035 99855 270125 99945
rect 270215 99855 270305 99945
rect 270395 99855 270485 99945
rect 270575 99855 270665 99945
rect 270755 99855 270845 99945
rect 270935 99855 271025 99945
rect 271115 99855 271205 99945
rect 271295 99855 271385 99945
rect 271475 99855 271565 99945
rect 271655 99855 271745 99945
rect 271835 99855 271925 99945
rect 272015 99855 272105 99945
rect 272195 99855 272285 99945
rect 272375 99855 272465 99945
rect 272555 99855 272645 99945
rect 272735 99855 272825 99945
rect 272915 99855 273005 99945
rect 273095 99855 273185 99945
rect 273275 99855 273365 99945
rect 273455 99855 273545 99945
rect 273635 99855 273725 99945
rect 273815 99855 273905 99945
rect 273995 99855 274085 99945
rect 274175 99855 274265 99945
rect 274355 99855 274450 99945
rect 265350 99765 274450 99855
rect 265350 99675 265445 99765
rect 265535 99675 265625 99765
rect 265715 99675 265805 99765
rect 265895 99675 265985 99765
rect 266075 99675 266165 99765
rect 266255 99675 266345 99765
rect 266435 99675 266525 99765
rect 266615 99675 266705 99765
rect 266795 99675 266885 99765
rect 266975 99675 267065 99765
rect 267155 99675 267245 99765
rect 267335 99675 267425 99765
rect 267515 99675 267605 99765
rect 267695 99675 267785 99765
rect 267875 99675 267965 99765
rect 268055 99675 268145 99765
rect 268235 99675 268325 99765
rect 268415 99675 268505 99765
rect 268595 99675 268685 99765
rect 268775 99675 268865 99765
rect 268955 99675 269045 99765
rect 269135 99675 269225 99765
rect 269315 99675 269405 99765
rect 269495 99675 269585 99765
rect 269675 99675 269765 99765
rect 269855 99675 269945 99765
rect 270035 99675 270125 99765
rect 270215 99675 270305 99765
rect 270395 99675 270485 99765
rect 270575 99675 270665 99765
rect 270755 99675 270845 99765
rect 270935 99675 271025 99765
rect 271115 99675 271205 99765
rect 271295 99675 271385 99765
rect 271475 99675 271565 99765
rect 271655 99675 271745 99765
rect 271835 99675 271925 99765
rect 272015 99675 272105 99765
rect 272195 99675 272285 99765
rect 272375 99675 272465 99765
rect 272555 99675 272645 99765
rect 272735 99675 272825 99765
rect 272915 99675 273005 99765
rect 273095 99675 273185 99765
rect 273275 99675 273365 99765
rect 273455 99675 273545 99765
rect 273635 99675 273725 99765
rect 273815 99675 273905 99765
rect 273995 99675 274085 99765
rect 274175 99675 274265 99765
rect 274355 99675 274450 99765
rect 265350 99585 274450 99675
rect 265350 99495 265445 99585
rect 265535 99495 265625 99585
rect 265715 99495 265805 99585
rect 265895 99495 265985 99585
rect 266075 99495 266165 99585
rect 266255 99495 266345 99585
rect 266435 99495 266525 99585
rect 266615 99495 266705 99585
rect 266795 99495 266885 99585
rect 266975 99495 267065 99585
rect 267155 99495 267245 99585
rect 267335 99495 267425 99585
rect 267515 99495 267605 99585
rect 267695 99495 267785 99585
rect 267875 99495 267965 99585
rect 268055 99495 268145 99585
rect 268235 99495 268325 99585
rect 268415 99495 268505 99585
rect 268595 99495 268685 99585
rect 268775 99495 268865 99585
rect 268955 99495 269045 99585
rect 269135 99495 269225 99585
rect 269315 99495 269405 99585
rect 269495 99495 269585 99585
rect 269675 99495 269765 99585
rect 269855 99495 269945 99585
rect 270035 99495 270125 99585
rect 270215 99495 270305 99585
rect 270395 99495 270485 99585
rect 270575 99495 270665 99585
rect 270755 99495 270845 99585
rect 270935 99495 271025 99585
rect 271115 99495 271205 99585
rect 271295 99495 271385 99585
rect 271475 99495 271565 99585
rect 271655 99495 271745 99585
rect 271835 99495 271925 99585
rect 272015 99495 272105 99585
rect 272195 99495 272285 99585
rect 272375 99495 272465 99585
rect 272555 99495 272645 99585
rect 272735 99495 272825 99585
rect 272915 99495 273005 99585
rect 273095 99495 273185 99585
rect 273275 99495 273365 99585
rect 273455 99495 273545 99585
rect 273635 99495 273725 99585
rect 273815 99495 273905 99585
rect 273995 99495 274085 99585
rect 274175 99495 274265 99585
rect 274355 99495 274450 99585
rect 265350 99350 274450 99495
<< m2contact >>
rect 106655 280325 106745 280415
rect 106835 280325 106925 280415
rect 107015 280325 107105 280415
rect 107195 280325 107285 280415
rect 107375 280325 107465 280415
rect 107555 280325 107645 280415
rect 107735 280325 107825 280415
rect 107915 280325 108005 280415
rect 108095 280325 108185 280415
rect 108275 280325 108365 280415
rect 108455 280325 108545 280415
rect 108635 280325 108725 280415
rect 108815 280325 108905 280415
rect 108995 280325 109085 280415
rect 109175 280325 109265 280415
rect 109355 280325 109445 280415
rect 109535 280325 109625 280415
rect 109715 280325 109805 280415
rect 109895 280325 109985 280415
rect 110075 280325 110165 280415
rect 110255 280325 110345 280415
rect 110435 280325 110525 280415
rect 110615 280325 110705 280415
rect 110795 280325 110885 280415
rect 110975 280325 111065 280415
rect 111155 280325 111245 280415
rect 111335 280325 111425 280415
rect 111515 280325 111605 280415
rect 111695 280325 111785 280415
rect 111875 280325 111965 280415
rect 112055 280325 112145 280415
rect 112235 280325 112325 280415
rect 112415 280325 112505 280415
rect 112595 280325 112685 280415
rect 112775 280325 112865 280415
rect 112955 280325 113045 280415
rect 106655 280145 106745 280235
rect 106835 280145 106925 280235
rect 107015 280145 107105 280235
rect 107195 280145 107285 280235
rect 107375 280145 107465 280235
rect 107555 280145 107645 280235
rect 107735 280145 107825 280235
rect 107915 280145 108005 280235
rect 108095 280145 108185 280235
rect 108275 280145 108365 280235
rect 108455 280145 108545 280235
rect 108635 280145 108725 280235
rect 108815 280145 108905 280235
rect 108995 280145 109085 280235
rect 109175 280145 109265 280235
rect 109355 280145 109445 280235
rect 109535 280145 109625 280235
rect 109715 280145 109805 280235
rect 109895 280145 109985 280235
rect 110075 280145 110165 280235
rect 110255 280145 110345 280235
rect 110435 280145 110525 280235
rect 110615 280145 110705 280235
rect 110795 280145 110885 280235
rect 110975 280145 111065 280235
rect 111155 280145 111245 280235
rect 111335 280145 111425 280235
rect 111515 280145 111605 280235
rect 111695 280145 111785 280235
rect 111875 280145 111965 280235
rect 112055 280145 112145 280235
rect 112235 280145 112325 280235
rect 112415 280145 112505 280235
rect 112595 280145 112685 280235
rect 112775 280145 112865 280235
rect 112955 280145 113045 280235
rect 106655 279965 106745 280055
rect 106835 279965 106925 280055
rect 107015 279965 107105 280055
rect 107195 279965 107285 280055
rect 107375 279965 107465 280055
rect 107555 279965 107645 280055
rect 107735 279965 107825 280055
rect 107915 279965 108005 280055
rect 108095 279965 108185 280055
rect 108275 279965 108365 280055
rect 108455 279965 108545 280055
rect 108635 279965 108725 280055
rect 108815 279965 108905 280055
rect 108995 279965 109085 280055
rect 109175 279965 109265 280055
rect 109355 279965 109445 280055
rect 109535 279965 109625 280055
rect 109715 279965 109805 280055
rect 109895 279965 109985 280055
rect 110075 279965 110165 280055
rect 110255 279965 110345 280055
rect 110435 279965 110525 280055
rect 110615 279965 110705 280055
rect 110795 279965 110885 280055
rect 110975 279965 111065 280055
rect 111155 279965 111245 280055
rect 111335 279965 111425 280055
rect 111515 279965 111605 280055
rect 111695 279965 111785 280055
rect 111875 279965 111965 280055
rect 112055 279965 112145 280055
rect 112235 279965 112325 280055
rect 112415 279965 112505 280055
rect 112595 279965 112685 280055
rect 112775 279965 112865 280055
rect 112955 279965 113045 280055
rect 106655 279785 106745 279875
rect 106835 279785 106925 279875
rect 107015 279785 107105 279875
rect 107195 279785 107285 279875
rect 107375 279785 107465 279875
rect 107555 279785 107645 279875
rect 107735 279785 107825 279875
rect 107915 279785 108005 279875
rect 108095 279785 108185 279875
rect 108275 279785 108365 279875
rect 108455 279785 108545 279875
rect 108635 279785 108725 279875
rect 108815 279785 108905 279875
rect 108995 279785 109085 279875
rect 109175 279785 109265 279875
rect 109355 279785 109445 279875
rect 109535 279785 109625 279875
rect 109715 279785 109805 279875
rect 109895 279785 109985 279875
rect 110075 279785 110165 279875
rect 110255 279785 110345 279875
rect 110435 279785 110525 279875
rect 110615 279785 110705 279875
rect 110795 279785 110885 279875
rect 110975 279785 111065 279875
rect 111155 279785 111245 279875
rect 111335 279785 111425 279875
rect 111515 279785 111605 279875
rect 111695 279785 111785 279875
rect 111875 279785 111965 279875
rect 112055 279785 112145 279875
rect 112235 279785 112325 279875
rect 112415 279785 112505 279875
rect 112595 279785 112685 279875
rect 112775 279785 112865 279875
rect 112955 279785 113045 279875
rect 265445 280355 265535 280445
rect 265625 280355 265715 280445
rect 265805 280355 265895 280445
rect 265985 280355 266075 280445
rect 266165 280355 266255 280445
rect 266345 280355 266435 280445
rect 266525 280355 266615 280445
rect 266705 280355 266795 280445
rect 266885 280355 266975 280445
rect 267065 280355 267155 280445
rect 267245 280355 267335 280445
rect 267425 280355 267515 280445
rect 267605 280355 267695 280445
rect 267785 280355 267875 280445
rect 267965 280355 268055 280445
rect 268145 280355 268235 280445
rect 268325 280355 268415 280445
rect 268505 280355 268595 280445
rect 268685 280355 268775 280445
rect 268865 280355 268955 280445
rect 269045 280355 269135 280445
rect 269225 280355 269315 280445
rect 269405 280355 269495 280445
rect 269585 280355 269675 280445
rect 269765 280355 269855 280445
rect 269945 280355 270035 280445
rect 270125 280355 270215 280445
rect 270305 280355 270395 280445
rect 270485 280355 270575 280445
rect 270665 280355 270755 280445
rect 270845 280355 270935 280445
rect 271025 280355 271115 280445
rect 271205 280355 271295 280445
rect 271385 280355 271475 280445
rect 271565 280355 271655 280445
rect 271745 280355 271835 280445
rect 271925 280355 272015 280445
rect 272105 280355 272195 280445
rect 272285 280355 272375 280445
rect 272465 280355 272555 280445
rect 272645 280355 272735 280445
rect 272825 280355 272915 280445
rect 273005 280355 273095 280445
rect 273185 280355 273275 280445
rect 273365 280355 273455 280445
rect 273545 280355 273635 280445
rect 273725 280355 273815 280445
rect 273905 280355 273995 280445
rect 274085 280355 274175 280445
rect 274265 280355 274355 280445
rect 265445 280175 265535 280265
rect 265625 280175 265715 280265
rect 265805 280175 265895 280265
rect 265985 280175 266075 280265
rect 266165 280175 266255 280265
rect 266345 280175 266435 280265
rect 266525 280175 266615 280265
rect 266705 280175 266795 280265
rect 266885 280175 266975 280265
rect 267065 280175 267155 280265
rect 267245 280175 267335 280265
rect 267425 280175 267515 280265
rect 267605 280175 267695 280265
rect 267785 280175 267875 280265
rect 267965 280175 268055 280265
rect 268145 280175 268235 280265
rect 268325 280175 268415 280265
rect 268505 280175 268595 280265
rect 268685 280175 268775 280265
rect 268865 280175 268955 280265
rect 269045 280175 269135 280265
rect 269225 280175 269315 280265
rect 269405 280175 269495 280265
rect 269585 280175 269675 280265
rect 269765 280175 269855 280265
rect 269945 280175 270035 280265
rect 270125 280175 270215 280265
rect 270305 280175 270395 280265
rect 270485 280175 270575 280265
rect 270665 280175 270755 280265
rect 270845 280175 270935 280265
rect 271025 280175 271115 280265
rect 271205 280175 271295 280265
rect 271385 280175 271475 280265
rect 271565 280175 271655 280265
rect 271745 280175 271835 280265
rect 271925 280175 272015 280265
rect 272105 280175 272195 280265
rect 272285 280175 272375 280265
rect 272465 280175 272555 280265
rect 272645 280175 272735 280265
rect 272825 280175 272915 280265
rect 273005 280175 273095 280265
rect 273185 280175 273275 280265
rect 273365 280175 273455 280265
rect 273545 280175 273635 280265
rect 273725 280175 273815 280265
rect 273905 280175 273995 280265
rect 274085 280175 274175 280265
rect 274265 280175 274355 280265
rect 265445 279995 265535 280085
rect 265625 279995 265715 280085
rect 265805 279995 265895 280085
rect 265985 279995 266075 280085
rect 266165 279995 266255 280085
rect 266345 279995 266435 280085
rect 266525 279995 266615 280085
rect 266705 279995 266795 280085
rect 266885 279995 266975 280085
rect 267065 279995 267155 280085
rect 267245 279995 267335 280085
rect 267425 279995 267515 280085
rect 267605 279995 267695 280085
rect 267785 279995 267875 280085
rect 267965 279995 268055 280085
rect 268145 279995 268235 280085
rect 268325 279995 268415 280085
rect 268505 279995 268595 280085
rect 268685 279995 268775 280085
rect 268865 279995 268955 280085
rect 269045 279995 269135 280085
rect 269225 279995 269315 280085
rect 269405 279995 269495 280085
rect 269585 279995 269675 280085
rect 269765 279995 269855 280085
rect 269945 279995 270035 280085
rect 270125 279995 270215 280085
rect 270305 279995 270395 280085
rect 270485 279995 270575 280085
rect 270665 279995 270755 280085
rect 270845 279995 270935 280085
rect 271025 279995 271115 280085
rect 271205 279995 271295 280085
rect 271385 279995 271475 280085
rect 271565 279995 271655 280085
rect 271745 279995 271835 280085
rect 271925 279995 272015 280085
rect 272105 279995 272195 280085
rect 272285 279995 272375 280085
rect 272465 279995 272555 280085
rect 272645 279995 272735 280085
rect 272825 279995 272915 280085
rect 273005 279995 273095 280085
rect 273185 279995 273275 280085
rect 273365 279995 273455 280085
rect 273545 279995 273635 280085
rect 273725 279995 273815 280085
rect 273905 279995 273995 280085
rect 274085 279995 274175 280085
rect 274265 279995 274355 280085
rect 265445 279815 265535 279905
rect 265625 279815 265715 279905
rect 265805 279815 265895 279905
rect 265985 279815 266075 279905
rect 266165 279815 266255 279905
rect 266345 279815 266435 279905
rect 266525 279815 266615 279905
rect 266705 279815 266795 279905
rect 266885 279815 266975 279905
rect 267065 279815 267155 279905
rect 267245 279815 267335 279905
rect 267425 279815 267515 279905
rect 267605 279815 267695 279905
rect 267785 279815 267875 279905
rect 267965 279815 268055 279905
rect 268145 279815 268235 279905
rect 268325 279815 268415 279905
rect 268505 279815 268595 279905
rect 268685 279815 268775 279905
rect 268865 279815 268955 279905
rect 269045 279815 269135 279905
rect 269225 279815 269315 279905
rect 269405 279815 269495 279905
rect 269585 279815 269675 279905
rect 269765 279815 269855 279905
rect 269945 279815 270035 279905
rect 270125 279815 270215 279905
rect 270305 279815 270395 279905
rect 270485 279815 270575 279905
rect 270665 279815 270755 279905
rect 270845 279815 270935 279905
rect 271025 279815 271115 279905
rect 271205 279815 271295 279905
rect 271385 279815 271475 279905
rect 271565 279815 271655 279905
rect 271745 279815 271835 279905
rect 271925 279815 272015 279905
rect 272105 279815 272195 279905
rect 272285 279815 272375 279905
rect 272465 279815 272555 279905
rect 272645 279815 272735 279905
rect 272825 279815 272915 279905
rect 273005 279815 273095 279905
rect 273185 279815 273275 279905
rect 273365 279815 273455 279905
rect 273545 279815 273635 279905
rect 273725 279815 273815 279905
rect 273905 279815 273995 279905
rect 274085 279815 274175 279905
rect 274265 279815 274355 279905
rect 265445 279635 265535 279725
rect 265625 279635 265715 279725
rect 265805 279635 265895 279725
rect 265985 279635 266075 279725
rect 266165 279635 266255 279725
rect 266345 279635 266435 279725
rect 266525 279635 266615 279725
rect 266705 279635 266795 279725
rect 266885 279635 266975 279725
rect 267065 279635 267155 279725
rect 267245 279635 267335 279725
rect 267425 279635 267515 279725
rect 267605 279635 267695 279725
rect 267785 279635 267875 279725
rect 267965 279635 268055 279725
rect 268145 279635 268235 279725
rect 268325 279635 268415 279725
rect 268505 279635 268595 279725
rect 268685 279635 268775 279725
rect 268865 279635 268955 279725
rect 269045 279635 269135 279725
rect 269225 279635 269315 279725
rect 269405 279635 269495 279725
rect 269585 279635 269675 279725
rect 269765 279635 269855 279725
rect 269945 279635 270035 279725
rect 270125 279635 270215 279725
rect 270305 279635 270395 279725
rect 270485 279635 270575 279725
rect 270665 279635 270755 279725
rect 270845 279635 270935 279725
rect 271025 279635 271115 279725
rect 271205 279635 271295 279725
rect 271385 279635 271475 279725
rect 271565 279635 271655 279725
rect 271745 279635 271835 279725
rect 271925 279635 272015 279725
rect 272105 279635 272195 279725
rect 272285 279635 272375 279725
rect 272465 279635 272555 279725
rect 272645 279635 272735 279725
rect 272825 279635 272915 279725
rect 273005 279635 273095 279725
rect 273185 279635 273275 279725
rect 273365 279635 273455 279725
rect 273545 279635 273635 279725
rect 273725 279635 273815 279725
rect 273905 279635 273995 279725
rect 274085 279635 274175 279725
rect 274265 279635 274355 279725
rect 265445 279455 265535 279545
rect 265625 279455 265715 279545
rect 265805 279455 265895 279545
rect 265985 279455 266075 279545
rect 266165 279455 266255 279545
rect 266345 279455 266435 279545
rect 266525 279455 266615 279545
rect 266705 279455 266795 279545
rect 266885 279455 266975 279545
rect 267065 279455 267155 279545
rect 267245 279455 267335 279545
rect 267425 279455 267515 279545
rect 267605 279455 267695 279545
rect 267785 279455 267875 279545
rect 267965 279455 268055 279545
rect 268145 279455 268235 279545
rect 268325 279455 268415 279545
rect 268505 279455 268595 279545
rect 268685 279455 268775 279545
rect 268865 279455 268955 279545
rect 269045 279455 269135 279545
rect 269225 279455 269315 279545
rect 269405 279455 269495 279545
rect 269585 279455 269675 279545
rect 269765 279455 269855 279545
rect 269945 279455 270035 279545
rect 270125 279455 270215 279545
rect 270305 279455 270395 279545
rect 270485 279455 270575 279545
rect 270665 279455 270755 279545
rect 270845 279455 270935 279545
rect 271025 279455 271115 279545
rect 271205 279455 271295 279545
rect 271385 279455 271475 279545
rect 271565 279455 271655 279545
rect 271745 279455 271835 279545
rect 271925 279455 272015 279545
rect 272105 279455 272195 279545
rect 272285 279455 272375 279545
rect 272465 279455 272555 279545
rect 272645 279455 272735 279545
rect 272825 279455 272915 279545
rect 273005 279455 273095 279545
rect 273185 279455 273275 279545
rect 273365 279455 273455 279545
rect 273545 279455 273635 279545
rect 273725 279455 273815 279545
rect 273905 279455 273995 279545
rect 274085 279455 274175 279545
rect 274265 279455 274355 279545
rect 106655 100265 106745 100355
rect 106835 100265 106925 100355
rect 107015 100265 107105 100355
rect 107195 100265 107285 100355
rect 107375 100265 107465 100355
rect 107555 100265 107645 100355
rect 107735 100265 107825 100355
rect 107915 100265 108005 100355
rect 108095 100265 108185 100355
rect 108275 100265 108365 100355
rect 108455 100265 108545 100355
rect 108635 100265 108725 100355
rect 108815 100265 108905 100355
rect 108995 100265 109085 100355
rect 109175 100265 109265 100355
rect 109355 100265 109445 100355
rect 109535 100265 109625 100355
rect 109715 100265 109805 100355
rect 109895 100265 109985 100355
rect 110075 100265 110165 100355
rect 110255 100265 110345 100355
rect 110435 100265 110525 100355
rect 110615 100265 110705 100355
rect 110795 100265 110885 100355
rect 110975 100265 111065 100355
rect 111155 100265 111245 100355
rect 111335 100265 111425 100355
rect 111515 100265 111605 100355
rect 111695 100265 111785 100355
rect 111875 100265 111965 100355
rect 112055 100265 112145 100355
rect 112235 100265 112325 100355
rect 112415 100265 112505 100355
rect 112595 100265 112685 100355
rect 112775 100265 112865 100355
rect 112955 100265 113045 100355
rect 106655 100085 106745 100175
rect 106835 100085 106925 100175
rect 107015 100085 107105 100175
rect 107195 100085 107285 100175
rect 107375 100085 107465 100175
rect 107555 100085 107645 100175
rect 107735 100085 107825 100175
rect 107915 100085 108005 100175
rect 108095 100085 108185 100175
rect 108275 100085 108365 100175
rect 108455 100085 108545 100175
rect 108635 100085 108725 100175
rect 108815 100085 108905 100175
rect 108995 100085 109085 100175
rect 109175 100085 109265 100175
rect 109355 100085 109445 100175
rect 109535 100085 109625 100175
rect 109715 100085 109805 100175
rect 109895 100085 109985 100175
rect 110075 100085 110165 100175
rect 110255 100085 110345 100175
rect 110435 100085 110525 100175
rect 110615 100085 110705 100175
rect 110795 100085 110885 100175
rect 110975 100085 111065 100175
rect 111155 100085 111245 100175
rect 111335 100085 111425 100175
rect 111515 100085 111605 100175
rect 111695 100085 111785 100175
rect 111875 100085 111965 100175
rect 112055 100085 112145 100175
rect 112235 100085 112325 100175
rect 112415 100085 112505 100175
rect 112595 100085 112685 100175
rect 112775 100085 112865 100175
rect 112955 100085 113045 100175
rect 106655 99905 106745 99995
rect 106835 99905 106925 99995
rect 107015 99905 107105 99995
rect 107195 99905 107285 99995
rect 107375 99905 107465 99995
rect 107555 99905 107645 99995
rect 107735 99905 107825 99995
rect 107915 99905 108005 99995
rect 108095 99905 108185 99995
rect 108275 99905 108365 99995
rect 108455 99905 108545 99995
rect 108635 99905 108725 99995
rect 108815 99905 108905 99995
rect 108995 99905 109085 99995
rect 109175 99905 109265 99995
rect 109355 99905 109445 99995
rect 109535 99905 109625 99995
rect 109715 99905 109805 99995
rect 109895 99905 109985 99995
rect 110075 99905 110165 99995
rect 110255 99905 110345 99995
rect 110435 99905 110525 99995
rect 110615 99905 110705 99995
rect 110795 99905 110885 99995
rect 110975 99905 111065 99995
rect 111155 99905 111245 99995
rect 111335 99905 111425 99995
rect 111515 99905 111605 99995
rect 111695 99905 111785 99995
rect 111875 99905 111965 99995
rect 112055 99905 112145 99995
rect 112235 99905 112325 99995
rect 112415 99905 112505 99995
rect 112595 99905 112685 99995
rect 112775 99905 112865 99995
rect 112955 99905 113045 99995
rect 106655 99725 106745 99815
rect 106835 99725 106925 99815
rect 107015 99725 107105 99815
rect 107195 99725 107285 99815
rect 107375 99725 107465 99815
rect 107555 99725 107645 99815
rect 107735 99725 107825 99815
rect 107915 99725 108005 99815
rect 108095 99725 108185 99815
rect 108275 99725 108365 99815
rect 108455 99725 108545 99815
rect 108635 99725 108725 99815
rect 108815 99725 108905 99815
rect 108995 99725 109085 99815
rect 109175 99725 109265 99815
rect 109355 99725 109445 99815
rect 109535 99725 109625 99815
rect 109715 99725 109805 99815
rect 109895 99725 109985 99815
rect 110075 99725 110165 99815
rect 110255 99725 110345 99815
rect 110435 99725 110525 99815
rect 110615 99725 110705 99815
rect 110795 99725 110885 99815
rect 110975 99725 111065 99815
rect 111155 99725 111245 99815
rect 111335 99725 111425 99815
rect 111515 99725 111605 99815
rect 111695 99725 111785 99815
rect 111875 99725 111965 99815
rect 112055 99725 112145 99815
rect 112235 99725 112325 99815
rect 112415 99725 112505 99815
rect 112595 99725 112685 99815
rect 112775 99725 112865 99815
rect 112955 99725 113045 99815
rect 106655 99545 106745 99635
rect 106835 99545 106925 99635
rect 107015 99545 107105 99635
rect 107195 99545 107285 99635
rect 107375 99545 107465 99635
rect 107555 99545 107645 99635
rect 107735 99545 107825 99635
rect 107915 99545 108005 99635
rect 108095 99545 108185 99635
rect 108275 99545 108365 99635
rect 108455 99545 108545 99635
rect 108635 99545 108725 99635
rect 108815 99545 108905 99635
rect 108995 99545 109085 99635
rect 109175 99545 109265 99635
rect 109355 99545 109445 99635
rect 109535 99545 109625 99635
rect 109715 99545 109805 99635
rect 109895 99545 109985 99635
rect 110075 99545 110165 99635
rect 110255 99545 110345 99635
rect 110435 99545 110525 99635
rect 110615 99545 110705 99635
rect 110795 99545 110885 99635
rect 110975 99545 111065 99635
rect 111155 99545 111245 99635
rect 111335 99545 111425 99635
rect 111515 99545 111605 99635
rect 111695 99545 111785 99635
rect 111875 99545 111965 99635
rect 112055 99545 112145 99635
rect 112235 99545 112325 99635
rect 112415 99545 112505 99635
rect 112595 99545 112685 99635
rect 112775 99545 112865 99635
rect 112955 99545 113045 99635
rect 265445 100215 265535 100305
rect 265625 100215 265715 100305
rect 265805 100215 265895 100305
rect 265985 100215 266075 100305
rect 266165 100215 266255 100305
rect 266345 100215 266435 100305
rect 266525 100215 266615 100305
rect 266705 100215 266795 100305
rect 266885 100215 266975 100305
rect 267065 100215 267155 100305
rect 267245 100215 267335 100305
rect 267425 100215 267515 100305
rect 267605 100215 267695 100305
rect 267785 100215 267875 100305
rect 267965 100215 268055 100305
rect 268145 100215 268235 100305
rect 268325 100215 268415 100305
rect 268505 100215 268595 100305
rect 268685 100215 268775 100305
rect 268865 100215 268955 100305
rect 269045 100215 269135 100305
rect 269225 100215 269315 100305
rect 269405 100215 269495 100305
rect 269585 100215 269675 100305
rect 269765 100215 269855 100305
rect 269945 100215 270035 100305
rect 270125 100215 270215 100305
rect 270305 100215 270395 100305
rect 270485 100215 270575 100305
rect 270665 100215 270755 100305
rect 270845 100215 270935 100305
rect 271025 100215 271115 100305
rect 271205 100215 271295 100305
rect 271385 100215 271475 100305
rect 271565 100215 271655 100305
rect 271745 100215 271835 100305
rect 271925 100215 272015 100305
rect 272105 100215 272195 100305
rect 272285 100215 272375 100305
rect 272465 100215 272555 100305
rect 272645 100215 272735 100305
rect 272825 100215 272915 100305
rect 273005 100215 273095 100305
rect 273185 100215 273275 100305
rect 273365 100215 273455 100305
rect 273545 100215 273635 100305
rect 273725 100215 273815 100305
rect 273905 100215 273995 100305
rect 274085 100215 274175 100305
rect 274265 100215 274355 100305
rect 265445 100035 265535 100125
rect 265625 100035 265715 100125
rect 265805 100035 265895 100125
rect 265985 100035 266075 100125
rect 266165 100035 266255 100125
rect 266345 100035 266435 100125
rect 266525 100035 266615 100125
rect 266705 100035 266795 100125
rect 266885 100035 266975 100125
rect 267065 100035 267155 100125
rect 267245 100035 267335 100125
rect 267425 100035 267515 100125
rect 267605 100035 267695 100125
rect 267785 100035 267875 100125
rect 267965 100035 268055 100125
rect 268145 100035 268235 100125
rect 268325 100035 268415 100125
rect 268505 100035 268595 100125
rect 268685 100035 268775 100125
rect 268865 100035 268955 100125
rect 269045 100035 269135 100125
rect 269225 100035 269315 100125
rect 269405 100035 269495 100125
rect 269585 100035 269675 100125
rect 269765 100035 269855 100125
rect 269945 100035 270035 100125
rect 270125 100035 270215 100125
rect 270305 100035 270395 100125
rect 270485 100035 270575 100125
rect 270665 100035 270755 100125
rect 270845 100035 270935 100125
rect 271025 100035 271115 100125
rect 271205 100035 271295 100125
rect 271385 100035 271475 100125
rect 271565 100035 271655 100125
rect 271745 100035 271835 100125
rect 271925 100035 272015 100125
rect 272105 100035 272195 100125
rect 272285 100035 272375 100125
rect 272465 100035 272555 100125
rect 272645 100035 272735 100125
rect 272825 100035 272915 100125
rect 273005 100035 273095 100125
rect 273185 100035 273275 100125
rect 273365 100035 273455 100125
rect 273545 100035 273635 100125
rect 273725 100035 273815 100125
rect 273905 100035 273995 100125
rect 274085 100035 274175 100125
rect 274265 100035 274355 100125
rect 265445 99855 265535 99945
rect 265625 99855 265715 99945
rect 265805 99855 265895 99945
rect 265985 99855 266075 99945
rect 266165 99855 266255 99945
rect 266345 99855 266435 99945
rect 266525 99855 266615 99945
rect 266705 99855 266795 99945
rect 266885 99855 266975 99945
rect 267065 99855 267155 99945
rect 267245 99855 267335 99945
rect 267425 99855 267515 99945
rect 267605 99855 267695 99945
rect 267785 99855 267875 99945
rect 267965 99855 268055 99945
rect 268145 99855 268235 99945
rect 268325 99855 268415 99945
rect 268505 99855 268595 99945
rect 268685 99855 268775 99945
rect 268865 99855 268955 99945
rect 269045 99855 269135 99945
rect 269225 99855 269315 99945
rect 269405 99855 269495 99945
rect 269585 99855 269675 99945
rect 269765 99855 269855 99945
rect 269945 99855 270035 99945
rect 270125 99855 270215 99945
rect 270305 99855 270395 99945
rect 270485 99855 270575 99945
rect 270665 99855 270755 99945
rect 270845 99855 270935 99945
rect 271025 99855 271115 99945
rect 271205 99855 271295 99945
rect 271385 99855 271475 99945
rect 271565 99855 271655 99945
rect 271745 99855 271835 99945
rect 271925 99855 272015 99945
rect 272105 99855 272195 99945
rect 272285 99855 272375 99945
rect 272465 99855 272555 99945
rect 272645 99855 272735 99945
rect 272825 99855 272915 99945
rect 273005 99855 273095 99945
rect 273185 99855 273275 99945
rect 273365 99855 273455 99945
rect 273545 99855 273635 99945
rect 273725 99855 273815 99945
rect 273905 99855 273995 99945
rect 274085 99855 274175 99945
rect 274265 99855 274355 99945
rect 265445 99675 265535 99765
rect 265625 99675 265715 99765
rect 265805 99675 265895 99765
rect 265985 99675 266075 99765
rect 266165 99675 266255 99765
rect 266345 99675 266435 99765
rect 266525 99675 266615 99765
rect 266705 99675 266795 99765
rect 266885 99675 266975 99765
rect 267065 99675 267155 99765
rect 267245 99675 267335 99765
rect 267425 99675 267515 99765
rect 267605 99675 267695 99765
rect 267785 99675 267875 99765
rect 267965 99675 268055 99765
rect 268145 99675 268235 99765
rect 268325 99675 268415 99765
rect 268505 99675 268595 99765
rect 268685 99675 268775 99765
rect 268865 99675 268955 99765
rect 269045 99675 269135 99765
rect 269225 99675 269315 99765
rect 269405 99675 269495 99765
rect 269585 99675 269675 99765
rect 269765 99675 269855 99765
rect 269945 99675 270035 99765
rect 270125 99675 270215 99765
rect 270305 99675 270395 99765
rect 270485 99675 270575 99765
rect 270665 99675 270755 99765
rect 270845 99675 270935 99765
rect 271025 99675 271115 99765
rect 271205 99675 271295 99765
rect 271385 99675 271475 99765
rect 271565 99675 271655 99765
rect 271745 99675 271835 99765
rect 271925 99675 272015 99765
rect 272105 99675 272195 99765
rect 272285 99675 272375 99765
rect 272465 99675 272555 99765
rect 272645 99675 272735 99765
rect 272825 99675 272915 99765
rect 273005 99675 273095 99765
rect 273185 99675 273275 99765
rect 273365 99675 273455 99765
rect 273545 99675 273635 99765
rect 273725 99675 273815 99765
rect 273905 99675 273995 99765
rect 274085 99675 274175 99765
rect 274265 99675 274355 99765
rect 265445 99495 265535 99585
rect 265625 99495 265715 99585
rect 265805 99495 265895 99585
rect 265985 99495 266075 99585
rect 266165 99495 266255 99585
rect 266345 99495 266435 99585
rect 266525 99495 266615 99585
rect 266705 99495 266795 99585
rect 266885 99495 266975 99585
rect 267065 99495 267155 99585
rect 267245 99495 267335 99585
rect 267425 99495 267515 99585
rect 267605 99495 267695 99585
rect 267785 99495 267875 99585
rect 267965 99495 268055 99585
rect 268145 99495 268235 99585
rect 268325 99495 268415 99585
rect 268505 99495 268595 99585
rect 268685 99495 268775 99585
rect 268865 99495 268955 99585
rect 269045 99495 269135 99585
rect 269225 99495 269315 99585
rect 269405 99495 269495 99585
rect 269585 99495 269675 99585
rect 269765 99495 269855 99585
rect 269945 99495 270035 99585
rect 270125 99495 270215 99585
rect 270305 99495 270395 99585
rect 270485 99495 270575 99585
rect 270665 99495 270755 99585
rect 270845 99495 270935 99585
rect 271025 99495 271115 99585
rect 271205 99495 271295 99585
rect 271385 99495 271475 99585
rect 271565 99495 271655 99585
rect 271745 99495 271835 99585
rect 271925 99495 272015 99585
rect 272105 99495 272195 99585
rect 272285 99495 272375 99585
rect 272465 99495 272555 99585
rect 272645 99495 272735 99585
rect 272825 99495 272915 99585
rect 273005 99495 273095 99585
rect 273185 99495 273275 99585
rect 273365 99495 273455 99585
rect 273545 99495 273635 99585
rect 273725 99495 273815 99585
rect 273905 99495 273995 99585
rect 274085 99495 274175 99585
rect 274265 99495 274355 99585
<< metal2 >>
rect 106550 280415 113150 280550
rect 106550 280325 106655 280415
rect 106745 280325 106835 280415
rect 106925 280325 107015 280415
rect 107105 280325 107195 280415
rect 107285 280325 107375 280415
rect 107465 280325 107555 280415
rect 107645 280325 107735 280415
rect 107825 280325 107915 280415
rect 108005 280325 108095 280415
rect 108185 280325 108275 280415
rect 108365 280325 108455 280415
rect 108545 280325 108635 280415
rect 108725 280325 108815 280415
rect 108905 280325 108995 280415
rect 109085 280325 109175 280415
rect 109265 280325 109355 280415
rect 109445 280325 109535 280415
rect 109625 280325 109715 280415
rect 109805 280325 109895 280415
rect 109985 280325 110075 280415
rect 110165 280325 110255 280415
rect 110345 280325 110435 280415
rect 110525 280325 110615 280415
rect 110705 280325 110795 280415
rect 110885 280325 110975 280415
rect 111065 280325 111155 280415
rect 111245 280325 111335 280415
rect 111425 280325 111515 280415
rect 111605 280325 111695 280415
rect 111785 280325 111875 280415
rect 111965 280325 112055 280415
rect 112145 280325 112235 280415
rect 112325 280325 112415 280415
rect 112505 280325 112595 280415
rect 112685 280325 112775 280415
rect 112865 280325 112955 280415
rect 113045 280325 113150 280415
rect 106550 280235 113150 280325
rect 106550 280145 106655 280235
rect 106745 280145 106835 280235
rect 106925 280145 107015 280235
rect 107105 280145 107195 280235
rect 107285 280145 107375 280235
rect 107465 280145 107555 280235
rect 107645 280145 107735 280235
rect 107825 280145 107915 280235
rect 108005 280145 108095 280235
rect 108185 280145 108275 280235
rect 108365 280145 108455 280235
rect 108545 280145 108635 280235
rect 108725 280145 108815 280235
rect 108905 280145 108995 280235
rect 109085 280145 109175 280235
rect 109265 280145 109355 280235
rect 109445 280145 109535 280235
rect 109625 280145 109715 280235
rect 109805 280145 109895 280235
rect 109985 280145 110075 280235
rect 110165 280145 110255 280235
rect 110345 280145 110435 280235
rect 110525 280145 110615 280235
rect 110705 280145 110795 280235
rect 110885 280145 110975 280235
rect 111065 280145 111155 280235
rect 111245 280145 111335 280235
rect 111425 280145 111515 280235
rect 111605 280145 111695 280235
rect 111785 280145 111875 280235
rect 111965 280145 112055 280235
rect 112145 280145 112235 280235
rect 112325 280145 112415 280235
rect 112505 280145 112595 280235
rect 112685 280145 112775 280235
rect 112865 280145 112955 280235
rect 113045 280145 113150 280235
rect 106550 280055 113150 280145
rect 106550 279965 106655 280055
rect 106745 279965 106835 280055
rect 106925 279965 107015 280055
rect 107105 279965 107195 280055
rect 107285 279965 107375 280055
rect 107465 279965 107555 280055
rect 107645 279965 107735 280055
rect 107825 279965 107915 280055
rect 108005 279965 108095 280055
rect 108185 279965 108275 280055
rect 108365 279965 108455 280055
rect 108545 279965 108635 280055
rect 108725 279965 108815 280055
rect 108905 279965 108995 280055
rect 109085 279965 109175 280055
rect 109265 279965 109355 280055
rect 109445 279965 109535 280055
rect 109625 279965 109715 280055
rect 109805 279965 109895 280055
rect 109985 279965 110075 280055
rect 110165 279965 110255 280055
rect 110345 279965 110435 280055
rect 110525 279965 110615 280055
rect 110705 279965 110795 280055
rect 110885 279965 110975 280055
rect 111065 279965 111155 280055
rect 111245 279965 111335 280055
rect 111425 279965 111515 280055
rect 111605 279965 111695 280055
rect 111785 279965 111875 280055
rect 111965 279965 112055 280055
rect 112145 279965 112235 280055
rect 112325 279965 112415 280055
rect 112505 279965 112595 280055
rect 112685 279965 112775 280055
rect 112865 279965 112955 280055
rect 113045 279965 113150 280055
rect 106550 279875 113150 279965
rect 106550 279785 106655 279875
rect 106745 279785 106835 279875
rect 106925 279785 107015 279875
rect 107105 279785 107195 279875
rect 107285 279785 107375 279875
rect 107465 279785 107555 279875
rect 107645 279785 107735 279875
rect 107825 279785 107915 279875
rect 108005 279785 108095 279875
rect 108185 279785 108275 279875
rect 108365 279785 108455 279875
rect 108545 279785 108635 279875
rect 108725 279785 108815 279875
rect 108905 279785 108995 279875
rect 109085 279785 109175 279875
rect 109265 279785 109355 279875
rect 109445 279785 109535 279875
rect 109625 279785 109715 279875
rect 109805 279785 109895 279875
rect 109985 279785 110075 279875
rect 110165 279785 110255 279875
rect 110345 279785 110435 279875
rect 110525 279785 110615 279875
rect 110705 279785 110795 279875
rect 110885 279785 110975 279875
rect 111065 279785 111155 279875
rect 111245 279785 111335 279875
rect 111425 279785 111515 279875
rect 111605 279785 111695 279875
rect 111785 279785 111875 279875
rect 111965 279785 112055 279875
rect 112145 279785 112235 279875
rect 112325 279785 112415 279875
rect 112505 279785 112595 279875
rect 112685 279785 112775 279875
rect 112865 279785 112955 279875
rect 113045 279785 113150 279875
rect 106550 279650 113150 279785
rect 120450 274550 120800 280550
rect 136450 275150 136800 280550
rect 152450 275750 152800 280550
rect 168450 276350 168800 280550
rect 184450 278450 184800 280550
rect 181650 278150 184800 278450
rect 168450 276050 178350 276350
rect 152450 275450 177350 275750
rect 136450 274850 176250 275150
rect 120450 274250 170850 274550
rect 100950 273650 137200 273950
rect 100950 264700 101250 273650
rect 99400 264350 101250 264700
rect 101550 273050 135350 273350
rect 101550 259500 101850 273050
rect 99400 259150 101850 259500
rect 102150 272450 131600 272750
rect 102150 232700 102450 272450
rect 99400 232350 102450 232700
rect 102750 271850 126350 272150
rect 102750 216700 103050 271850
rect 99400 216350 103050 216700
rect 103350 271250 111050 271550
rect 126050 271250 126350 271850
rect 131250 271300 131600 272450
rect 135050 271250 135350 273050
rect 103350 200750 103650 271250
rect 110750 271150 111050 271250
rect 136900 271200 137200 273650
rect 170500 271250 170850 274250
rect 175850 271250 176250 274850
rect 176950 271250 177350 275450
rect 177950 271250 178350 276050
rect 181650 271250 181950 278150
rect 200450 277850 200800 280550
rect 182850 277550 200800 277850
rect 182850 271250 183150 277550
rect 216450 277250 216800 280500
rect 185450 276950 216800 277250
rect 185450 271250 185750 276950
rect 232450 276650 232800 280550
rect 187015 276350 232800 276650
rect 187015 271249 187296 276350
rect 248450 276050 248800 280550
rect 265350 280445 274450 280550
rect 265350 280355 265445 280445
rect 265535 280355 265625 280445
rect 265715 280355 265805 280445
rect 265895 280355 265985 280445
rect 266075 280355 266165 280445
rect 266255 280355 266345 280445
rect 266435 280355 266525 280445
rect 266615 280355 266705 280445
rect 266795 280355 266885 280445
rect 266975 280355 267065 280445
rect 267155 280355 267245 280445
rect 267335 280355 267425 280445
rect 267515 280355 267605 280445
rect 267695 280355 267785 280445
rect 267875 280355 267965 280445
rect 268055 280355 268145 280445
rect 268235 280355 268325 280445
rect 268415 280355 268505 280445
rect 268595 280355 268685 280445
rect 268775 280355 268865 280445
rect 268955 280355 269045 280445
rect 269135 280355 269225 280445
rect 269315 280355 269405 280445
rect 269495 280355 269585 280445
rect 269675 280355 269765 280445
rect 269855 280355 269945 280445
rect 270035 280355 270125 280445
rect 270215 280355 270305 280445
rect 270395 280355 270485 280445
rect 270575 280355 270665 280445
rect 270755 280355 270845 280445
rect 270935 280355 271025 280445
rect 271115 280355 271205 280445
rect 271295 280355 271385 280445
rect 271475 280355 271565 280445
rect 271655 280355 271745 280445
rect 271835 280355 271925 280445
rect 272015 280355 272105 280445
rect 272195 280355 272285 280445
rect 272375 280355 272465 280445
rect 272555 280355 272645 280445
rect 272735 280355 272825 280445
rect 272915 280355 273005 280445
rect 273095 280355 273185 280445
rect 273275 280355 273365 280445
rect 273455 280355 273545 280445
rect 273635 280355 273725 280445
rect 273815 280355 273905 280445
rect 273995 280355 274085 280445
rect 274175 280355 274265 280445
rect 274355 280355 274450 280445
rect 265350 280265 274450 280355
rect 265350 280175 265445 280265
rect 265535 280175 265625 280265
rect 265715 280175 265805 280265
rect 265895 280175 265985 280265
rect 266075 280175 266165 280265
rect 266255 280175 266345 280265
rect 266435 280175 266525 280265
rect 266615 280175 266705 280265
rect 266795 280175 266885 280265
rect 266975 280175 267065 280265
rect 267155 280175 267245 280265
rect 267335 280175 267425 280265
rect 267515 280175 267605 280265
rect 267695 280175 267785 280265
rect 267875 280175 267965 280265
rect 268055 280175 268145 280265
rect 268235 280175 268325 280265
rect 268415 280175 268505 280265
rect 268595 280175 268685 280265
rect 268775 280175 268865 280265
rect 268955 280175 269045 280265
rect 269135 280175 269225 280265
rect 269315 280175 269405 280265
rect 269495 280175 269585 280265
rect 269675 280175 269765 280265
rect 269855 280175 269945 280265
rect 270035 280175 270125 280265
rect 270215 280175 270305 280265
rect 270395 280175 270485 280265
rect 270575 280175 270665 280265
rect 270755 280175 270845 280265
rect 270935 280175 271025 280265
rect 271115 280175 271205 280265
rect 271295 280175 271385 280265
rect 271475 280175 271565 280265
rect 271655 280175 271745 280265
rect 271835 280175 271925 280265
rect 272015 280175 272105 280265
rect 272195 280175 272285 280265
rect 272375 280175 272465 280265
rect 272555 280175 272645 280265
rect 272735 280175 272825 280265
rect 272915 280175 273005 280265
rect 273095 280175 273185 280265
rect 273275 280175 273365 280265
rect 273455 280175 273545 280265
rect 273635 280175 273725 280265
rect 273815 280175 273905 280265
rect 273995 280175 274085 280265
rect 274175 280175 274265 280265
rect 274355 280175 274450 280265
rect 265350 280085 274450 280175
rect 265350 279995 265445 280085
rect 265535 279995 265625 280085
rect 265715 279995 265805 280085
rect 265895 279995 265985 280085
rect 266075 279995 266165 280085
rect 266255 279995 266345 280085
rect 266435 279995 266525 280085
rect 266615 279995 266705 280085
rect 266795 279995 266885 280085
rect 266975 279995 267065 280085
rect 267155 279995 267245 280085
rect 267335 279995 267425 280085
rect 267515 279995 267605 280085
rect 267695 279995 267785 280085
rect 267875 279995 267965 280085
rect 268055 279995 268145 280085
rect 268235 279995 268325 280085
rect 268415 279995 268505 280085
rect 268595 279995 268685 280085
rect 268775 279995 268865 280085
rect 268955 279995 269045 280085
rect 269135 279995 269225 280085
rect 269315 279995 269405 280085
rect 269495 279995 269585 280085
rect 269675 279995 269765 280085
rect 269855 279995 269945 280085
rect 270035 279995 270125 280085
rect 270215 279995 270305 280085
rect 270395 279995 270485 280085
rect 270575 279995 270665 280085
rect 270755 279995 270845 280085
rect 270935 279995 271025 280085
rect 271115 279995 271205 280085
rect 271295 279995 271385 280085
rect 271475 279995 271565 280085
rect 271655 279995 271745 280085
rect 271835 279995 271925 280085
rect 272015 279995 272105 280085
rect 272195 279995 272285 280085
rect 272375 279995 272465 280085
rect 272555 279995 272645 280085
rect 272735 279995 272825 280085
rect 272915 279995 273005 280085
rect 273095 279995 273185 280085
rect 273275 279995 273365 280085
rect 273455 279995 273545 280085
rect 273635 279995 273725 280085
rect 273815 279995 273905 280085
rect 273995 279995 274085 280085
rect 274175 279995 274265 280085
rect 274355 279995 274450 280085
rect 265350 279905 274450 279995
rect 265350 279815 265445 279905
rect 265535 279815 265625 279905
rect 265715 279815 265805 279905
rect 265895 279815 265985 279905
rect 266075 279815 266165 279905
rect 266255 279815 266345 279905
rect 266435 279815 266525 279905
rect 266615 279815 266705 279905
rect 266795 279815 266885 279905
rect 266975 279815 267065 279905
rect 267155 279815 267245 279905
rect 267335 279815 267425 279905
rect 267515 279815 267605 279905
rect 267695 279815 267785 279905
rect 267875 279815 267965 279905
rect 268055 279815 268145 279905
rect 268235 279815 268325 279905
rect 268415 279815 268505 279905
rect 268595 279815 268685 279905
rect 268775 279815 268865 279905
rect 268955 279815 269045 279905
rect 269135 279815 269225 279905
rect 269315 279815 269405 279905
rect 269495 279815 269585 279905
rect 269675 279815 269765 279905
rect 269855 279815 269945 279905
rect 270035 279815 270125 279905
rect 270215 279815 270305 279905
rect 270395 279815 270485 279905
rect 270575 279815 270665 279905
rect 270755 279815 270845 279905
rect 270935 279815 271025 279905
rect 271115 279815 271205 279905
rect 271295 279815 271385 279905
rect 271475 279815 271565 279905
rect 271655 279815 271745 279905
rect 271835 279815 271925 279905
rect 272015 279815 272105 279905
rect 272195 279815 272285 279905
rect 272375 279815 272465 279905
rect 272555 279815 272645 279905
rect 272735 279815 272825 279905
rect 272915 279815 273005 279905
rect 273095 279815 273185 279905
rect 273275 279815 273365 279905
rect 273455 279815 273545 279905
rect 273635 279815 273725 279905
rect 273815 279815 273905 279905
rect 273995 279815 274085 279905
rect 274175 279815 274265 279905
rect 274355 279815 274450 279905
rect 265350 279725 274450 279815
rect 265350 279635 265445 279725
rect 265535 279635 265625 279725
rect 265715 279635 265805 279725
rect 265895 279635 265985 279725
rect 266075 279635 266165 279725
rect 266255 279635 266345 279725
rect 266435 279635 266525 279725
rect 266615 279635 266705 279725
rect 266795 279635 266885 279725
rect 266975 279635 267065 279725
rect 267155 279635 267245 279725
rect 267335 279635 267425 279725
rect 267515 279635 267605 279725
rect 267695 279635 267785 279725
rect 267875 279635 267965 279725
rect 268055 279635 268145 279725
rect 268235 279635 268325 279725
rect 268415 279635 268505 279725
rect 268595 279635 268685 279725
rect 268775 279635 268865 279725
rect 268955 279635 269045 279725
rect 269135 279635 269225 279725
rect 269315 279635 269405 279725
rect 269495 279635 269585 279725
rect 269675 279635 269765 279725
rect 269855 279635 269945 279725
rect 270035 279635 270125 279725
rect 270215 279635 270305 279725
rect 270395 279635 270485 279725
rect 270575 279635 270665 279725
rect 270755 279635 270845 279725
rect 270935 279635 271025 279725
rect 271115 279635 271205 279725
rect 271295 279635 271385 279725
rect 271475 279635 271565 279725
rect 271655 279635 271745 279725
rect 271835 279635 271925 279725
rect 272015 279635 272105 279725
rect 272195 279635 272285 279725
rect 272375 279635 272465 279725
rect 272555 279635 272645 279725
rect 272735 279635 272825 279725
rect 272915 279635 273005 279725
rect 273095 279635 273185 279725
rect 273275 279635 273365 279725
rect 273455 279635 273545 279725
rect 273635 279635 273725 279725
rect 273815 279635 273905 279725
rect 273995 279635 274085 279725
rect 274175 279635 274265 279725
rect 274355 279635 274450 279725
rect 265350 279545 274450 279635
rect 265350 279455 265445 279545
rect 265535 279455 265625 279545
rect 265715 279455 265805 279545
rect 265895 279455 265985 279545
rect 266075 279455 266165 279545
rect 266255 279455 266345 279545
rect 266435 279455 266525 279545
rect 266615 279455 266705 279545
rect 266795 279455 266885 279545
rect 266975 279455 267065 279545
rect 267155 279455 267245 279545
rect 267335 279455 267425 279545
rect 267515 279455 267605 279545
rect 267695 279455 267785 279545
rect 267875 279455 267965 279545
rect 268055 279455 268145 279545
rect 268235 279455 268325 279545
rect 268415 279455 268505 279545
rect 268595 279455 268685 279545
rect 268775 279455 268865 279545
rect 268955 279455 269045 279545
rect 269135 279455 269225 279545
rect 269315 279455 269405 279545
rect 269495 279455 269585 279545
rect 269675 279455 269765 279545
rect 269855 279455 269945 279545
rect 270035 279455 270125 279545
rect 270215 279455 270305 279545
rect 270395 279455 270485 279545
rect 270575 279455 270665 279545
rect 270755 279455 270845 279545
rect 270935 279455 271025 279545
rect 271115 279455 271205 279545
rect 271295 279455 271385 279545
rect 271475 279455 271565 279545
rect 271655 279455 271745 279545
rect 271835 279455 271925 279545
rect 272015 279455 272105 279545
rect 272195 279455 272285 279545
rect 272375 279455 272465 279545
rect 272555 279455 272645 279545
rect 272735 279455 272825 279545
rect 272915 279455 273005 279545
rect 273095 279455 273185 279545
rect 273275 279455 273365 279545
rect 273455 279455 273545 279545
rect 273635 279455 273725 279545
rect 273815 279455 273905 279545
rect 273995 279455 274085 279545
rect 274175 279455 274265 279545
rect 274355 279455 274450 279545
rect 265350 279350 274450 279455
rect 189986 275750 248800 276050
rect 189989 271238 190289 275750
rect 190630 275156 280250 275450
rect 190630 275150 191996 275156
rect 192575 275150 280250 275156
rect 190633 271216 190933 275150
rect 192575 274828 279650 274850
rect 192098 274555 279650 274828
rect 192098 274550 193556 274555
rect 193959 274550 279650 274555
rect 192100 274300 192400 274550
rect 192100 274250 192394 274300
rect 192098 273950 192394 274250
rect 192100 273650 192394 273950
rect 192098 273350 192394 273650
rect 192100 273050 192394 273350
rect 192098 272750 192394 273050
rect 192100 272450 192394 272750
rect 192098 272150 192394 272450
rect 192100 271850 192394 272150
rect 192098 271550 192394 271850
rect 192100 271200 192394 271550
rect 193604 274250 193900 274264
rect 193604 273950 279050 274250
rect 193604 273725 193900 273950
rect 193604 271200 193888 273725
rect 194801 273350 278450 273650
rect 194801 273345 195100 273350
rect 194807 273161 195100 273345
rect 194807 271200 195098 273161
rect 196301 272750 277850 273050
rect 196301 272515 196600 272750
rect 196301 271934 196597 272515
rect 199597 272150 277250 272450
rect 196301 271401 196592 271934
rect 199600 271863 199900 272150
rect 199600 271850 199899 271863
rect 199597 271550 199899 271850
rect 201091 271550 276650 271850
rect 196301 271200 196597 271401
rect 199600 271300 199899 271550
rect 199600 271200 199900 271300
rect 201100 271200 201400 271550
rect 99400 200350 103650 200750
rect 104250 194465 104650 194550
rect 104250 194375 104315 194465
rect 104405 194375 104495 194465
rect 104585 194375 104650 194465
rect 104250 194285 104650 194375
rect 104250 194195 104315 194285
rect 104405 194195 104495 194285
rect 104585 194195 104650 194285
rect 104250 194150 104650 194195
rect 102150 194105 104650 194150
rect 102150 194015 104315 194105
rect 104405 194015 104495 194105
rect 104585 194015 104650 194105
rect 102150 193925 104650 194015
rect 102150 193835 104315 193925
rect 104405 193835 104495 193925
rect 104585 193835 104650 193925
rect 102150 193750 104650 193835
rect 100050 184925 100350 185050
rect 100050 184835 100155 184925
rect 100245 184835 100350 184925
rect 100050 184745 100350 184835
rect 100050 184700 100155 184745
rect 99400 184655 100155 184700
rect 100245 184655 100350 184745
rect 99400 184565 100350 184655
rect 99400 184475 100155 184565
rect 100245 184475 100350 184565
rect 99400 184350 100350 184475
rect 99400 179370 100950 179500
rect 99400 179280 100400 179370
rect 100490 179280 100580 179370
rect 100670 179280 100760 179370
rect 100850 179280 100950 179370
rect 99400 179150 100950 179280
rect 99400 163370 101550 163500
rect 99400 163280 100975 163370
rect 101065 163280 101155 163370
rect 101245 163280 101335 163370
rect 101425 163280 101550 163370
rect 99400 163150 101550 163280
rect 99400 147370 101200 147500
rect 99400 147280 100485 147370
rect 100575 147280 100665 147370
rect 100755 147280 100845 147370
rect 100935 147280 101025 147370
rect 101115 147280 101200 147370
rect 99400 147150 101200 147280
rect 99400 131485 101300 131550
rect 99400 131395 100610 131485
rect 100700 131395 100790 131485
rect 100880 131395 100970 131485
rect 101060 131395 101150 131485
rect 101240 131395 101300 131485
rect 99400 131305 101300 131395
rect 99400 131215 100610 131305
rect 100700 131215 100790 131305
rect 100880 131215 100970 131305
rect 101060 131215 101150 131305
rect 101240 131215 101300 131305
rect 99400 131150 101300 131215
rect 99400 115370 101450 115500
rect 99400 115280 100875 115370
rect 100965 115280 101055 115370
rect 101145 115280 101235 115370
rect 101325 115280 101450 115370
rect 99400 115150 101450 115280
rect 102152 101250 102448 193750
rect 104250 190565 104650 190650
rect 104250 190475 104315 190565
rect 104405 190475 104495 190565
rect 104585 190475 104650 190565
rect 104250 190385 104650 190475
rect 104250 190295 104315 190385
rect 104405 190295 104495 190385
rect 104585 190295 104650 190385
rect 104250 190250 104650 190295
rect 102750 190205 104650 190250
rect 102750 190115 104315 190205
rect 104405 190115 104495 190205
rect 104585 190115 104650 190205
rect 102750 190025 104650 190115
rect 102750 189935 104315 190025
rect 104405 189935 104495 190025
rect 104585 189935 104650 190025
rect 102750 189850 104650 189935
rect 102750 101850 103050 189850
rect 104250 182165 104650 182250
rect 104250 182075 104315 182165
rect 104405 182075 104495 182165
rect 104585 182075 104650 182165
rect 104250 181985 104650 182075
rect 104250 181895 104315 181985
rect 104405 181895 104495 181985
rect 104585 181895 104650 181985
rect 104250 181850 104650 181895
rect 103350 181805 104650 181850
rect 103350 181715 104315 181805
rect 104405 181715 104495 181805
rect 104585 181715 104650 181805
rect 103350 181625 104650 181715
rect 103350 181535 104315 181625
rect 104405 181535 104495 181625
rect 104585 181535 104650 181625
rect 103350 181450 104650 181535
rect 103350 102450 103650 181450
rect 276350 168800 276650 271550
rect 276950 184800 277250 272150
rect 277550 200800 277850 272750
rect 278150 227600 278450 273350
rect 278750 232800 279050 273950
rect 279350 248800 279650 274550
rect 279950 264800 280250 275150
rect 279950 264440 280550 264800
rect 279350 248450 280550 248800
rect 278750 232450 280550 232800
rect 278150 227250 280550 227600
rect 277550 200450 280550 200800
rect 276950 184450 280550 184800
rect 276350 168450 280550 168800
rect 279050 163940 279350 164000
rect 279050 163850 279155 163940
rect 279245 163850 279350 163940
rect 279050 163760 279350 163850
rect 279050 163670 279155 163760
rect 279245 163670 279350 163760
rect 279050 163600 279350 163670
rect 279050 163580 280550 163600
rect 279050 163490 279155 163580
rect 279245 163490 280550 163580
rect 279050 163400 280550 163490
rect 279050 163310 279155 163400
rect 279245 163310 280550 163400
rect 279050 163250 280550 163310
rect 278450 137025 278750 137150
rect 278450 136935 278555 137025
rect 278645 136935 278750 137025
rect 278450 136845 278750 136935
rect 278450 136755 278555 136845
rect 278645 136800 278750 136845
rect 278645 136755 280550 136800
rect 278450 136665 280550 136755
rect 278450 136575 278555 136665
rect 278645 136575 280550 136665
rect 278450 136450 280550 136575
rect 277850 131825 278150 131950
rect 277850 131735 277955 131825
rect 278045 131735 278150 131825
rect 277850 131645 278150 131735
rect 277850 131555 277955 131645
rect 278045 131600 278150 131645
rect 278045 131555 280550 131600
rect 277850 131465 280550 131555
rect 277850 131375 277955 131465
rect 278045 131375 280550 131465
rect 277850 131250 280550 131375
rect 277250 115800 277550 115900
rect 277250 115710 277355 115800
rect 277445 115710 277550 115800
rect 277250 115620 277550 115710
rect 277250 115530 277355 115620
rect 277445 115600 277550 115620
rect 277445 115530 280550 115600
rect 277250 115440 280550 115530
rect 277250 115350 277355 115440
rect 277445 115350 280550 115440
rect 277250 115250 280550 115350
rect 103350 102150 179600 102450
rect 102750 101550 152800 101850
rect 102150 100950 136800 101250
rect 131250 100525 131600 100600
rect 106550 100355 113150 100450
rect 106550 100265 106655 100355
rect 106745 100265 106835 100355
rect 106925 100265 107015 100355
rect 107105 100265 107195 100355
rect 107285 100265 107375 100355
rect 107465 100265 107555 100355
rect 107645 100265 107735 100355
rect 107825 100265 107915 100355
rect 108005 100265 108095 100355
rect 108185 100265 108275 100355
rect 108365 100265 108455 100355
rect 108545 100265 108635 100355
rect 108725 100265 108815 100355
rect 108905 100265 108995 100355
rect 109085 100265 109175 100355
rect 109265 100265 109355 100355
rect 109445 100265 109535 100355
rect 109625 100265 109715 100355
rect 109805 100265 109895 100355
rect 109985 100265 110075 100355
rect 110165 100265 110255 100355
rect 110345 100265 110435 100355
rect 110525 100265 110615 100355
rect 110705 100265 110795 100355
rect 110885 100265 110975 100355
rect 111065 100265 111155 100355
rect 111245 100265 111335 100355
rect 111425 100265 111515 100355
rect 111605 100265 111695 100355
rect 111785 100265 111875 100355
rect 111965 100265 112055 100355
rect 112145 100265 112235 100355
rect 112325 100265 112415 100355
rect 112505 100265 112595 100355
rect 112685 100265 112775 100355
rect 112865 100265 112955 100355
rect 113045 100265 113150 100355
rect 106550 100175 113150 100265
rect 106550 100085 106655 100175
rect 106745 100085 106835 100175
rect 106925 100085 107015 100175
rect 107105 100085 107195 100175
rect 107285 100085 107375 100175
rect 107465 100085 107555 100175
rect 107645 100085 107735 100175
rect 107825 100085 107915 100175
rect 108005 100085 108095 100175
rect 108185 100085 108275 100175
rect 108365 100085 108455 100175
rect 108545 100085 108635 100175
rect 108725 100085 108815 100175
rect 108905 100085 108995 100175
rect 109085 100085 109175 100175
rect 109265 100085 109355 100175
rect 109445 100085 109535 100175
rect 109625 100085 109715 100175
rect 109805 100085 109895 100175
rect 109985 100085 110075 100175
rect 110165 100085 110255 100175
rect 110345 100085 110435 100175
rect 110525 100085 110615 100175
rect 110705 100085 110795 100175
rect 110885 100085 110975 100175
rect 111065 100085 111155 100175
rect 111245 100085 111335 100175
rect 111425 100085 111515 100175
rect 111605 100085 111695 100175
rect 111785 100085 111875 100175
rect 111965 100085 112055 100175
rect 112145 100085 112235 100175
rect 112325 100085 112415 100175
rect 112505 100085 112595 100175
rect 112685 100085 112775 100175
rect 112865 100085 112955 100175
rect 113045 100085 113150 100175
rect 106550 99995 113150 100085
rect 106550 99905 106655 99995
rect 106745 99905 106835 99995
rect 106925 99905 107015 99995
rect 107105 99905 107195 99995
rect 107285 99905 107375 99995
rect 107465 99905 107555 99995
rect 107645 99905 107735 99995
rect 107825 99905 107915 99995
rect 108005 99905 108095 99995
rect 108185 99905 108275 99995
rect 108365 99905 108455 99995
rect 108545 99905 108635 99995
rect 108725 99905 108815 99995
rect 108905 99905 108995 99995
rect 109085 99905 109175 99995
rect 109265 99905 109355 99995
rect 109445 99905 109535 99995
rect 109625 99905 109715 99995
rect 109805 99905 109895 99995
rect 109985 99905 110075 99995
rect 110165 99905 110255 99995
rect 110345 99905 110435 99995
rect 110525 99905 110615 99995
rect 110705 99905 110795 99995
rect 110885 99905 110975 99995
rect 111065 99905 111155 99995
rect 111245 99905 111335 99995
rect 111425 99905 111515 99995
rect 111605 99905 111695 99995
rect 111785 99905 111875 99995
rect 111965 99905 112055 99995
rect 112145 99905 112235 99995
rect 112325 99905 112415 99995
rect 112505 99905 112595 99995
rect 112685 99905 112775 99995
rect 112865 99905 112955 99995
rect 113045 99905 113150 99995
rect 106550 99815 113150 99905
rect 106550 99725 106655 99815
rect 106745 99725 106835 99815
rect 106925 99725 107015 99815
rect 107105 99725 107195 99815
rect 107285 99725 107375 99815
rect 107465 99725 107555 99815
rect 107645 99725 107735 99815
rect 107825 99725 107915 99815
rect 108005 99725 108095 99815
rect 108185 99725 108275 99815
rect 108365 99725 108455 99815
rect 108545 99725 108635 99815
rect 108725 99725 108815 99815
rect 108905 99725 108995 99815
rect 109085 99725 109175 99815
rect 109265 99725 109355 99815
rect 109445 99725 109535 99815
rect 109625 99725 109715 99815
rect 109805 99725 109895 99815
rect 109985 99725 110075 99815
rect 110165 99725 110255 99815
rect 110345 99725 110435 99815
rect 110525 99725 110615 99815
rect 110705 99725 110795 99815
rect 110885 99725 110975 99815
rect 111065 99725 111155 99815
rect 111245 99725 111335 99815
rect 111425 99725 111515 99815
rect 111605 99725 111695 99815
rect 111785 99725 111875 99815
rect 111965 99725 112055 99815
rect 112145 99725 112235 99815
rect 112325 99725 112415 99815
rect 112505 99725 112595 99815
rect 112685 99725 112775 99815
rect 112865 99725 112955 99815
rect 113045 99725 113150 99815
rect 106550 99635 113150 99725
rect 106550 99545 106655 99635
rect 106745 99545 106835 99635
rect 106925 99545 107015 99635
rect 107105 99545 107195 99635
rect 107285 99545 107375 99635
rect 107465 99545 107555 99635
rect 107645 99545 107735 99635
rect 107825 99545 107915 99635
rect 108005 99545 108095 99635
rect 108185 99545 108275 99635
rect 108365 99545 108455 99635
rect 108545 99545 108635 99635
rect 108725 99545 108815 99635
rect 108905 99545 108995 99635
rect 109085 99545 109175 99635
rect 109265 99545 109355 99635
rect 109445 99545 109535 99635
rect 109625 99545 109715 99635
rect 109805 99545 109895 99635
rect 109985 99545 110075 99635
rect 110165 99545 110255 99635
rect 110345 99545 110435 99635
rect 110525 99545 110615 99635
rect 110705 99545 110795 99635
rect 110885 99545 110975 99635
rect 111065 99545 111155 99635
rect 111245 99545 111335 99635
rect 111425 99545 111515 99635
rect 111605 99545 111695 99635
rect 111785 99545 111875 99635
rect 111965 99545 112055 99635
rect 112145 99545 112235 99635
rect 112325 99545 112415 99635
rect 112505 99545 112595 99635
rect 112685 99545 112775 99635
rect 112865 99545 112955 99635
rect 113045 99545 113150 99635
rect 106550 99450 113150 99545
rect 131250 100435 131380 100525
rect 131470 100435 131600 100525
rect 131250 100345 131600 100435
rect 131250 100255 131380 100345
rect 131470 100255 131600 100345
rect 131250 100165 131600 100255
rect 131250 100075 131380 100165
rect 131470 100075 131600 100165
rect 131250 99400 131600 100075
rect 136450 99400 136800 100950
rect 152450 99400 152800 101550
rect 179250 99400 179600 102150
rect 185150 100850 185450 102350
rect 184450 100550 185450 100850
rect 184450 99400 184800 100550
rect 208550 100250 208850 102450
rect 259250 102445 260000 102550
rect 259250 102355 259310 102445
rect 259400 102355 259490 102445
rect 259580 102355 259670 102445
rect 259760 102355 259850 102445
rect 259940 102355 260000 102445
rect 259250 102250 260000 102355
rect 208550 99950 211600 100250
rect 211250 99400 211600 99950
rect 259250 99400 259650 102250
rect 265350 100305 274450 100450
rect 265350 100215 265445 100305
rect 265535 100215 265625 100305
rect 265715 100215 265805 100305
rect 265895 100215 265985 100305
rect 266075 100215 266165 100305
rect 266255 100215 266345 100305
rect 266435 100215 266525 100305
rect 266615 100215 266705 100305
rect 266795 100215 266885 100305
rect 266975 100215 267065 100305
rect 267155 100215 267245 100305
rect 267335 100215 267425 100305
rect 267515 100215 267605 100305
rect 267695 100215 267785 100305
rect 267875 100215 267965 100305
rect 268055 100215 268145 100305
rect 268235 100215 268325 100305
rect 268415 100215 268505 100305
rect 268595 100215 268685 100305
rect 268775 100215 268865 100305
rect 268955 100215 269045 100305
rect 269135 100215 269225 100305
rect 269315 100215 269405 100305
rect 269495 100215 269585 100305
rect 269675 100215 269765 100305
rect 269855 100215 269945 100305
rect 270035 100215 270125 100305
rect 270215 100215 270305 100305
rect 270395 100215 270485 100305
rect 270575 100215 270665 100305
rect 270755 100215 270845 100305
rect 270935 100215 271025 100305
rect 271115 100215 271205 100305
rect 271295 100215 271385 100305
rect 271475 100215 271565 100305
rect 271655 100215 271745 100305
rect 271835 100215 271925 100305
rect 272015 100215 272105 100305
rect 272195 100215 272285 100305
rect 272375 100215 272465 100305
rect 272555 100215 272645 100305
rect 272735 100215 272825 100305
rect 272915 100215 273005 100305
rect 273095 100215 273185 100305
rect 273275 100215 273365 100305
rect 273455 100215 273545 100305
rect 273635 100215 273725 100305
rect 273815 100215 273905 100305
rect 273995 100215 274085 100305
rect 274175 100215 274265 100305
rect 274355 100215 274450 100305
rect 265350 100125 274450 100215
rect 265350 100035 265445 100125
rect 265535 100035 265625 100125
rect 265715 100035 265805 100125
rect 265895 100035 265985 100125
rect 266075 100035 266165 100125
rect 266255 100035 266345 100125
rect 266435 100035 266525 100125
rect 266615 100035 266705 100125
rect 266795 100035 266885 100125
rect 266975 100035 267065 100125
rect 267155 100035 267245 100125
rect 267335 100035 267425 100125
rect 267515 100035 267605 100125
rect 267695 100035 267785 100125
rect 267875 100035 267965 100125
rect 268055 100035 268145 100125
rect 268235 100035 268325 100125
rect 268415 100035 268505 100125
rect 268595 100035 268685 100125
rect 268775 100035 268865 100125
rect 268955 100035 269045 100125
rect 269135 100035 269225 100125
rect 269315 100035 269405 100125
rect 269495 100035 269585 100125
rect 269675 100035 269765 100125
rect 269855 100035 269945 100125
rect 270035 100035 270125 100125
rect 270215 100035 270305 100125
rect 270395 100035 270485 100125
rect 270575 100035 270665 100125
rect 270755 100035 270845 100125
rect 270935 100035 271025 100125
rect 271115 100035 271205 100125
rect 271295 100035 271385 100125
rect 271475 100035 271565 100125
rect 271655 100035 271745 100125
rect 271835 100035 271925 100125
rect 272015 100035 272105 100125
rect 272195 100035 272285 100125
rect 272375 100035 272465 100125
rect 272555 100035 272645 100125
rect 272735 100035 272825 100125
rect 272915 100035 273005 100125
rect 273095 100035 273185 100125
rect 273275 100035 273365 100125
rect 273455 100035 273545 100125
rect 273635 100035 273725 100125
rect 273815 100035 273905 100125
rect 273995 100035 274085 100125
rect 274175 100035 274265 100125
rect 274355 100035 274450 100125
rect 265350 99945 274450 100035
rect 265350 99855 265445 99945
rect 265535 99855 265625 99945
rect 265715 99855 265805 99945
rect 265895 99855 265985 99945
rect 266075 99855 266165 99945
rect 266255 99855 266345 99945
rect 266435 99855 266525 99945
rect 266615 99855 266705 99945
rect 266795 99855 266885 99945
rect 266975 99855 267065 99945
rect 267155 99855 267245 99945
rect 267335 99855 267425 99945
rect 267515 99855 267605 99945
rect 267695 99855 267785 99945
rect 267875 99855 267965 99945
rect 268055 99855 268145 99945
rect 268235 99855 268325 99945
rect 268415 99855 268505 99945
rect 268595 99855 268685 99945
rect 268775 99855 268865 99945
rect 268955 99855 269045 99945
rect 269135 99855 269225 99945
rect 269315 99855 269405 99945
rect 269495 99855 269585 99945
rect 269675 99855 269765 99945
rect 269855 99855 269945 99945
rect 270035 99855 270125 99945
rect 270215 99855 270305 99945
rect 270395 99855 270485 99945
rect 270575 99855 270665 99945
rect 270755 99855 270845 99945
rect 270935 99855 271025 99945
rect 271115 99855 271205 99945
rect 271295 99855 271385 99945
rect 271475 99855 271565 99945
rect 271655 99855 271745 99945
rect 271835 99855 271925 99945
rect 272015 99855 272105 99945
rect 272195 99855 272285 99945
rect 272375 99855 272465 99945
rect 272555 99855 272645 99945
rect 272735 99855 272825 99945
rect 272915 99855 273005 99945
rect 273095 99855 273185 99945
rect 273275 99855 273365 99945
rect 273455 99855 273545 99945
rect 273635 99855 273725 99945
rect 273815 99855 273905 99945
rect 273995 99855 274085 99945
rect 274175 99855 274265 99945
rect 274355 99855 274450 99945
rect 265350 99765 274450 99855
rect 265350 99675 265445 99765
rect 265535 99675 265625 99765
rect 265715 99675 265805 99765
rect 265895 99675 265985 99765
rect 266075 99675 266165 99765
rect 266255 99675 266345 99765
rect 266435 99675 266525 99765
rect 266615 99675 266705 99765
rect 266795 99675 266885 99765
rect 266975 99675 267065 99765
rect 267155 99675 267245 99765
rect 267335 99675 267425 99765
rect 267515 99675 267605 99765
rect 267695 99675 267785 99765
rect 267875 99675 267965 99765
rect 268055 99675 268145 99765
rect 268235 99675 268325 99765
rect 268415 99675 268505 99765
rect 268595 99675 268685 99765
rect 268775 99675 268865 99765
rect 268955 99675 269045 99765
rect 269135 99675 269225 99765
rect 269315 99675 269405 99765
rect 269495 99675 269585 99765
rect 269675 99675 269765 99765
rect 269855 99675 269945 99765
rect 270035 99675 270125 99765
rect 270215 99675 270305 99765
rect 270395 99675 270485 99765
rect 270575 99675 270665 99765
rect 270755 99675 270845 99765
rect 270935 99675 271025 99765
rect 271115 99675 271205 99765
rect 271295 99675 271385 99765
rect 271475 99675 271565 99765
rect 271655 99675 271745 99765
rect 271835 99675 271925 99765
rect 272015 99675 272105 99765
rect 272195 99675 272285 99765
rect 272375 99675 272465 99765
rect 272555 99675 272645 99765
rect 272735 99675 272825 99765
rect 272915 99675 273005 99765
rect 273095 99675 273185 99765
rect 273275 99675 273365 99765
rect 273455 99675 273545 99765
rect 273635 99675 273725 99765
rect 273815 99675 273905 99765
rect 273995 99675 274085 99765
rect 274175 99675 274265 99765
rect 274355 99675 274450 99765
rect 265350 99585 274450 99675
rect 265350 99495 265445 99585
rect 265535 99495 265625 99585
rect 265715 99495 265805 99585
rect 265895 99495 265985 99585
rect 266075 99495 266165 99585
rect 266255 99495 266345 99585
rect 266435 99495 266525 99585
rect 266615 99495 266705 99585
rect 266795 99495 266885 99585
rect 266975 99495 267065 99585
rect 267155 99495 267245 99585
rect 267335 99495 267425 99585
rect 267515 99495 267605 99585
rect 267695 99495 267785 99585
rect 267875 99495 267965 99585
rect 268055 99495 268145 99585
rect 268235 99495 268325 99585
rect 268415 99495 268505 99585
rect 268595 99495 268685 99585
rect 268775 99495 268865 99585
rect 268955 99495 269045 99585
rect 269135 99495 269225 99585
rect 269315 99495 269405 99585
rect 269495 99495 269585 99585
rect 269675 99495 269765 99585
rect 269855 99495 269945 99585
rect 270035 99495 270125 99585
rect 270215 99495 270305 99585
rect 270395 99495 270485 99585
rect 270575 99495 270665 99585
rect 270755 99495 270845 99585
rect 270935 99495 271025 99585
rect 271115 99495 271205 99585
rect 271295 99495 271385 99585
rect 271475 99495 271565 99585
rect 271655 99495 271745 99585
rect 271835 99495 271925 99585
rect 272015 99495 272105 99585
rect 272195 99495 272285 99585
rect 272375 99495 272465 99585
rect 272555 99495 272645 99585
rect 272735 99495 272825 99585
rect 272915 99495 273005 99585
rect 273095 99495 273185 99585
rect 273275 99495 273365 99585
rect 273455 99495 273545 99585
rect 273635 99495 273725 99585
rect 273815 99495 273905 99585
rect 273995 99495 274085 99585
rect 274175 99495 274265 99585
rect 274355 99495 274450 99585
rect 265350 99350 274450 99495
<< m3contact >>
rect 104315 194375 104405 194465
rect 104495 194375 104585 194465
rect 104315 194195 104405 194285
rect 104495 194195 104585 194285
rect 104315 194015 104405 194105
rect 104495 194015 104585 194105
rect 104315 193835 104405 193925
rect 104495 193835 104585 193925
rect 100155 184835 100245 184925
rect 100155 184655 100245 184745
rect 100155 184475 100245 184565
rect 100400 179280 100490 179370
rect 100580 179280 100670 179370
rect 100760 179280 100850 179370
rect 100975 163280 101065 163370
rect 101155 163280 101245 163370
rect 101335 163280 101425 163370
rect 100485 147280 100575 147370
rect 100665 147280 100755 147370
rect 100845 147280 100935 147370
rect 101025 147280 101115 147370
rect 100610 131395 100700 131485
rect 100790 131395 100880 131485
rect 100970 131395 101060 131485
rect 101150 131395 101240 131485
rect 100610 131215 100700 131305
rect 100790 131215 100880 131305
rect 100970 131215 101060 131305
rect 101150 131215 101240 131305
rect 100875 115280 100965 115370
rect 101055 115280 101145 115370
rect 101235 115280 101325 115370
rect 104315 190475 104405 190565
rect 104495 190475 104585 190565
rect 104315 190295 104405 190385
rect 104495 190295 104585 190385
rect 104315 190115 104405 190205
rect 104495 190115 104585 190205
rect 104315 189935 104405 190025
rect 104495 189935 104585 190025
rect 104315 182075 104405 182165
rect 104495 182075 104585 182165
rect 104315 181895 104405 181985
rect 104495 181895 104585 181985
rect 104315 181715 104405 181805
rect 104495 181715 104585 181805
rect 104315 181535 104405 181625
rect 104495 181535 104585 181625
rect 279155 163850 279245 163940
rect 279155 163670 279245 163760
rect 279155 163490 279245 163580
rect 279155 163310 279245 163400
rect 278555 136935 278645 137025
rect 278555 136755 278645 136845
rect 278555 136575 278645 136665
rect 277955 131735 278045 131825
rect 277955 131555 278045 131645
rect 277955 131375 278045 131465
rect 277355 115710 277445 115800
rect 277355 115530 277445 115620
rect 277355 115350 277445 115440
rect 131380 100435 131470 100525
rect 131380 100255 131470 100345
rect 131380 100075 131470 100165
rect 259310 102355 259400 102445
rect 259490 102355 259580 102445
rect 259670 102355 259760 102445
rect 259850 102355 259940 102445
<< metal3 >>
rect 100050 269255 104450 269350
rect 100050 269135 105410 269255
rect 100050 269050 104450 269135
rect 100050 184925 100350 269050
rect 100050 184835 100155 184925
rect 100245 184835 100350 184925
rect 100050 184745 100350 184835
rect 100050 184655 100155 184745
rect 100245 184655 100350 184745
rect 100050 184565 100350 184655
rect 100050 184475 100155 184565
rect 100245 184475 100350 184565
rect 100050 184350 100350 184475
rect 100650 242150 104350 242450
rect 100650 179500 100950 242150
rect 100300 179370 100950 179500
rect 100300 179280 100400 179370
rect 100490 179280 100580 179370
rect 100670 179280 100760 179370
rect 100850 179280 100950 179370
rect 100300 179150 100950 179280
rect 101250 241450 104350 241750
rect 101250 163500 101550 241450
rect 100850 163370 101550 163500
rect 100850 163280 100975 163370
rect 101065 163280 101155 163370
rect 101245 163280 101335 163370
rect 101425 163280 101550 163370
rect 100850 163150 101550 163280
rect 101850 233350 104450 233650
rect 101850 147500 102150 233350
rect 100400 147370 102150 147500
rect 100400 147280 100485 147370
rect 100575 147280 100665 147370
rect 100755 147280 100845 147370
rect 100935 147280 101025 147370
rect 101115 147280 102150 147370
rect 100400 147150 102150 147280
rect 102450 221650 104350 221950
rect 102450 131550 102750 221650
rect 100550 131485 102750 131550
rect 100550 131395 100610 131485
rect 100700 131395 100790 131485
rect 100880 131395 100970 131485
rect 101060 131395 101150 131485
rect 101240 131395 102750 131485
rect 100550 131305 102750 131395
rect 100550 131215 100610 131305
rect 100700 131215 100790 131305
rect 100880 131215 100970 131305
rect 101060 131215 101150 131305
rect 101240 131215 102750 131305
rect 100550 131150 102750 131215
rect 103050 210750 104350 211150
rect 103050 115500 103350 210750
rect 100750 115370 103350 115500
rect 100750 115280 100875 115370
rect 100965 115280 101055 115370
rect 101145 115280 101235 115370
rect 101325 115280 103350 115370
rect 100750 115150 103350 115280
rect 103650 209850 104350 210250
rect 276150 209850 279350 210250
rect 103650 101550 103950 209850
rect 276150 205950 278750 206350
rect 276150 202050 278150 202450
rect 104250 194465 104650 194550
rect 104250 194375 104315 194465
rect 104405 194375 104495 194465
rect 104585 194375 104650 194465
rect 104250 194285 104650 194375
rect 104250 194195 104315 194285
rect 104405 194195 104495 194285
rect 104585 194195 104650 194285
rect 104250 194105 104650 194195
rect 104250 194015 104315 194105
rect 104405 194015 104495 194105
rect 104585 194015 104650 194105
rect 104250 193925 104650 194015
rect 104250 193835 104315 193925
rect 104405 193835 104495 193925
rect 104585 193835 104650 193925
rect 104250 193750 104650 193835
rect 276150 193650 277550 194050
rect 104250 190565 104650 190650
rect 104250 190475 104315 190565
rect 104405 190475 104495 190565
rect 104585 190475 104650 190565
rect 104250 190385 104650 190475
rect 104250 190295 104315 190385
rect 104405 190295 104495 190385
rect 104585 190295 104650 190385
rect 104250 190205 104650 190295
rect 104250 190115 104315 190205
rect 104405 190115 104495 190205
rect 104585 190115 104650 190205
rect 104250 190025 104650 190115
rect 104250 189935 104315 190025
rect 104405 189935 104495 190025
rect 104585 189935 104650 190025
rect 104250 189850 104650 189935
rect 104250 182165 104650 182250
rect 104250 182075 104315 182165
rect 104405 182075 104495 182165
rect 104585 182075 104650 182165
rect 104250 181985 104650 182075
rect 104250 181895 104315 181985
rect 104405 181895 104495 181985
rect 104585 181895 104650 181985
rect 104250 181805 104650 181895
rect 104250 181715 104315 181805
rect 104405 181715 104495 181805
rect 104585 181715 104650 181805
rect 104250 181625 104650 181715
rect 104250 181535 104315 181625
rect 104405 181535 104495 181625
rect 104585 181535 104650 181625
rect 104250 181450 104650 181535
rect 276150 178950 276950 179350
rect 276650 102550 276950 178950
rect 277250 115800 277550 193650
rect 277850 131825 278150 202050
rect 278450 137025 278750 205950
rect 279050 163940 279350 209850
rect 279050 163850 279155 163940
rect 279245 163850 279350 163940
rect 279050 163760 279350 163850
rect 279050 163670 279155 163760
rect 279245 163670 279350 163760
rect 279050 163580 279350 163670
rect 279050 163490 279155 163580
rect 279245 163490 279350 163580
rect 279050 163400 279350 163490
rect 279050 163310 279155 163400
rect 279245 163310 279350 163400
rect 279050 163250 279350 163310
rect 278450 136935 278555 137025
rect 278645 136935 278750 137025
rect 278450 136845 278750 136935
rect 278450 136755 278555 136845
rect 278645 136755 278750 136845
rect 278450 136665 278750 136755
rect 278450 136575 278555 136665
rect 278645 136575 278750 136665
rect 278450 136450 278750 136575
rect 277850 131735 277955 131825
rect 278045 131735 278150 131825
rect 277850 131645 278150 131735
rect 277850 131555 277955 131645
rect 278045 131555 278150 131645
rect 277850 131465 278150 131555
rect 277850 131375 277955 131465
rect 278045 131375 278150 131465
rect 277850 131250 278150 131375
rect 277250 115710 277355 115800
rect 277445 115710 277550 115800
rect 277250 115620 277550 115710
rect 277250 115530 277355 115620
rect 277445 115530 277550 115620
rect 277250 115440 277550 115530
rect 277250 115350 277355 115440
rect 277445 115350 277550 115440
rect 277250 115250 277550 115350
rect 259250 102445 276950 102550
rect 259250 102355 259310 102445
rect 259400 102355 259490 102445
rect 259580 102355 259670 102445
rect 259760 102355 259850 102445
rect 259940 102355 276950 102445
rect 259250 102250 276950 102355
rect 103650 101250 131600 101550
rect 131250 100525 131600 101250
rect 131250 100435 131380 100525
rect 131470 100435 131600 100525
rect 131250 100345 131600 100435
rect 131250 100255 131380 100345
rect 131470 100255 131600 100345
rect 131250 100165 131600 100255
rect 131250 100075 131380 100165
rect 131470 100075 131600 100165
rect 131250 100000 131600 100075
<< comment >>
rect 0 0 380000 380000
<< end >>

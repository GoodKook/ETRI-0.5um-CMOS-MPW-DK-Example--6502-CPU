magic
tech scmos
magscale 1 2
timestamp 1709120482
<< checkpaint >>
rect 2068 11288 2155 11289
rect -103 11144 11446 11288
rect -106 11056 11446 11144
rect -103 9355 11446 11056
rect -107 9324 11446 9355
rect -108 9217 11446 9324
rect -103 8764 11446 9217
rect -107 8676 11446 8764
rect -103 7984 11446 8676
rect -107 7896 11446 7984
rect -103 7263 11446 7896
rect -107 7156 11446 7263
rect -105 7116 11446 7156
rect -103 6164 11446 7116
rect -107 6076 11446 6164
rect -103 5904 11446 6076
rect -106 5816 11446 5904
rect -103 5344 11446 5816
rect -105 5256 11446 5344
rect -103 -64 11446 5256
<< metal1 >>
rect -63 10938 -3 11198
rect 11310 11182 11403 11198
rect 9087 11117 9173 11123
rect 3387 11037 3453 11043
rect 6747 11037 6913 11043
rect -63 10922 30 10938
rect 347 10933 350 10947
rect -63 10418 -3 10922
rect 7367 10837 7473 10843
rect 7087 10817 7193 10823
rect 7467 10817 7533 10823
rect 8267 10817 8453 10823
rect 7367 10797 7413 10803
rect 6227 10737 6293 10743
rect 6367 10737 6393 10743
rect 10807 10737 10993 10743
rect 11343 10678 11403 11182
rect 11310 10662 11403 10678
rect 2467 10597 2473 10603
rect 2487 10597 2593 10603
rect 9007 10597 9033 10603
rect 5667 10577 5753 10583
rect 9547 10537 9573 10543
rect 2487 10517 2693 10523
rect 3427 10517 3553 10523
rect 4487 10517 4593 10523
rect 4707 10517 4873 10523
rect 6767 10517 6853 10523
rect 8627 10517 8773 10523
rect 10727 10517 10773 10523
rect -63 10402 30 10418
rect -63 9898 -3 10402
rect 3097 10383 3103 10403
rect 3067 10377 3103 10383
rect 4387 10317 4473 10323
rect 1487 10297 1593 10303
rect 8427 10297 8533 10303
rect 9207 10297 9413 10303
rect 3487 10277 3593 10283
rect 8007 10277 8133 10283
rect 5233 10243 5247 10253
rect 5233 10240 5353 10243
rect 5237 10237 5353 10240
rect 9327 10237 9353 10243
rect 207 10217 353 10223
rect 5267 10217 5353 10223
rect 5487 10217 5613 10223
rect 7747 10217 7793 10223
rect 9347 10217 9393 10223
rect 4407 10197 4433 10203
rect 11343 10158 11403 10662
rect 11310 10142 11403 10158
rect 1167 10097 1293 10103
rect 2867 10097 2893 10103
rect 1087 10077 1233 10083
rect 6987 10077 7053 10083
rect 8947 10077 9093 10083
rect 2547 10063 2560 10067
rect 2547 10053 2563 10063
rect 4787 10057 4853 10063
rect 5547 10057 5613 10063
rect 7827 10057 7933 10063
rect 2557 10027 2563 10053
rect 2547 10017 2563 10027
rect 2547 10013 2560 10017
rect 1127 9997 1193 10003
rect 2267 9997 2453 10003
rect 2747 9997 2793 10003
rect 2807 9997 2873 10003
rect 3147 9997 3193 10003
rect 4787 9997 4933 10003
rect 6907 9997 7073 10003
rect 8327 9997 8433 10003
rect 10047 9997 10073 10003
rect 1207 9977 1293 9983
rect -63 9882 30 9898
rect -63 9378 -3 9882
rect 397 9863 403 9883
rect 347 9857 403 9863
rect 5727 9857 5773 9863
rect 367 9777 453 9783
rect 1327 9777 1373 9783
rect 3407 9777 3493 9783
rect 4627 9777 4773 9783
rect 2440 9763 2453 9767
rect 2437 9753 2453 9763
rect 5707 9757 5813 9763
rect 7587 9757 7693 9763
rect 2437 9727 2443 9753
rect 2327 9717 2373 9723
rect 2437 9717 2453 9727
rect 2440 9713 2453 9717
rect 3707 9717 3753 9723
rect 6267 9717 6293 9723
rect 6847 9717 6953 9723
rect 7087 9717 7173 9723
rect 7347 9717 7453 9723
rect 7787 9697 7833 9703
rect 11343 9638 11403 10142
rect 11310 9622 11403 9638
rect 1107 9577 1173 9583
rect 1427 9557 1473 9563
rect 3307 9557 3413 9563
rect 4467 9557 4513 9563
rect 10407 9557 10593 9563
rect 2907 9537 2993 9543
rect 9327 9537 9433 9543
rect 5047 9517 5113 9523
rect 7467 9517 7513 9523
rect 2267 9497 2313 9503
rect 5033 9503 5047 9513
rect 5007 9500 5047 9503
rect 5007 9497 5043 9500
rect 5927 9497 6033 9503
rect 227 9477 413 9483
rect 1327 9477 1493 9483
rect 3887 9477 3953 9483
rect 4007 9477 4113 9483
rect 4467 9477 4613 9483
rect 7167 9477 7233 9483
rect 9487 9477 9533 9483
rect 9767 9477 9933 9483
rect 9987 9477 10093 9483
rect 10227 9477 10353 9483
rect 2967 9457 2993 9463
rect 9147 9457 9213 9463
rect 4767 9397 4873 9403
rect -63 9362 30 9378
rect -63 9315 -3 9362
rect 3747 9337 3773 9343
rect 3787 9337 3873 9343
rect -63 9307 -55 9315
rect -54 9307 -3 9315
rect -63 8858 -3 9307
rect 4947 9297 5013 9303
rect 3227 9277 3293 9283
rect 1287 9257 1313 9263
rect 2867 9257 2913 9263
rect 4067 9257 4133 9263
rect 4247 9257 4373 9263
rect 5427 9257 5473 9263
rect 2847 9237 2893 9243
rect 3007 9243 3020 9247
rect 4100 9243 4113 9247
rect 3007 9233 3023 9243
rect 3017 9207 3023 9233
rect 3007 9197 3023 9207
rect 4097 9233 4113 9243
rect 5187 9237 5273 9243
rect 4097 9207 4103 9233
rect 4097 9197 4113 9207
rect 3007 9193 3020 9197
rect 4100 9193 4113 9197
rect 5707 9197 5753 9203
rect 2387 9177 2453 9183
rect 2587 9177 2653 9183
rect 3527 9177 3673 9183
rect 5127 9177 5213 9183
rect 5267 9177 5313 9183
rect 5667 9177 5733 9183
rect 8507 9177 8613 9183
rect 6107 9157 6213 9163
rect 5167 9137 5273 9143
rect 11343 9118 11403 9622
rect 11310 9102 11403 9118
rect 5007 9057 5073 9063
rect 1427 9037 1513 9043
rect 4687 9037 4853 9043
rect 120 9023 133 9027
rect 117 9013 133 9023
rect 4987 9017 5013 9023
rect 117 8987 123 9013
rect 5287 8997 5323 9003
rect 5317 8987 5323 8997
rect 117 8977 133 8987
rect 120 8973 133 8977
rect 5317 8977 5333 8987
rect 5320 8973 5333 8977
rect 2687 8957 2813 8963
rect 4947 8957 5113 8963
rect 5207 8957 5253 8963
rect 5667 8957 5753 8963
rect 5867 8957 6073 8963
rect 7507 8957 7633 8963
rect 3587 8917 3673 8923
rect 4747 8877 4833 8883
rect -63 8842 30 8858
rect -63 8338 -3 8842
rect 2067 8817 2093 8823
rect 8497 8823 8503 8843
rect 8427 8817 8503 8823
rect 8687 8817 8713 8823
rect 4927 8797 5013 8803
rect 4887 8777 4913 8783
rect 2947 8737 2993 8743
rect 4027 8737 4073 8743
rect 4247 8737 4313 8743
rect 4967 8737 5033 8743
rect 5387 8737 5473 8743
rect 5487 8737 5513 8743
rect 5787 8737 5953 8743
rect 6107 8737 6193 8743
rect 3947 8717 4033 8723
rect 4167 8723 4180 8727
rect 4520 8723 4533 8727
rect 4167 8713 4183 8723
rect 4177 8687 4183 8713
rect 4517 8713 4533 8723
rect 4717 8717 4773 8723
rect 4167 8677 4183 8687
rect 4167 8673 4180 8677
rect 4517 8683 4523 8713
rect 4717 8686 4723 8717
rect 4407 8677 4523 8683
rect 4887 8677 4953 8683
rect 5127 8677 5193 8683
rect 5347 8677 5473 8683
rect 2787 8657 2813 8663
rect 2827 8657 2873 8663
rect 4647 8657 4813 8663
rect 6107 8657 6133 8663
rect 2727 8637 2833 8643
rect 5787 8637 5813 8643
rect 6307 8637 6333 8643
rect 3207 8617 3313 8623
rect 5667 8617 5693 8623
rect 11343 8598 11403 9102
rect 11310 8582 11403 8598
rect 4067 8557 4133 8563
rect 6307 8557 6413 8563
rect 4247 8537 4333 8543
rect 6347 8537 6393 8543
rect 227 8517 293 8523
rect 3347 8517 3473 8523
rect 4027 8517 4173 8523
rect 4487 8517 4513 8523
rect 4987 8517 5153 8523
rect 6287 8517 6353 8523
rect 3587 8497 3693 8503
rect 9367 8497 9473 8503
rect 3127 8457 3213 8463
rect 3847 8457 3933 8463
rect 4147 8457 4193 8463
rect 4747 8457 4853 8463
rect 5667 8457 5753 8463
rect 6107 8457 6133 8463
rect 10287 8457 10373 8463
rect 1347 8437 1393 8443
rect 4967 8437 4993 8443
rect 5087 8437 5133 8443
rect 5627 8437 5833 8443
rect 6107 8437 6153 8443
rect 7527 8437 7613 8443
rect 8287 8437 8313 8443
rect 10007 8437 10113 8443
rect 10307 8437 10433 8443
rect 5027 8357 5093 8363
rect -63 8322 30 8338
rect -63 7818 -3 8322
rect 397 8307 403 8323
rect 387 8297 403 8307
rect 3817 8300 3913 8303
rect 3813 8297 3913 8300
rect 387 8293 400 8297
rect 3813 8287 3827 8297
rect 10607 8277 10693 8283
rect 3107 8243 3120 8247
rect 3107 8240 3123 8243
rect 3107 8233 3127 8240
rect 3113 8227 3127 8233
rect 1347 8217 1473 8223
rect 1727 8217 1813 8223
rect 3567 8217 3673 8223
rect 4007 8217 4213 8223
rect 5107 8217 5193 8223
rect 6227 8217 6393 8223
rect 7127 8217 7233 8223
rect 10587 8217 10713 8223
rect 3827 8197 3933 8203
rect 6347 8197 6373 8203
rect 4107 8157 4193 8163
rect 7087 8157 7193 8163
rect 8247 8157 8353 8163
rect 8447 8157 8493 8163
rect 2427 8137 2573 8143
rect 5787 8137 5933 8143
rect 5987 8137 6133 8143
rect 6267 8137 6393 8143
rect 8567 8137 8593 8143
rect 10087 8137 10133 8143
rect 10187 8137 10273 8143
rect 1127 8117 1253 8123
rect 6447 8117 6593 8123
rect 7367 8117 7473 8123
rect 11343 8078 11403 8582
rect 11310 8062 11403 8078
rect 2907 8040 2983 8043
rect 2907 8037 2987 8040
rect 2973 8027 2987 8037
rect 5467 8037 5553 8043
rect 5507 8017 5613 8023
rect 2387 7997 2533 8003
rect 2687 7997 2733 8003
rect 3747 7997 3933 8003
rect 4707 7997 4793 8003
rect 5207 7997 5293 8003
rect 5907 7997 6033 8003
rect 9907 7997 9953 8003
rect 5007 7977 5073 7983
rect 6447 7977 6493 7983
rect 4093 7943 4107 7953
rect 4047 7940 4107 7943
rect 4047 7937 4103 7940
rect 1847 7917 1913 7923
rect 2307 7917 2533 7923
rect 3067 7917 3153 7923
rect 3767 7917 3813 7923
rect 3827 7917 3973 7923
rect 4167 7917 4193 7923
rect 4807 7917 4913 7923
rect 5307 7917 5393 7923
rect 4027 7897 4173 7903
rect 4527 7897 4633 7903
rect 8847 7877 8913 7883
rect 2687 7837 2753 7843
rect 3207 7837 3233 7843
rect 3327 7837 3373 7843
rect 4047 7837 4153 7843
rect 5007 7837 5033 7843
rect -63 7802 30 7818
rect -63 7298 -3 7802
rect 2777 7783 2783 7803
rect 11317 7787 11323 7803
rect 2707 7777 2783 7783
rect 11307 7777 11323 7787
rect 11307 7773 11320 7777
rect 4327 7737 4373 7743
rect 10087 7717 10213 7723
rect 1007 7697 1073 7703
rect 2887 7697 3073 7703
rect 3187 7697 3313 7703
rect 4147 7697 4233 7703
rect 4367 7697 4453 7703
rect 4807 7697 4933 7703
rect 7207 7697 7253 7703
rect 7267 7697 7293 7703
rect 8747 7697 8853 7703
rect 8867 7697 8913 7703
rect 9667 7697 9813 7703
rect 10127 7697 10253 7703
rect 10367 7697 10453 7703
rect 10587 7697 10773 7703
rect 2667 7683 2680 7687
rect 2667 7673 2683 7683
rect 4547 7677 4613 7683
rect 5427 7683 5440 7687
rect 5427 7673 5443 7683
rect 10607 7683 10620 7687
rect 10700 7683 10713 7687
rect 10607 7680 10623 7683
rect 10607 7673 10627 7680
rect 1827 7637 1853 7643
rect 2677 7643 2683 7673
rect 2677 7637 2793 7643
rect 5047 7637 5113 7643
rect 5437 7643 5443 7673
rect 10613 7666 10627 7673
rect 10697 7673 10713 7683
rect 10697 7647 10703 7673
rect 5417 7640 5443 7643
rect 5413 7637 5443 7640
rect 5413 7627 5427 7637
rect 7287 7637 7353 7643
rect 7647 7637 7733 7643
rect 10697 7637 10713 7647
rect 10700 7633 10713 7637
rect 2427 7617 2493 7623
rect 2507 7617 2573 7623
rect 3167 7617 3273 7623
rect 4807 7617 4873 7623
rect 7287 7617 7373 7623
rect 7627 7617 7693 7623
rect 7707 7617 7733 7623
rect 9687 7617 9773 7623
rect 9787 7617 9833 7623
rect 10627 7617 10733 7623
rect 5447 7597 5573 7603
rect 7027 7577 7093 7583
rect 11343 7558 11403 8062
rect 11310 7542 11403 7558
rect 447 7497 553 7503
rect 9627 7500 9723 7503
rect 9627 7497 9727 7500
rect 9713 7487 9727 7497
rect 1527 7477 1633 7483
rect 2627 7477 2793 7483
rect 4987 7477 5023 7483
rect 1640 7463 1653 7467
rect 1637 7460 1653 7463
rect 1633 7453 1653 7460
rect 5017 7463 5023 7477
rect 6087 7477 6233 7483
rect 7547 7477 7633 7483
rect 10927 7477 11113 7483
rect 5017 7457 5043 7463
rect 1633 7446 1647 7453
rect 5037 7447 5043 7457
rect 5467 7463 5480 7467
rect 5467 7453 5483 7463
rect 5037 7446 5060 7447
rect 5037 7437 5053 7446
rect 5040 7433 5053 7437
rect 5477 7427 5483 7453
rect 5467 7417 5483 7427
rect 5467 7413 5480 7417
rect 8447 7417 8533 7423
rect 2027 7397 2093 7403
rect 4967 7397 5173 7403
rect 5727 7397 5833 7403
rect 6847 7397 6973 7403
rect 8987 7397 9033 7403
rect 9187 7397 9253 7403
rect 10747 7397 10853 7403
rect 1987 7377 2073 7383
rect 5667 7377 5733 7383
rect 8907 7377 8953 7383
rect 10507 7377 10633 7383
rect 5307 7357 5353 7363
rect -63 7282 30 7298
rect -63 6778 -3 7282
rect 1437 7263 1443 7283
rect 1387 7257 1443 7263
rect 2047 7257 2133 7263
rect 9807 7257 9893 7263
rect 4187 7177 4293 7183
rect 9947 7177 9993 7183
rect 707 7157 753 7163
rect 767 7157 813 7163
rect 3927 7157 4053 7163
rect 5180 7163 5193 7167
rect 5177 7153 5193 7163
rect 5177 7127 5183 7153
rect 7567 7137 7593 7143
rect 2727 7117 2853 7123
rect 5177 7117 5193 7127
rect 5180 7113 5193 7117
rect 5580 7123 5593 7127
rect 5577 7113 5593 7123
rect 5747 7117 5793 7123
rect 6507 7117 6593 7123
rect 6687 7117 6793 7123
rect 7827 7117 7873 7123
rect 3467 7097 3513 7103
rect 5577 7083 5583 7113
rect 5607 7097 5693 7103
rect 6667 7097 6753 7103
rect 9647 7097 9733 7103
rect 5577 7077 5613 7083
rect 8887 7077 8913 7083
rect 3207 7057 3313 7063
rect 11343 7038 11403 7542
rect 11310 7022 11403 7038
rect 5227 6997 5313 7003
rect 5467 6997 5593 7003
rect 5247 6977 5293 6983
rect 6107 6977 6253 6983
rect 2507 6957 2633 6963
rect 4107 6957 4173 6963
rect 4367 6957 4393 6963
rect 4607 6957 4733 6963
rect 4987 6957 5173 6963
rect 5847 6957 5933 6963
rect 7127 6957 7173 6963
rect 8867 6957 9053 6963
rect 4347 6937 4413 6943
rect 7627 6937 7673 6943
rect 9487 6937 9513 6943
rect 6347 6897 6433 6903
rect 7367 6897 7413 6903
rect 7547 6897 7613 6903
rect 3807 6877 3843 6883
rect 2533 6863 2547 6873
rect 3837 6867 3843 6877
rect 3887 6877 3913 6883
rect 6327 6877 6433 6883
rect 7387 6877 7453 6883
rect 8927 6877 9033 6883
rect 9607 6877 9653 6883
rect 2533 6860 2573 6863
rect 2537 6857 2573 6860
rect 3727 6857 3833 6863
rect 3887 6857 3993 6863
rect 6367 6857 6453 6863
rect 2667 6837 2693 6843
rect 4253 6843 4267 6853
rect 4167 6840 4267 6843
rect 4167 6837 4263 6840
rect -63 6762 30 6778
rect -63 6258 -3 6762
rect 11147 6737 11193 6743
rect 3073 6703 3087 6713
rect 2927 6700 3087 6703
rect 2927 6697 3083 6700
rect 5487 6697 5533 6703
rect 2287 6657 2393 6663
rect 9867 6657 9913 6663
rect 3207 6637 3293 6643
rect 10687 6617 10713 6623
rect 5447 6597 5473 6603
rect 7987 6597 8113 6603
rect 8647 6597 8753 6603
rect 9107 6597 9153 6603
rect 2047 6577 2113 6583
rect 3847 6577 3933 6583
rect 5467 6577 5553 6583
rect 6447 6577 6473 6583
rect 6667 6577 6693 6583
rect 8847 6577 8893 6583
rect 8907 6577 8933 6583
rect 9367 6577 9453 6583
rect 11007 6577 11033 6583
rect 3867 6557 3933 6563
rect 8007 6557 8093 6563
rect 3167 6537 3273 6543
rect 11343 6518 11403 7022
rect 11310 6502 11403 6518
rect 2547 6457 2573 6463
rect 2667 6437 2793 6443
rect 4087 6437 4213 6443
rect 4347 6437 4513 6443
rect 8307 6437 8393 6443
rect 2967 6417 3013 6423
rect 3907 6417 3973 6423
rect 8107 6423 8120 6427
rect 8813 6423 8827 6433
rect 8107 6413 8123 6423
rect 8813 6420 8853 6423
rect 8817 6417 8853 6420
rect 9727 6417 9813 6423
rect 9827 6417 9853 6423
rect 2967 6377 3013 6383
rect 447 6357 533 6363
rect 2567 6357 2613 6363
rect 2727 6357 2773 6363
rect 3647 6357 3693 6363
rect 3787 6357 3813 6363
rect 4587 6357 4713 6363
rect 5147 6357 5212 6363
rect 5247 6357 5373 6363
rect 6207 6357 6273 6363
rect 6427 6357 6633 6363
rect 6687 6357 6773 6363
rect 6787 6357 6813 6363
rect 8117 6366 8123 6413
rect 8307 6357 8513 6363
rect 9707 6357 9913 6363
rect 2560 6346 2580 6347
rect 2427 6337 2553 6343
rect 2567 6343 2580 6346
rect 2567 6337 2583 6343
rect 2567 6333 2580 6337
rect 6327 6337 6373 6343
rect -63 6242 30 6258
rect -63 5738 -3 6242
rect 5937 6223 5943 6243
rect 5937 6217 5973 6223
rect 6947 6217 6993 6223
rect 8537 6223 8543 6243
rect 8537 6217 8593 6223
rect 10377 6223 10383 6243
rect 10377 6217 10433 6223
rect 7667 6177 7733 6183
rect 1407 6137 1573 6143
rect 3687 6137 3893 6143
rect 5907 6137 6013 6143
rect 6867 6137 6893 6143
rect 8307 6137 8453 6143
rect 8807 6137 8953 6143
rect 10247 6137 10313 6143
rect 10427 6137 10533 6143
rect 1187 6117 1213 6123
rect 5300 6123 5313 6127
rect 5297 6113 5313 6123
rect 5927 6117 5993 6123
rect 6527 6117 6553 6123
rect 7007 6117 7073 6123
rect 9727 6123 9740 6127
rect 9727 6113 9743 6123
rect 10927 6117 10973 6123
rect 2693 6087 2707 6093
rect 5297 6087 5303 6113
rect 9737 6087 9743 6113
rect 2693 6083 2713 6087
rect 2567 6077 2713 6083
rect 2700 6073 2713 6077
rect 3507 6077 3533 6083
rect 5297 6077 5313 6087
rect 5300 6073 5313 6077
rect 6527 6077 6553 6083
rect 9587 6080 9623 6083
rect 9587 6077 9627 6080
rect 9613 6067 9627 6077
rect 9727 6077 9743 6087
rect 9727 6073 9740 6077
rect 9947 6077 10053 6083
rect 1687 6057 1773 6063
rect 3767 6057 3893 6063
rect 3947 6057 4073 6063
rect 6547 6057 6673 6063
rect 10747 6057 10793 6063
rect 8127 6017 8253 6023
rect 11107 6017 11193 6023
rect 11343 5998 11403 6502
rect 11310 5982 11403 5998
rect 10887 5937 10973 5943
rect 5027 5917 5053 5923
rect 7647 5917 7713 5923
rect 1447 5897 1513 5903
rect 2607 5897 2653 5903
rect 4620 5903 4633 5907
rect 4617 5893 4633 5903
rect 6047 5897 6093 5903
rect 7827 5903 7840 5907
rect 7827 5893 7843 5903
rect 7887 5897 7953 5903
rect 11107 5903 11120 5907
rect 11107 5893 11123 5903
rect 1887 5840 2083 5843
rect 1887 5837 2087 5840
rect 2073 5827 2087 5837
rect 3127 5837 3153 5843
rect 3867 5837 3973 5843
rect 4617 5843 4623 5893
rect 7837 5867 7843 5893
rect 11117 5867 11123 5893
rect 6747 5857 6813 5863
rect 7827 5857 7843 5867
rect 7827 5853 7840 5857
rect 11107 5857 11123 5867
rect 11107 5853 11120 5857
rect 4617 5837 4653 5843
rect 6247 5837 6333 5843
rect 10867 5837 10973 5843
rect 11087 5837 11233 5843
rect 6487 5757 6613 5763
rect -63 5722 30 5738
rect -63 5218 -3 5722
rect 727 5617 873 5623
rect 1107 5617 1153 5623
rect 1807 5617 1873 5623
rect 2067 5617 2153 5623
rect 2607 5617 2773 5623
rect 3287 5617 3313 5623
rect 4147 5617 4193 5623
rect 5067 5617 5103 5623
rect 4487 5597 4513 5603
rect 5097 5603 5103 5617
rect 5127 5617 5173 5623
rect 5827 5617 5893 5623
rect 6027 5617 6113 5623
rect 6927 5617 6953 5623
rect 5097 5600 5123 5603
rect 5097 5597 5127 5600
rect 5113 5587 5127 5597
rect 11277 5567 11283 5633
rect 11297 5627 11303 5653
rect 4147 5557 4173 5563
rect 7207 5557 7313 5563
rect 11277 5566 11300 5567
rect 11277 5557 11293 5566
rect 11280 5553 11293 5557
rect 1147 5537 1293 5543
rect 1547 5537 1693 5543
rect 9427 5537 9593 5543
rect 1947 5497 1993 5503
rect 11343 5478 11403 5982
rect 11310 5462 11403 5478
rect 2667 5437 2793 5443
rect 2867 5437 2993 5443
rect 5807 5437 5913 5443
rect 7847 5417 7893 5423
rect 1507 5377 1593 5383
rect 2313 5383 2327 5393
rect 2297 5380 2327 5383
rect 2413 5383 2427 5393
rect 6267 5397 6393 5403
rect 2413 5380 2513 5383
rect 2297 5377 2323 5380
rect 2417 5377 2513 5380
rect 2297 5343 2303 5377
rect 6227 5377 6313 5383
rect 8307 5383 8320 5387
rect 8307 5373 8323 5383
rect 10187 5377 10283 5383
rect 8317 5347 8323 5373
rect 2297 5337 2323 5343
rect 1127 5317 1373 5323
rect 1547 5317 1653 5323
rect 2317 5323 2323 5337
rect 2767 5337 2793 5343
rect 8147 5337 8213 5343
rect 8307 5337 8323 5347
rect 10277 5347 10283 5377
rect 10277 5337 10293 5347
rect 8307 5333 8320 5337
rect 10280 5333 10293 5337
rect 2127 5317 2303 5323
rect 2317 5317 2373 5323
rect 2247 5297 2273 5303
rect 2297 5303 2303 5317
rect 5787 5317 5813 5323
rect 6067 5317 6153 5323
rect 6207 5317 6413 5323
rect 6767 5317 6833 5323
rect 7867 5317 7993 5323
rect 8287 5317 8393 5323
rect 9207 5317 9233 5323
rect 2297 5297 2333 5303
rect 3047 5297 3193 5303
rect 4227 5297 4253 5303
rect 2207 5277 2293 5283
rect 6813 5263 6827 5273
rect 6767 5260 6827 5263
rect 6767 5257 6823 5260
rect 2687 5237 2773 5243
rect 6707 5237 6793 5243
rect 6927 5237 7013 5243
rect -63 5202 30 5218
rect -63 4698 -3 5202
rect 2127 5177 2253 5183
rect 2587 5177 2673 5183
rect 2147 5157 2233 5163
rect 10727 5157 10773 5163
rect 6533 5123 6547 5133
rect 6533 5120 6693 5123
rect 6537 5117 6693 5120
rect 9927 5117 9953 5123
rect 527 5097 733 5103
rect 1647 5097 1733 5103
rect 1987 5097 2053 5103
rect 2567 5097 2713 5103
rect 2987 5097 3053 5103
rect 3067 5097 3193 5103
rect 5087 5097 5153 5103
rect 6307 5097 6413 5103
rect 6587 5097 6693 5103
rect 8827 5097 8913 5103
rect 10907 5097 11013 5103
rect 11147 5097 11233 5103
rect 2460 5083 2473 5087
rect 2457 5073 2473 5083
rect 2587 5077 2673 5083
rect 6547 5077 6653 5083
rect 2457 5027 2463 5073
rect 2787 5037 2813 5043
rect 4540 5043 4553 5047
rect 4537 5040 4553 5043
rect 4533 5033 4553 5040
rect 5047 5037 5113 5043
rect 5667 5037 5813 5043
rect 8647 5037 8733 5043
rect 8867 5040 8983 5043
rect 8867 5037 8987 5040
rect 4533 5027 4547 5033
rect 8973 5027 8987 5037
rect 1907 5017 2053 5023
rect 2847 5017 2933 5023
rect 4587 5017 4653 5023
rect 4967 5017 5033 5023
rect 10827 5017 10973 5023
rect 2333 4983 2347 4993
rect 2333 4980 2393 4983
rect 2337 4977 2393 4980
rect 4127 4977 4153 4983
rect 6113 4983 6127 4993
rect 6113 4980 6233 4983
rect 6117 4977 6233 4980
rect 11343 4958 11403 5462
rect 11310 4942 11403 4958
rect 2687 4917 2773 4923
rect 7247 4917 7313 4923
rect 5367 4897 5473 4903
rect 1907 4877 1993 4883
rect 2187 4877 2273 4883
rect 6227 4877 6313 4883
rect 6487 4877 6613 4883
rect 7237 4877 7333 4883
rect 2187 4857 2293 4863
rect 4887 4857 4993 4863
rect 6087 4857 6173 4863
rect 7237 4847 7243 4877
rect 8147 4857 8263 4863
rect 8257 4827 8263 4857
rect 8887 4857 8913 4863
rect 8257 4817 8273 4827
rect 8260 4813 8273 4817
rect 2447 4797 2573 4803
rect 2947 4797 2973 4803
rect 6227 4797 6273 4803
rect 11127 4797 11313 4803
rect 1947 4777 2073 4783
rect 3327 4777 3393 4783
rect 11147 4777 11173 4783
rect 1687 4757 1773 4763
rect -63 4682 30 4698
rect -63 4178 -3 4682
rect 2087 4657 2213 4663
rect 6897 4663 6903 4683
rect 6847 4657 6903 4663
rect 7287 4657 7313 4663
rect 1887 4617 1953 4623
rect 3067 4617 3113 4623
rect 6767 4617 6833 4623
rect 2067 4597 2273 4603
rect 9607 4597 9653 4603
rect 667 4577 753 4583
rect 1607 4577 1673 4583
rect 1787 4577 1853 4583
rect 1947 4577 2013 4583
rect 2967 4577 3113 4583
rect 4867 4577 4893 4583
rect 6087 4577 6193 4583
rect 6567 4577 6613 4583
rect 5867 4557 5993 4563
rect 9327 4557 9393 4563
rect 11247 4557 11293 4563
rect 7267 4537 7313 4543
rect 3627 4517 3733 4523
rect 5707 4517 5753 4523
rect 2967 4477 3053 4483
rect 6627 4457 6713 4463
rect 11343 4438 11403 4942
rect 11310 4422 11403 4438
rect 3787 4397 3893 4403
rect 3867 4357 3913 4363
rect 8407 4357 8473 4363
rect 2940 4343 2953 4347
rect 2937 4333 2953 4343
rect 3767 4337 3873 4343
rect 4907 4337 5013 4343
rect 2937 4327 2943 4333
rect 2920 4326 2943 4327
rect 2927 4317 2943 4326
rect 2927 4313 2940 4317
rect 2407 4297 2523 4303
rect 2517 4283 2523 4297
rect 3547 4297 3633 4303
rect 7427 4297 7453 4303
rect 2517 4277 2553 4283
rect 3047 4277 3233 4283
rect 3527 4277 3553 4283
rect 4427 4277 4573 4283
rect 4787 4277 4833 4283
rect 4987 4277 5073 4283
rect 6147 4277 6193 4283
rect 6627 4277 6833 4283
rect 6887 4277 7053 4283
rect 7167 4277 7233 4283
rect 2407 4257 2513 4263
rect 6087 4257 6173 4263
rect 2227 4217 2253 4223
rect 3193 4203 3207 4213
rect 3107 4200 3207 4203
rect 3107 4197 3203 4200
rect 4487 4197 4553 4203
rect 7207 4197 7293 4203
rect -63 4162 30 4178
rect -63 3658 -3 4162
rect 4567 4137 4673 4143
rect 11317 4143 11323 4163
rect 11247 4137 11323 4143
rect 1687 4097 1713 4103
rect 3107 4077 3133 4083
rect 1087 4057 1333 4063
rect 2687 4057 2753 4063
rect 3247 4057 3393 4063
rect 3707 4057 3833 4063
rect 4227 4057 4293 4063
rect 5727 4057 5893 4063
rect 6927 4057 7093 4063
rect 8087 4057 8213 4063
rect 3027 4037 3133 4043
rect 3360 4043 3373 4047
rect 3357 4033 3373 4043
rect 3357 4007 3363 4033
rect 7687 4037 7713 4043
rect 3477 4017 3573 4023
rect 3477 4007 3483 4017
rect 2807 4000 2943 4003
rect 2807 3997 2947 4000
rect 3357 3997 3373 4007
rect 2933 3987 2947 3997
rect 3360 3993 3373 3997
rect 3467 3997 3483 4007
rect 3467 3993 3480 3997
rect 4347 3997 4453 4003
rect 6947 3997 7033 4003
rect 8887 3997 8913 4003
rect 9007 3997 9053 4003
rect 1247 3977 1273 3983
rect 1647 3977 1713 3983
rect 4907 3977 4953 3983
rect 9867 3977 9953 3983
rect 3887 3957 4033 3963
rect 6653 3943 6667 3953
rect 6653 3940 6793 3943
rect 6657 3937 6793 3940
rect 11343 3918 11403 4422
rect 11310 3902 11403 3918
rect 2787 3877 2873 3883
rect 5787 3877 5853 3883
rect 1227 3860 1323 3863
rect 1227 3857 1327 3860
rect 1313 3847 1327 3857
rect 2747 3857 2853 3863
rect 3167 3857 3273 3863
rect 3893 3863 3907 3873
rect 3893 3860 4013 3863
rect 3897 3857 4013 3860
rect 2587 3837 2693 3843
rect 3427 3837 3533 3843
rect 4107 3837 4133 3843
rect 7637 3837 7693 3843
rect 567 3817 633 3823
rect 3447 3817 3553 3823
rect 3707 3817 3793 3823
rect 7440 3823 7453 3827
rect 7437 3813 7453 3823
rect 7437 3787 7443 3813
rect 2307 3777 2373 3783
rect 2537 3777 2573 3783
rect 2537 3767 2543 3777
rect 2767 3777 2853 3783
rect 3187 3777 3253 3783
rect 7437 3777 7453 3787
rect 7440 3773 7453 3777
rect 1227 3757 1293 3763
rect 2187 3757 2233 3763
rect 2347 3757 2373 3763
rect 2527 3757 2543 3767
rect 2527 3753 2540 3757
rect 2567 3757 2693 3763
rect 4107 3757 4213 3763
rect 7087 3757 7153 3763
rect 7167 3757 7253 3763
rect 7637 3763 7643 3837
rect 8427 3837 8573 3843
rect 10467 3837 10573 3843
rect 7660 3823 7673 3827
rect 7657 3813 7673 3823
rect 7657 3787 7663 3813
rect 7657 3777 7673 3787
rect 7660 3773 7673 3777
rect 9207 3777 9313 3783
rect 9327 3777 9353 3783
rect 10907 3777 11013 3783
rect 7637 3757 7693 3763
rect 9107 3757 9293 3763
rect 10887 3757 10993 3763
rect 11007 3757 11073 3763
rect 7147 3737 7193 3743
rect 3027 3717 3053 3723
rect 2967 3677 2993 3683
rect -63 3642 30 3658
rect -63 3138 -3 3642
rect 2947 3617 3013 3623
rect 4527 3617 4573 3623
rect 1887 3577 1913 3583
rect 3347 3577 3473 3583
rect 2267 3557 2453 3563
rect 4907 3557 5033 3563
rect 9927 3557 10033 3563
rect 1907 3537 1973 3543
rect 2507 3537 2633 3543
rect 3087 3537 3113 3543
rect 3547 3537 3673 3543
rect 3807 3537 3913 3543
rect 3967 3537 4093 3543
rect 4787 3537 4833 3543
rect 7707 3537 7753 3543
rect 1407 3517 1473 3523
rect 1487 3517 1513 3523
rect 3460 3523 3473 3527
rect 3457 3513 3473 3523
rect 5587 3517 5653 3523
rect 9093 3523 9107 3533
rect 8987 3520 9107 3523
rect 8987 3517 9103 3520
rect 9647 3517 9773 3523
rect 3457 3487 3463 3513
rect 1167 3477 1293 3483
rect 2987 3477 3013 3483
rect 3347 3477 3373 3483
rect 3457 3477 3473 3487
rect 3460 3473 3473 3477
rect 4347 3477 4393 3483
rect 4687 3477 4753 3483
rect 1067 3457 1093 3463
rect 1227 3457 1293 3463
rect 3547 3457 3593 3463
rect 1827 3437 1933 3443
rect 2867 3437 3033 3443
rect 3787 3437 3813 3443
rect 8987 3437 9113 3443
rect 10187 3437 10233 3443
rect 3447 3417 3473 3423
rect 9647 3417 9773 3423
rect 11343 3398 11403 3902
rect 11310 3382 11403 3398
rect 1827 3357 1913 3363
rect 2727 3357 2773 3363
rect 3027 3357 3093 3363
rect 4407 3357 4533 3363
rect 10687 3357 10713 3363
rect 4147 3337 4173 3343
rect 1047 3317 1213 3323
rect 1587 3317 1673 3323
rect 3667 3317 3733 3323
rect 4607 3317 4733 3323
rect 6687 3317 6833 3323
rect 9227 3317 9313 3323
rect 1047 3297 1093 3303
rect 1607 3297 1653 3303
rect 9687 3303 9700 3307
rect 10020 3303 10033 3307
rect 9687 3293 9703 3303
rect 9697 3267 9703 3293
rect 1927 3257 1953 3263
rect 2987 3257 3053 3263
rect 7587 3257 7673 3263
rect 9687 3257 9703 3267
rect 10017 3293 10033 3303
rect 11107 3297 11153 3303
rect 10017 3263 10023 3293
rect 11307 3283 11320 3287
rect 11307 3273 11323 3283
rect 10017 3257 10043 3263
rect 9687 3253 9700 3257
rect 10037 3247 10043 3257
rect 1927 3237 1973 3243
rect 2607 3237 2653 3243
rect 2767 3237 2893 3243
rect 3107 3237 3153 3243
rect 3687 3237 3733 3243
rect 3967 3237 4093 3243
rect 4847 3237 4933 3243
rect 8327 3237 8413 3243
rect 9067 3237 9113 3243
rect 9167 3237 9293 3243
rect 9407 3237 9553 3243
rect 9787 3237 9813 3243
rect 9987 3237 10013 3243
rect 10037 3237 10053 3247
rect 10040 3233 10053 3237
rect 11247 3237 11293 3243
rect 1607 3217 1633 3223
rect 3833 3203 3847 3213
rect 3927 3217 4033 3223
rect 3727 3200 3847 3203
rect 3727 3197 3843 3200
rect 3573 3183 3587 3193
rect 3487 3180 3587 3183
rect 3487 3177 3583 3180
rect 2287 3157 2333 3163
rect 8967 3157 9073 3163
rect 9507 3157 9553 3163
rect -63 3122 30 3138
rect 11317 3137 11323 3273
rect -63 2618 -3 3122
rect 9967 3097 9993 3103
rect 4147 3077 4193 3083
rect 2307 3057 2373 3063
rect 2507 3057 2633 3063
rect 2767 3057 2893 3063
rect 1807 3037 1913 3043
rect 2017 3037 2153 3043
rect 1067 3017 1113 3023
rect 2017 3023 2023 3037
rect 2347 3037 2393 3043
rect 9767 3037 9793 3043
rect 1987 3017 2023 3023
rect 2157 3017 2193 3023
rect 1567 2997 1673 3003
rect 2157 3003 2163 3017
rect 2267 3017 2333 3023
rect 3687 3017 3713 3023
rect 4987 3017 5113 3023
rect 5427 3017 5453 3023
rect 6107 3017 6233 3023
rect 9787 3017 9833 3023
rect 2260 3006 2280 3007
rect 2137 2997 2163 3003
rect 2137 2967 2143 2997
rect 2267 3003 2280 3006
rect 2380 3003 2393 3007
rect 2267 2993 2283 3003
rect 2277 2983 2283 2993
rect 2377 2993 2393 3003
rect 3967 2997 4013 3003
rect 5247 2997 5353 3003
rect 2377 2983 2383 2993
rect 2277 2977 2383 2983
rect 927 2957 993 2963
rect 1087 2957 1213 2963
rect 1827 2957 1913 2963
rect 2137 2957 2153 2967
rect 2140 2953 2153 2957
rect 2307 2957 2353 2963
rect 2507 2957 2613 2963
rect 3227 2957 3273 2963
rect 5227 2957 5253 2963
rect 5927 2957 6033 2963
rect 447 2937 593 2943
rect 3407 2937 3493 2943
rect 3667 2937 3773 2943
rect 427 2917 493 2923
rect 1567 2897 1673 2903
rect 2987 2897 3113 2903
rect 3887 2897 4013 2903
rect 4167 2897 4253 2903
rect 4427 2897 4473 2903
rect 4807 2897 4893 2903
rect 5307 2897 5353 2903
rect 11343 2878 11403 3382
rect 11310 2862 11403 2878
rect 4747 2837 4793 2843
rect 4047 2797 4173 2803
rect 6407 2797 6453 2803
rect 8207 2797 8293 2803
rect 10487 2797 10533 2803
rect 4707 2777 4813 2783
rect 9747 2783 9760 2787
rect 9747 2780 9763 2783
rect 9747 2773 9767 2780
rect 9753 2766 9767 2773
rect 11097 2777 11213 2783
rect 11097 2747 11103 2777
rect 6847 2737 6893 2743
rect 11087 2737 11103 2747
rect 11087 2733 11100 2737
rect 127 2717 193 2723
rect 3627 2717 3693 2723
rect 3847 2717 3953 2723
rect 4747 2717 4833 2723
rect 9727 2717 9833 2723
rect 10007 2717 10093 2723
rect 4287 2637 4353 2643
rect -63 2602 30 2618
rect -63 2098 -3 2602
rect 4847 2577 4913 2583
rect 10577 2583 10583 2603
rect 10577 2577 10653 2583
rect 11007 2577 11073 2583
rect 2147 2557 2213 2563
rect 8327 2557 8433 2563
rect 747 2537 793 2543
rect 1627 2537 1673 2543
rect 2107 2537 2253 2543
rect 8327 2537 8473 2543
rect 2527 2517 2553 2523
rect 2567 2517 2673 2523
rect 4117 2517 4233 2523
rect 727 2497 813 2503
rect 1587 2497 1713 2503
rect 1967 2497 1993 2503
rect 4117 2503 4123 2517
rect 4087 2497 4123 2503
rect 4587 2497 4613 2503
rect 8747 2497 8793 2503
rect 8967 2497 9013 2503
rect 9647 2497 9753 2503
rect 4607 2477 4713 2483
rect 7507 2477 7553 2483
rect 8547 2477 8573 2483
rect 11047 2477 11133 2483
rect 1887 2437 1933 2443
rect 2987 2437 3093 2443
rect 8587 2437 8673 2443
rect 10647 2437 10693 2443
rect 1887 2417 2013 2423
rect 4787 2417 4893 2423
rect 4887 2397 4933 2403
rect 2107 2377 2213 2383
rect 5227 2377 5333 2383
rect 11343 2358 11403 2862
rect 11310 2342 11403 2358
rect 7947 2317 7993 2323
rect 1107 2297 1253 2303
rect 2547 2297 2613 2303
rect 5047 2297 5093 2303
rect 5787 2297 5853 2303
rect 7887 2297 7993 2303
rect 9567 2297 9613 2303
rect 10887 2297 10913 2303
rect 267 2277 393 2283
rect 447 2277 553 2283
rect 5287 2277 5333 2283
rect 6487 2277 6533 2283
rect 10207 2277 10293 2283
rect 10727 2277 10813 2283
rect 1827 2263 1840 2267
rect 1827 2253 1843 2263
rect 4587 2257 4693 2263
rect 6247 2257 6333 2263
rect 8007 2257 8033 2263
rect 9567 2257 9713 2263
rect 767 2197 793 2203
rect 867 2197 1013 2203
rect 1837 2203 1843 2253
rect 2047 2217 2113 2223
rect 8887 2217 8993 2223
rect 1807 2197 1843 2203
rect 2267 2197 2453 2203
rect 2947 2197 3033 2203
rect 3057 2183 3063 2213
rect 3947 2197 4013 2203
rect 5227 2197 5313 2203
rect 5467 2197 5513 2203
rect 5527 2197 5633 2203
rect 8847 2197 9033 2203
rect 9987 2197 10013 2203
rect 10447 2197 10513 2203
rect 10727 2197 10813 2203
rect 10867 2197 10973 2203
rect 2967 2177 3063 2183
rect 10007 2177 10033 2183
rect 1847 2157 1933 2163
rect 2747 2157 2853 2163
rect 967 2137 993 2143
rect 5247 2117 5293 2123
rect -63 2082 30 2098
rect -63 1578 -3 2082
rect 3147 2057 3273 2063
rect 6567 2037 6673 2043
rect 1547 2017 1693 2023
rect 11027 1997 11173 2003
rect 2567 1977 2633 1983
rect 3367 1977 3393 1983
rect 3507 1977 3573 1983
rect 1127 1957 1233 1963
rect 1393 1963 1407 1973
rect 7287 1977 7373 1983
rect 8807 1977 8853 1983
rect 9767 1977 9793 1983
rect 10307 1977 10333 1983
rect 1347 1960 1407 1963
rect 1347 1957 1403 1960
rect 3627 1957 3733 1963
rect 4087 1957 4193 1963
rect 4747 1957 4813 1963
rect 6147 1957 6233 1963
rect 9667 1957 9733 1963
rect 9980 1963 9993 1967
rect 9977 1953 9993 1963
rect 10567 1963 10580 1967
rect 10567 1953 10583 1963
rect 3147 1917 3253 1923
rect 8987 1917 9073 1923
rect 9667 1917 9713 1923
rect 9977 1923 9983 1953
rect 10577 1927 10583 1953
rect 9867 1917 9983 1923
rect 10567 1917 10583 1927
rect 10567 1913 10580 1917
rect 5647 1877 5753 1883
rect 5907 1857 5933 1863
rect 7447 1857 7573 1863
rect 11343 1838 11403 2342
rect 11310 1822 11403 1838
rect 3307 1757 3453 1763
rect 9197 1760 9333 1763
rect 9193 1757 9333 1760
rect 9193 1747 9207 1757
rect 9927 1757 10073 1763
rect 6967 1737 7073 1743
rect 10340 1746 10360 1747
rect 10347 1743 10360 1746
rect 10347 1733 10363 1743
rect 2027 1697 2093 1703
rect 9207 1697 9233 1703
rect 9527 1697 9573 1703
rect 1107 1677 1233 1683
rect 2067 1677 2153 1683
rect 2667 1677 2793 1683
rect 3087 1677 3193 1683
rect 5767 1677 5973 1683
rect 7027 1677 7093 1683
rect 10127 1677 10273 1683
rect 10357 1683 10363 1733
rect 10327 1677 10363 1683
rect 1067 1637 1213 1643
rect 1287 1637 1333 1643
rect 3807 1597 3913 1603
rect -63 1562 30 1578
rect -63 1058 -3 1562
rect 9127 1537 9233 1543
rect 8447 1517 8473 1523
rect 4933 1503 4947 1513
rect 4847 1500 4947 1503
rect 4847 1497 4943 1500
rect 8847 1497 8953 1503
rect 3787 1477 3933 1483
rect 3287 1457 3393 1463
rect 5047 1457 5093 1463
rect 5947 1457 5993 1463
rect 8047 1457 8073 1463
rect 9087 1457 9213 1463
rect 9707 1457 9833 1463
rect 10187 1457 10333 1463
rect 10847 1457 10953 1463
rect 8857 1400 8993 1403
rect 8853 1397 8993 1400
rect 8853 1387 8867 1397
rect 10667 1397 10733 1403
rect 1827 1377 1853 1383
rect 5067 1377 5093 1383
rect 10187 1377 10333 1383
rect 1307 1357 1453 1363
rect 7057 1360 7173 1363
rect 7053 1357 7173 1360
rect 7053 1347 7067 1357
rect 11343 1318 11403 1822
rect 11310 1302 11403 1318
rect 2007 1277 2133 1283
rect 10387 1277 10473 1283
rect 3647 1237 3793 1243
rect 3847 1237 3953 1243
rect 6167 1237 6273 1243
rect 8807 1237 8873 1243
rect 9027 1237 9113 1243
rect 4767 1217 4873 1223
rect 10147 1217 10213 1223
rect 3617 1180 3693 1183
rect 3613 1177 3693 1180
rect 3613 1167 3627 1177
rect 11087 1177 11133 1183
rect 2347 1157 2373 1163
rect 6147 1157 6233 1163
rect 8407 1157 8473 1163
rect 8627 1157 8713 1163
rect 11067 1157 11213 1163
rect 10107 1137 10253 1143
rect 5747 1117 5853 1123
rect 9247 1117 9373 1123
rect -63 1042 30 1058
rect -63 538 -3 1042
rect 3387 957 3533 963
rect 8907 957 9013 963
rect 1487 937 1573 943
rect 2687 937 2813 943
rect 3327 937 3413 943
rect 3427 937 3493 943
rect 4227 937 4313 943
rect 4607 937 4633 943
rect 7267 937 7313 943
rect 10987 937 11053 943
rect 4307 917 4413 923
rect 11007 877 11033 883
rect 11343 798 11403 1302
rect 11310 782 11403 798
rect 5547 717 5613 723
rect 6487 717 6613 723
rect 7867 717 7953 723
rect 9087 717 9213 723
rect 9407 717 9433 723
rect 9487 717 9653 723
rect 4993 703 5007 713
rect 4947 700 5007 703
rect 4947 697 5003 700
rect 8447 677 8493 683
rect 847 637 913 643
rect 4367 637 4413 643
rect 4867 637 4953 643
rect 4967 637 5013 643
rect 6227 637 6393 643
rect 7867 637 7933 643
rect 5787 617 5933 623
rect 10647 597 10733 603
rect 7947 557 8073 563
rect -63 522 30 538
rect -63 18 -3 522
rect 2207 417 2393 423
rect 2647 417 2753 423
rect 3447 417 3673 423
rect 3747 417 3913 423
rect 8467 417 8573 423
rect 10307 417 10353 423
rect 227 397 333 403
rect 10507 397 10533 403
rect 6207 357 6233 363
rect 467 337 573 343
rect 3247 337 3313 343
rect 4187 337 4213 343
rect 5527 337 5553 343
rect 10007 337 10073 343
rect 10207 297 10273 303
rect 11343 278 11403 782
rect 11310 262 11403 278
rect 8127 197 8293 203
rect 8347 137 8473 143
rect 9247 137 9333 143
rect 2727 117 2833 123
rect 9247 117 9333 123
rect 9707 117 9833 123
rect -63 2 30 18
rect 11343 2 11403 262
<< m2contact >>
rect 9073 11113 9087 11127
rect 9173 11113 9187 11127
rect 3373 11033 3387 11047
rect 3453 11033 3467 11047
rect 6733 11033 6747 11047
rect 6913 11033 6927 11047
rect 333 10933 347 10947
rect 1053 10913 1067 10927
rect 2613 10913 2627 10927
rect 4573 10913 4587 10927
rect 7353 10833 7367 10847
rect 7473 10833 7487 10847
rect 7073 10813 7087 10827
rect 7193 10813 7207 10827
rect 7453 10813 7467 10827
rect 7533 10813 7547 10827
rect 8253 10814 8267 10828
rect 8453 10813 8467 10827
rect 7353 10793 7367 10807
rect 7413 10793 7427 10807
rect 6213 10733 6227 10747
rect 6293 10733 6307 10747
rect 6353 10733 6367 10747
rect 6393 10733 6407 10747
rect 10793 10733 10807 10747
rect 10993 10733 11007 10747
rect 2453 10593 2467 10607
rect 2473 10593 2487 10607
rect 2593 10593 2607 10607
rect 8993 10593 9007 10607
rect 9033 10593 9047 10607
rect 5653 10573 5667 10587
rect 5753 10573 5767 10587
rect 9533 10533 9547 10547
rect 9573 10533 9587 10547
rect 2473 10513 2487 10527
rect 2693 10513 2707 10527
rect 3413 10513 3427 10527
rect 3553 10513 3567 10527
rect 4473 10513 4487 10527
rect 4593 10513 4607 10527
rect 4693 10513 4707 10527
rect 4873 10513 4887 10527
rect 6753 10513 6767 10527
rect 6853 10513 6867 10527
rect 8613 10513 8627 10527
rect 8773 10513 8787 10527
rect 10713 10513 10727 10527
rect 10773 10513 10787 10527
rect 653 10393 667 10407
rect 973 10393 987 10407
rect 1433 10393 1447 10407
rect 3053 10373 3067 10387
rect 3573 10393 3587 10407
rect 4433 10393 4447 10407
rect 5313 10393 5327 10407
rect 4373 10313 4387 10327
rect 4473 10313 4487 10327
rect 1473 10293 1487 10307
rect 1593 10293 1607 10307
rect 8413 10293 8427 10307
rect 8533 10293 8547 10307
rect 9193 10293 9207 10307
rect 9413 10292 9427 10306
rect 3473 10273 3487 10287
rect 3593 10273 3607 10287
rect 7993 10273 8007 10287
rect 8133 10273 8147 10287
rect 5233 10253 5247 10267
rect 5353 10233 5367 10247
rect 9313 10233 9327 10247
rect 9353 10233 9367 10247
rect 193 10213 207 10227
rect 353 10213 367 10227
rect 5253 10212 5267 10226
rect 5353 10212 5367 10226
rect 5473 10213 5487 10227
rect 5613 10213 5627 10227
rect 7733 10213 7747 10227
rect 7793 10213 7807 10227
rect 9333 10213 9347 10227
rect 9393 10213 9407 10227
rect 4393 10193 4407 10207
rect 4433 10193 4447 10207
rect 1153 10093 1167 10107
rect 1293 10093 1307 10107
rect 2853 10093 2867 10107
rect 2893 10093 2907 10107
rect 1073 10073 1087 10087
rect 1233 10073 1247 10087
rect 6973 10073 6987 10087
rect 7053 10073 7067 10087
rect 8933 10072 8947 10086
rect 9093 10073 9107 10087
rect 2533 10053 2547 10067
rect 4773 10053 4787 10067
rect 4853 10053 4867 10067
rect 5533 10053 5547 10067
rect 5613 10053 5627 10067
rect 7813 10053 7827 10067
rect 7933 10053 7947 10067
rect 2533 10013 2547 10027
rect 1113 9993 1127 10007
rect 1193 9993 1207 10007
rect 2253 9993 2267 10007
rect 2453 9993 2467 10007
rect 2733 9993 2747 10007
rect 2793 9993 2807 10007
rect 2873 9993 2887 10007
rect 3133 9993 3147 10007
rect 3193 9993 3207 10007
rect 4773 9993 4787 10007
rect 4933 9993 4947 10007
rect 6893 9993 6907 10007
rect 7073 9993 7087 10007
rect 8313 9993 8327 10007
rect 8433 9993 8447 10007
rect 10033 9993 10047 10007
rect 10073 9993 10087 10007
rect 1193 9972 1207 9986
rect 1293 9973 1307 9987
rect 333 9853 347 9867
rect 2433 9873 2447 9887
rect 5713 9853 5727 9867
rect 5773 9853 5787 9867
rect 353 9773 367 9787
rect 453 9773 467 9787
rect 1313 9773 1327 9787
rect 1373 9774 1387 9788
rect 3393 9773 3407 9787
rect 3493 9773 3507 9787
rect 4613 9773 4627 9787
rect 4773 9773 4787 9787
rect 2453 9753 2467 9767
rect 5693 9753 5707 9767
rect 5813 9753 5827 9767
rect 7573 9753 7587 9767
rect 7693 9753 7707 9767
rect 2313 9713 2327 9727
rect 2373 9713 2387 9727
rect 2453 9713 2467 9727
rect 3693 9713 3707 9727
rect 3753 9713 3767 9727
rect 6253 9713 6267 9727
rect 6293 9713 6307 9727
rect 6833 9713 6847 9727
rect 6953 9713 6967 9727
rect 7073 9713 7087 9727
rect 7173 9713 7187 9727
rect 7333 9713 7347 9727
rect 7453 9713 7467 9727
rect 7773 9693 7787 9707
rect 7833 9693 7847 9707
rect 1093 9573 1107 9587
rect 1173 9573 1187 9587
rect 1413 9553 1427 9567
rect 1473 9553 1487 9567
rect 3293 9552 3307 9566
rect 3413 9553 3427 9567
rect 4453 9553 4467 9567
rect 4513 9553 4527 9567
rect 10393 9553 10407 9567
rect 10593 9553 10607 9567
rect 2893 9533 2907 9547
rect 2993 9533 3007 9547
rect 9313 9533 9327 9547
rect 9433 9533 9447 9547
rect 5033 9513 5047 9527
rect 5113 9513 5127 9527
rect 7453 9513 7467 9527
rect 7513 9513 7527 9527
rect 2253 9493 2267 9507
rect 2313 9493 2327 9507
rect 4993 9493 5007 9507
rect 5913 9493 5927 9507
rect 6033 9493 6047 9507
rect 213 9473 227 9487
rect 413 9473 427 9487
rect 1313 9473 1327 9487
rect 1493 9473 1507 9487
rect 3873 9473 3887 9487
rect 3953 9473 3967 9487
rect 3993 9473 4007 9487
rect 4113 9473 4127 9487
rect 4453 9473 4467 9487
rect 4613 9473 4627 9487
rect 7153 9473 7167 9487
rect 7233 9473 7247 9487
rect 9473 9473 9487 9487
rect 9533 9473 9547 9487
rect 9753 9473 9767 9487
rect 9933 9471 9947 9485
rect 9973 9471 9987 9485
rect 10093 9473 10107 9487
rect 10213 9473 10227 9487
rect 10353 9473 10367 9487
rect 2953 9453 2967 9467
rect 2993 9452 3007 9466
rect 9133 9453 9147 9467
rect 9213 9453 9227 9467
rect 4753 9393 4767 9407
rect 4873 9393 4887 9407
rect 833 9353 847 9367
rect 1513 9353 1527 9367
rect 4913 9353 4927 9367
rect 9493 9353 9507 9367
rect 9713 9353 9727 9367
rect 10373 9353 10387 9367
rect 11253 9353 11267 9367
rect 3733 9333 3747 9347
rect 3773 9333 3787 9347
rect 3873 9333 3887 9347
rect 4933 9293 4947 9307
rect 5013 9293 5027 9307
rect 3213 9273 3227 9287
rect 3293 9273 3307 9287
rect 1273 9253 1287 9267
rect 1313 9253 1327 9267
rect 2853 9253 2867 9267
rect 2913 9253 2927 9267
rect 4053 9252 4067 9266
rect 4133 9254 4147 9268
rect 4233 9253 4247 9267
rect 4373 9253 4387 9267
rect 5413 9253 5427 9267
rect 5473 9253 5487 9267
rect 2833 9233 2847 9247
rect 2893 9233 2907 9247
rect 2993 9233 3007 9247
rect 2993 9193 3007 9207
rect 4113 9233 4127 9247
rect 5173 9233 5187 9247
rect 5273 9233 5287 9247
rect 4113 9193 4127 9207
rect 5693 9193 5707 9207
rect 5753 9193 5767 9207
rect 2373 9173 2387 9187
rect 2453 9173 2467 9187
rect 2573 9173 2587 9187
rect 2653 9173 2667 9187
rect 3513 9173 3527 9187
rect 3673 9173 3687 9187
rect 5113 9173 5127 9187
rect 5213 9173 5227 9187
rect 5253 9173 5267 9187
rect 5313 9171 5327 9185
rect 5653 9173 5667 9187
rect 5733 9172 5747 9186
rect 8493 9173 8507 9187
rect 8613 9173 8627 9187
rect 6093 9153 6107 9167
rect 6213 9153 6227 9167
rect 5153 9133 5167 9147
rect 5273 9133 5287 9147
rect 4993 9052 5007 9066
rect 5073 9053 5087 9067
rect 1413 9033 1427 9047
rect 1513 9033 1527 9047
rect 4673 9033 4687 9047
rect 4853 9033 4867 9047
rect 133 9013 147 9027
rect 4973 9013 4987 9027
rect 5013 9013 5027 9027
rect 5273 8993 5287 9007
rect 133 8973 147 8987
rect 5333 8973 5347 8987
rect 2673 8953 2687 8967
rect 2813 8953 2827 8967
rect 4933 8951 4947 8965
rect 5113 8953 5127 8967
rect 5193 8951 5207 8965
rect 5253 8953 5267 8967
rect 5653 8953 5667 8967
rect 5753 8953 5767 8967
rect 5853 8953 5867 8967
rect 6073 8951 6087 8965
rect 7493 8953 7507 8967
rect 7633 8953 7647 8967
rect 3573 8913 3587 8927
rect 3673 8913 3687 8927
rect 4733 8872 4747 8886
rect 4833 8873 4847 8887
rect 1033 8833 1047 8847
rect 3013 8833 3027 8847
rect 6933 8833 6947 8847
rect 2053 8813 2067 8827
rect 2093 8813 2107 8827
rect 8413 8813 8427 8827
rect 8653 8833 8667 8847
rect 9273 8833 9287 8847
rect 9613 8833 9627 8847
rect 10293 8833 10307 8847
rect 11313 8833 11327 8847
rect 8673 8813 8687 8827
rect 8713 8813 8727 8827
rect 4913 8793 4927 8807
rect 5013 8793 5027 8807
rect 4873 8773 4887 8787
rect 4913 8772 4927 8786
rect 2933 8733 2947 8747
rect 2993 8733 3007 8747
rect 4013 8733 4027 8747
rect 4073 8734 4087 8748
rect 4233 8733 4247 8747
rect 4313 8734 4327 8748
rect 4953 8733 4967 8747
rect 5033 8733 5047 8747
rect 5373 8733 5387 8747
rect 5473 8733 5487 8747
rect 5513 8733 5527 8747
rect 5773 8733 5787 8747
rect 5953 8733 5967 8747
rect 6093 8733 6107 8747
rect 6193 8734 6207 8748
rect 3933 8713 3947 8727
rect 4033 8713 4047 8727
rect 4153 8713 4167 8727
rect 4533 8713 4547 8727
rect 4153 8673 4167 8687
rect 4393 8673 4407 8687
rect 4773 8713 4787 8727
rect 4713 8672 4727 8686
rect 4873 8673 4887 8687
rect 4953 8673 4967 8687
rect 5113 8673 5127 8687
rect 5193 8673 5207 8687
rect 5333 8673 5347 8687
rect 5473 8673 5487 8687
rect 2773 8653 2787 8667
rect 2813 8653 2827 8667
rect 2873 8653 2887 8667
rect 4633 8653 4647 8667
rect 4813 8651 4827 8665
rect 6093 8653 6107 8667
rect 6133 8652 6147 8666
rect 2713 8633 2727 8647
rect 2833 8633 2847 8647
rect 5773 8632 5787 8646
rect 5813 8633 5827 8647
rect 6293 8633 6307 8647
rect 6333 8633 6347 8647
rect 3193 8613 3207 8627
rect 3313 8613 3327 8627
rect 5653 8613 5667 8627
rect 5693 8612 5707 8626
rect 4053 8553 4067 8567
rect 4133 8553 4147 8567
rect 6293 8553 6307 8567
rect 6413 8553 6427 8567
rect 4233 8533 4247 8547
rect 4333 8533 4347 8547
rect 6333 8533 6347 8547
rect 6393 8533 6407 8547
rect 213 8513 227 8527
rect 293 8513 307 8527
rect 3333 8513 3347 8527
rect 3473 8513 3487 8527
rect 4013 8514 4027 8528
rect 4173 8513 4187 8527
rect 4473 8513 4487 8527
rect 4513 8512 4527 8526
rect 4973 8513 4987 8527
rect 5153 8513 5167 8527
rect 6273 8513 6287 8527
rect 6353 8513 6367 8527
rect 3573 8493 3587 8507
rect 3693 8493 3707 8507
rect 9353 8493 9367 8507
rect 9473 8493 9487 8507
rect 3113 8453 3127 8467
rect 3213 8453 3227 8467
rect 3833 8453 3847 8467
rect 3933 8453 3947 8467
rect 4133 8453 4147 8467
rect 4193 8453 4207 8467
rect 4733 8453 4747 8467
rect 4853 8453 4867 8467
rect 5653 8453 5667 8467
rect 5753 8453 5767 8467
rect 6093 8453 6107 8467
rect 6133 8453 6147 8467
rect 10273 8453 10287 8467
rect 10373 8453 10387 8467
rect 1333 8433 1347 8447
rect 1393 8433 1407 8447
rect 4953 8433 4967 8447
rect 4993 8433 5007 8447
rect 5073 8433 5087 8447
rect 5133 8433 5147 8447
rect 5613 8433 5627 8447
rect 5833 8433 5847 8447
rect 6093 8432 6107 8446
rect 6153 8433 6167 8447
rect 7513 8432 7527 8446
rect 7613 8433 7627 8447
rect 8273 8433 8287 8447
rect 8313 8432 8327 8446
rect 9993 8433 10007 8447
rect 10113 8433 10127 8447
rect 10293 8433 10307 8447
rect 10433 8433 10447 8447
rect 5013 8353 5027 8367
rect 5093 8353 5107 8367
rect 6833 8313 6847 8327
rect 7433 8313 7447 8327
rect 7973 8313 7987 8327
rect 8093 8313 8107 8327
rect 8773 8313 8787 8327
rect 9953 8313 9967 8327
rect 10593 8313 10607 8327
rect 11313 8313 11327 8327
rect 373 8293 387 8307
rect 3913 8293 3927 8307
rect 3813 8273 3827 8287
rect 10593 8273 10607 8287
rect 10693 8273 10707 8287
rect 3093 8233 3107 8247
rect 1333 8213 1347 8227
rect 1473 8213 1487 8227
rect 1713 8213 1727 8227
rect 1813 8213 1827 8227
rect 3113 8213 3127 8227
rect 3553 8213 3567 8227
rect 3673 8213 3687 8227
rect 3993 8214 4007 8228
rect 4213 8214 4227 8228
rect 5093 8213 5107 8227
rect 5193 8213 5207 8227
rect 6213 8213 6227 8227
rect 6393 8213 6407 8227
rect 7113 8213 7127 8227
rect 7233 8213 7247 8227
rect 10573 8213 10587 8227
rect 10713 8213 10727 8227
rect 3813 8193 3827 8207
rect 3933 8193 3947 8207
rect 6333 8192 6347 8206
rect 6373 8193 6387 8207
rect 4093 8153 4107 8167
rect 4193 8153 4207 8167
rect 7073 8153 7087 8167
rect 7193 8153 7207 8167
rect 8233 8153 8247 8167
rect 8353 8153 8367 8167
rect 8433 8153 8447 8167
rect 8493 8153 8507 8167
rect 2413 8133 2427 8147
rect 2573 8133 2587 8147
rect 5773 8133 5787 8147
rect 5933 8133 5947 8147
rect 5973 8133 5987 8147
rect 6133 8133 6147 8147
rect 6253 8133 6267 8147
rect 6393 8133 6407 8147
rect 8553 8133 8567 8147
rect 8593 8133 8607 8147
rect 10073 8131 10087 8145
rect 10133 8133 10147 8147
rect 10173 8133 10187 8147
rect 10273 8133 10287 8147
rect 1113 8113 1127 8127
rect 1253 8113 1267 8127
rect 6433 8113 6447 8127
rect 6593 8113 6607 8127
rect 7353 8112 7367 8126
rect 7473 8113 7487 8127
rect 2893 8033 2907 8047
rect 5453 8033 5467 8047
rect 5553 8033 5567 8047
rect 2973 8013 2987 8027
rect 5493 8013 5507 8027
rect 5613 8013 5627 8027
rect 2373 7993 2387 8007
rect 2533 7994 2547 8008
rect 2673 7993 2687 8007
rect 2733 7993 2747 8007
rect 3733 7993 3747 8007
rect 3933 7993 3947 8007
rect 4693 7993 4707 8007
rect 4793 7993 4807 8007
rect 5193 7993 5207 8007
rect 5293 7993 5307 8007
rect 5893 7993 5907 8007
rect 6033 7993 6047 8007
rect 9893 7993 9907 8007
rect 9953 7993 9967 8007
rect 4993 7973 5007 7987
rect 5073 7973 5087 7987
rect 6433 7973 6447 7987
rect 6493 7973 6507 7987
rect 4093 7953 4107 7967
rect 4033 7933 4047 7947
rect 1833 7913 1847 7927
rect 1913 7913 1927 7927
rect 2293 7913 2307 7927
rect 2533 7913 2547 7927
rect 3053 7913 3067 7927
rect 3153 7913 3167 7927
rect 3753 7913 3767 7927
rect 3813 7913 3827 7927
rect 3973 7911 3987 7925
rect 4153 7913 4167 7927
rect 4193 7911 4207 7925
rect 4793 7913 4807 7927
rect 4913 7913 4927 7927
rect 5293 7913 5307 7927
rect 5393 7913 5407 7927
rect 4013 7893 4027 7907
rect 4173 7893 4187 7907
rect 4513 7892 4527 7906
rect 4633 7893 4647 7907
rect 8833 7873 8847 7887
rect 8913 7873 8927 7887
rect 2673 7833 2687 7847
rect 2753 7832 2767 7846
rect 3193 7833 3207 7847
rect 3233 7833 3247 7847
rect 3313 7833 3327 7847
rect 3373 7833 3387 7847
rect 4033 7833 4047 7847
rect 4153 7833 4167 7847
rect 4993 7833 5007 7847
rect 5033 7833 5047 7847
rect 1013 7793 1027 7807
rect 2513 7793 2527 7807
rect 2693 7773 2707 7787
rect 3253 7793 3267 7807
rect 6913 7793 6927 7807
rect 9013 7793 9027 7807
rect 9673 7793 9687 7807
rect 10273 7793 10287 7807
rect 11293 7773 11307 7787
rect 4313 7733 4327 7747
rect 4373 7732 4387 7746
rect 10073 7713 10087 7727
rect 10213 7713 10227 7727
rect 993 7693 1007 7707
rect 1073 7693 1087 7707
rect 2873 7693 2887 7707
rect 3073 7693 3087 7707
rect 3173 7693 3187 7707
rect 3313 7693 3327 7707
rect 4133 7693 4147 7707
rect 4233 7693 4247 7707
rect 4353 7692 4367 7706
rect 4453 7693 4467 7707
rect 4793 7693 4807 7707
rect 4933 7693 4947 7707
rect 7193 7693 7207 7707
rect 7253 7693 7267 7707
rect 7293 7693 7307 7707
rect 8733 7693 8747 7707
rect 8853 7693 8867 7707
rect 8913 7693 8927 7707
rect 9653 7693 9667 7707
rect 9813 7693 9827 7707
rect 10113 7693 10127 7707
rect 10253 7693 10267 7707
rect 10353 7693 10367 7707
rect 10453 7693 10467 7707
rect 10573 7693 10587 7707
rect 10773 7693 10787 7707
rect 2653 7673 2667 7687
rect 4533 7673 4547 7687
rect 4613 7673 4627 7687
rect 5413 7673 5427 7687
rect 10593 7673 10607 7687
rect 1813 7633 1827 7647
rect 1853 7633 1867 7647
rect 2793 7633 2807 7647
rect 5033 7633 5047 7647
rect 5113 7633 5127 7647
rect 10613 7652 10627 7666
rect 10713 7673 10727 7687
rect 7273 7633 7287 7647
rect 7353 7633 7367 7647
rect 7633 7633 7647 7647
rect 7733 7633 7747 7647
rect 10713 7633 10727 7647
rect 2413 7613 2427 7627
rect 2493 7613 2507 7627
rect 2573 7613 2587 7627
rect 3153 7613 3167 7627
rect 3273 7613 3287 7627
rect 4793 7613 4807 7627
rect 4873 7612 4887 7626
rect 5413 7613 5427 7627
rect 7273 7612 7287 7626
rect 7373 7613 7387 7627
rect 7613 7613 7627 7627
rect 7693 7613 7707 7627
rect 7733 7612 7747 7626
rect 9673 7613 9687 7627
rect 9773 7613 9787 7627
rect 9833 7613 9847 7627
rect 10613 7613 10627 7627
rect 10733 7613 10747 7627
rect 5433 7593 5447 7607
rect 5573 7593 5587 7607
rect 7013 7573 7027 7587
rect 7093 7573 7107 7587
rect 433 7493 447 7507
rect 553 7493 567 7507
rect 9613 7493 9627 7507
rect 1513 7473 1527 7487
rect 1633 7473 1647 7487
rect 2613 7473 2627 7487
rect 2793 7473 2807 7487
rect 4973 7473 4987 7487
rect 1653 7453 1667 7467
rect 6073 7473 6087 7487
rect 6233 7473 6247 7487
rect 7533 7472 7547 7486
rect 7633 7473 7647 7487
rect 9713 7473 9727 7487
rect 10913 7473 10927 7487
rect 11113 7473 11127 7487
rect 1633 7432 1647 7446
rect 5453 7453 5467 7467
rect 5053 7432 5067 7446
rect 5453 7413 5467 7427
rect 8433 7413 8447 7427
rect 8533 7413 8547 7427
rect 2013 7393 2027 7407
rect 2093 7393 2107 7407
rect 4953 7393 4967 7407
rect 5173 7393 5187 7407
rect 5713 7393 5727 7407
rect 5833 7393 5847 7407
rect 6833 7393 6847 7407
rect 6973 7393 6987 7407
rect 8973 7393 8987 7407
rect 9033 7393 9047 7407
rect 9173 7393 9187 7407
rect 9253 7393 9267 7407
rect 10733 7393 10747 7407
rect 10853 7393 10867 7407
rect 1973 7373 1987 7387
rect 2073 7373 2087 7387
rect 5653 7373 5667 7387
rect 5733 7373 5747 7387
rect 8893 7373 8907 7387
rect 8953 7373 8967 7387
rect 10493 7373 10507 7387
rect 10633 7373 10647 7387
rect 5293 7353 5307 7367
rect 5353 7352 5367 7366
rect 1373 7253 1387 7267
rect 2113 7273 2127 7287
rect 4933 7273 4947 7287
rect 7733 7273 7747 7287
rect 8373 7273 8387 7287
rect 9893 7273 9907 7287
rect 2033 7253 2047 7267
rect 2133 7253 2147 7267
rect 9793 7253 9807 7267
rect 9893 7252 9907 7266
rect 4173 7173 4187 7187
rect 4293 7172 4307 7186
rect 9933 7173 9947 7187
rect 9993 7173 10007 7187
rect 693 7153 707 7167
rect 753 7153 767 7167
rect 813 7153 827 7167
rect 3913 7153 3927 7167
rect 4053 7153 4067 7167
rect 5193 7153 5207 7167
rect 7553 7133 7567 7147
rect 7593 7133 7607 7147
rect 2713 7113 2727 7127
rect 2853 7113 2867 7127
rect 5193 7113 5207 7127
rect 5593 7113 5607 7127
rect 5733 7113 5747 7127
rect 5793 7113 5807 7127
rect 6493 7113 6507 7127
rect 6593 7113 6607 7127
rect 6673 7113 6687 7127
rect 6793 7113 6807 7127
rect 7813 7113 7827 7127
rect 7873 7113 7887 7127
rect 3453 7093 3467 7107
rect 3513 7092 3527 7106
rect 5593 7092 5607 7106
rect 5693 7093 5707 7107
rect 6653 7093 6667 7107
rect 6753 7093 6767 7107
rect 9633 7093 9647 7107
rect 9733 7093 9747 7107
rect 5613 7073 5627 7087
rect 8873 7073 8887 7087
rect 8913 7072 8927 7086
rect 3193 7053 3207 7067
rect 3313 7053 3327 7067
rect 5213 6993 5227 7007
rect 5313 6993 5327 7007
rect 5453 6993 5467 7007
rect 5593 6993 5607 7007
rect 5233 6973 5247 6987
rect 5293 6973 5307 6987
rect 6093 6973 6107 6987
rect 6253 6973 6267 6987
rect 2493 6953 2507 6967
rect 2633 6953 2647 6967
rect 4093 6953 4107 6967
rect 4173 6953 4187 6967
rect 4353 6953 4367 6967
rect 4393 6953 4407 6967
rect 4593 6953 4607 6967
rect 4733 6953 4747 6967
rect 4973 6953 4987 6967
rect 5173 6953 5187 6967
rect 5833 6954 5847 6968
rect 5933 6953 5947 6967
rect 7113 6953 7127 6967
rect 7173 6953 7187 6967
rect 8853 6953 8867 6967
rect 9053 6953 9067 6967
rect 4333 6933 4347 6947
rect 4413 6933 4427 6947
rect 7613 6933 7627 6947
rect 7673 6933 7687 6947
rect 9473 6933 9487 6947
rect 9513 6933 9527 6947
rect 6333 6893 6347 6907
rect 6433 6893 6447 6907
rect 7353 6893 7367 6907
rect 7413 6893 7427 6907
rect 7533 6893 7547 6907
rect 7613 6893 7627 6907
rect 2533 6873 2547 6887
rect 3793 6873 3807 6887
rect 3873 6873 3887 6887
rect 3913 6873 3927 6887
rect 6313 6873 6327 6887
rect 6433 6872 6447 6886
rect 7373 6873 7387 6887
rect 7453 6873 7467 6887
rect 8913 6873 8927 6887
rect 9033 6873 9047 6887
rect 9593 6873 9607 6887
rect 9653 6873 9667 6887
rect 2573 6852 2587 6866
rect 3713 6852 3727 6866
rect 3833 6853 3847 6867
rect 3873 6852 3887 6866
rect 3993 6853 4007 6867
rect 4253 6853 4267 6867
rect 6353 6853 6367 6867
rect 6453 6853 6467 6867
rect 2653 6833 2667 6847
rect 2693 6833 2707 6847
rect 4153 6833 4167 6847
rect 573 6753 587 6767
rect 1273 6753 1287 6767
rect 3293 6753 3307 6767
rect 4513 6753 4527 6767
rect 7213 6753 7227 6767
rect 9533 6753 9547 6767
rect 9873 6753 9887 6767
rect 10673 6753 10687 6767
rect 10893 6753 10907 6767
rect 11133 6733 11147 6747
rect 11193 6733 11207 6747
rect 3073 6713 3087 6727
rect 2913 6693 2927 6707
rect 5473 6693 5487 6707
rect 5533 6693 5547 6707
rect 2273 6653 2287 6667
rect 2393 6653 2407 6667
rect 9853 6653 9867 6667
rect 9913 6653 9927 6667
rect 3193 6633 3207 6647
rect 3293 6633 3307 6647
rect 10673 6613 10687 6627
rect 10713 6613 10727 6627
rect 5433 6593 5447 6607
rect 5473 6593 5487 6607
rect 7973 6593 7987 6607
rect 8113 6593 8127 6607
rect 8633 6593 8647 6607
rect 8753 6593 8767 6607
rect 9093 6593 9107 6607
rect 9153 6593 9167 6607
rect 2033 6573 2047 6587
rect 2113 6573 2127 6587
rect 3833 6573 3847 6587
rect 3933 6573 3947 6587
rect 5453 6572 5467 6586
rect 5553 6573 5567 6587
rect 6433 6573 6447 6587
rect 6473 6572 6487 6586
rect 6653 6572 6667 6586
rect 6693 6573 6707 6587
rect 8833 6573 8847 6587
rect 8893 6573 8907 6587
rect 8933 6573 8947 6587
rect 9353 6573 9367 6587
rect 9453 6573 9467 6587
rect 10993 6573 11007 6587
rect 11033 6573 11047 6587
rect 3853 6553 3867 6567
rect 3933 6552 3947 6566
rect 7993 6553 8007 6567
rect 8093 6552 8107 6566
rect 3153 6533 3167 6547
rect 3273 6533 3287 6547
rect 2533 6453 2547 6467
rect 2573 6453 2587 6467
rect 2653 6433 2667 6447
rect 2793 6433 2807 6447
rect 4073 6433 4087 6447
rect 4213 6433 4227 6447
rect 4333 6433 4347 6447
rect 4513 6433 4527 6447
rect 8293 6433 8307 6447
rect 8393 6433 8407 6447
rect 8813 6433 8827 6447
rect 2953 6413 2967 6427
rect 3013 6413 3027 6427
rect 3893 6413 3907 6427
rect 3973 6412 3987 6426
rect 8093 6413 8107 6427
rect 8853 6413 8867 6427
rect 9713 6413 9727 6427
rect 9813 6413 9827 6427
rect 9853 6413 9867 6427
rect 2953 6373 2967 6387
rect 3013 6373 3027 6387
rect 433 6353 447 6367
rect 533 6353 547 6367
rect 2553 6353 2567 6367
rect 2613 6353 2627 6367
rect 2713 6352 2727 6366
rect 2773 6353 2787 6367
rect 3633 6353 3647 6367
rect 3693 6353 3707 6367
rect 3773 6353 3787 6367
rect 3813 6353 3827 6367
rect 4573 6351 4587 6365
rect 4713 6353 4727 6367
rect 5133 6353 5147 6367
rect 5212 6353 5226 6367
rect 5233 6353 5247 6367
rect 5373 6353 5387 6367
rect 6193 6353 6207 6367
rect 6273 6353 6287 6367
rect 6413 6353 6427 6367
rect 6633 6353 6647 6367
rect 6673 6353 6687 6367
rect 6773 6353 6787 6367
rect 6813 6353 6827 6367
rect 8113 6352 8127 6366
rect 8293 6353 8307 6367
rect 8513 6353 8527 6367
rect 9693 6353 9707 6367
rect 9913 6353 9927 6367
rect 2413 6333 2427 6347
rect 2553 6332 2567 6346
rect 6313 6333 6327 6347
rect 6373 6333 6387 6347
rect 1293 6233 1307 6247
rect 1933 6233 1947 6247
rect 7973 6233 7987 6247
rect 5973 6213 5987 6227
rect 6933 6213 6947 6227
rect 6993 6213 7007 6227
rect 8593 6213 8607 6227
rect 10433 6213 10447 6227
rect 7653 6173 7667 6187
rect 7733 6172 7747 6186
rect 1393 6133 1407 6147
rect 1573 6133 1587 6147
rect 3673 6133 3687 6147
rect 3893 6133 3907 6147
rect 5893 6133 5907 6147
rect 6013 6133 6027 6147
rect 6853 6133 6867 6147
rect 6893 6134 6907 6148
rect 8293 6133 8307 6147
rect 8453 6133 8467 6147
rect 8793 6133 8807 6147
rect 8953 6133 8967 6147
rect 10233 6133 10247 6147
rect 10313 6134 10327 6148
rect 10413 6133 10427 6147
rect 10533 6133 10547 6147
rect 1173 6113 1187 6127
rect 1213 6113 1227 6127
rect 5313 6113 5327 6127
rect 5913 6113 5927 6127
rect 5993 6113 6007 6127
rect 6513 6113 6527 6127
rect 6553 6113 6567 6127
rect 6993 6113 7007 6127
rect 7073 6113 7087 6127
rect 9713 6113 9727 6127
rect 10913 6113 10927 6127
rect 10973 6113 10987 6127
rect 2693 6093 2707 6107
rect 2553 6073 2567 6087
rect 2713 6073 2727 6087
rect 3493 6073 3507 6087
rect 3533 6073 3547 6087
rect 5313 6073 5327 6087
rect 6513 6073 6527 6087
rect 6553 6073 6567 6087
rect 9573 6073 9587 6087
rect 9713 6073 9727 6087
rect 9933 6073 9947 6087
rect 10053 6073 10067 6087
rect 1673 6053 1687 6067
rect 1773 6053 1787 6067
rect 3753 6053 3767 6067
rect 3893 6051 3907 6065
rect 3933 6053 3947 6067
rect 4073 6053 4087 6067
rect 6533 6053 6547 6067
rect 6673 6053 6687 6067
rect 9613 6053 9627 6067
rect 10733 6053 10747 6067
rect 10793 6053 10807 6067
rect 8113 6013 8127 6027
rect 8253 6013 8267 6027
rect 11093 6013 11107 6027
rect 11193 6012 11207 6026
rect 10873 5933 10887 5947
rect 10973 5932 10987 5946
rect 5013 5913 5027 5927
rect 5053 5913 5067 5927
rect 7633 5912 7647 5926
rect 7713 5913 7727 5927
rect 1433 5893 1447 5907
rect 1513 5893 1527 5907
rect 2593 5893 2607 5907
rect 2653 5893 2667 5907
rect 4633 5893 4647 5907
rect 6033 5893 6047 5907
rect 6093 5893 6107 5907
rect 7813 5893 7827 5907
rect 7873 5893 7887 5907
rect 7953 5893 7967 5907
rect 11093 5893 11107 5907
rect 1873 5833 1887 5847
rect 3113 5833 3127 5847
rect 3153 5833 3167 5847
rect 3853 5833 3867 5847
rect 3973 5833 3987 5847
rect 6733 5853 6747 5867
rect 6813 5853 6827 5867
rect 7813 5853 7827 5867
rect 11093 5853 11107 5867
rect 4653 5833 4667 5847
rect 6233 5831 6247 5845
rect 6333 5833 6347 5847
rect 10853 5831 10867 5845
rect 10973 5833 10987 5847
rect 11073 5833 11087 5847
rect 11233 5833 11247 5847
rect 2073 5813 2087 5827
rect 6473 5753 6487 5767
rect 6613 5753 6627 5767
rect 553 5713 567 5727
rect 4453 5713 4467 5727
rect 4693 5713 4707 5727
rect 5773 5713 5787 5727
rect 9233 5713 9247 5727
rect 9373 5713 9387 5727
rect 10053 5713 10067 5727
rect 11313 5713 11327 5727
rect 11293 5653 11307 5667
rect 11273 5633 11287 5647
rect 713 5613 727 5627
rect 873 5613 887 5627
rect 1093 5613 1107 5627
rect 1153 5613 1167 5627
rect 1793 5613 1807 5627
rect 1873 5613 1887 5627
rect 2053 5613 2067 5627
rect 2153 5613 2167 5627
rect 2593 5613 2607 5627
rect 2773 5613 2787 5627
rect 3273 5613 3287 5627
rect 3313 5613 3327 5627
rect 4133 5613 4147 5627
rect 4193 5612 4207 5626
rect 5053 5613 5067 5627
rect 4473 5593 4487 5607
rect 4513 5593 4527 5607
rect 5113 5613 5127 5627
rect 5173 5612 5187 5626
rect 5813 5613 5827 5627
rect 5893 5613 5907 5627
rect 6013 5613 6027 5627
rect 6113 5613 6127 5627
rect 6913 5613 6927 5627
rect 6953 5613 6967 5627
rect 5113 5573 5127 5587
rect 11293 5613 11307 5627
rect 4133 5553 4147 5567
rect 4173 5553 4187 5567
rect 7193 5553 7207 5567
rect 7313 5553 7327 5567
rect 11293 5552 11307 5566
rect 1133 5533 1147 5547
rect 1293 5533 1307 5547
rect 1533 5533 1547 5547
rect 1693 5533 1707 5547
rect 9413 5533 9427 5547
rect 9593 5533 9607 5547
rect 1933 5493 1947 5507
rect 1993 5493 2007 5507
rect 2653 5433 2667 5447
rect 2793 5433 2807 5447
rect 2853 5433 2867 5447
rect 2993 5433 3007 5447
rect 5793 5433 5807 5447
rect 5913 5433 5927 5447
rect 7833 5412 7847 5426
rect 7893 5413 7907 5427
rect 2313 5393 2327 5407
rect 1493 5373 1507 5387
rect 1593 5373 1607 5387
rect 2413 5393 2427 5407
rect 6253 5392 6267 5406
rect 6393 5394 6407 5408
rect 2513 5373 2527 5387
rect 6213 5373 6227 5387
rect 6313 5373 6327 5387
rect 8293 5373 8307 5387
rect 10173 5373 10187 5387
rect 1113 5313 1127 5327
rect 1373 5313 1387 5327
rect 1533 5313 1547 5327
rect 1653 5313 1667 5327
rect 2113 5313 2127 5327
rect 2753 5333 2767 5347
rect 2793 5333 2807 5347
rect 8133 5333 8147 5347
rect 8213 5333 8227 5347
rect 8293 5333 8307 5347
rect 10293 5333 10307 5347
rect 2233 5293 2247 5307
rect 2273 5293 2287 5307
rect 2373 5313 2387 5327
rect 5773 5313 5787 5327
rect 5813 5313 5827 5327
rect 6053 5313 6067 5327
rect 6153 5313 6167 5327
rect 6193 5313 6207 5327
rect 6413 5313 6427 5327
rect 6753 5313 6767 5327
rect 6833 5311 6847 5325
rect 7853 5313 7867 5327
rect 7993 5311 8007 5325
rect 8273 5313 8287 5327
rect 8393 5313 8407 5327
rect 9193 5313 9207 5327
rect 9233 5313 9247 5327
rect 2333 5293 2347 5307
rect 3033 5293 3047 5307
rect 3193 5293 3207 5307
rect 4213 5292 4227 5306
rect 4253 5293 4267 5307
rect 2193 5272 2207 5286
rect 2293 5273 2307 5287
rect 6813 5273 6827 5287
rect 6753 5253 6767 5267
rect 2673 5233 2687 5247
rect 2773 5233 2787 5247
rect 6693 5233 6707 5247
rect 6793 5233 6807 5247
rect 6913 5233 6927 5247
rect 7013 5233 7027 5247
rect 4153 5193 4167 5207
rect 5013 5193 5027 5207
rect 5953 5193 5967 5207
rect 7753 5193 7767 5207
rect 9513 5193 9527 5207
rect 9633 5193 9647 5207
rect 10633 5193 10647 5207
rect 10713 5193 10727 5207
rect 11173 5193 11187 5207
rect 2113 5173 2127 5187
rect 2253 5173 2267 5187
rect 2573 5173 2587 5187
rect 2673 5173 2687 5187
rect 2133 5153 2147 5167
rect 2233 5153 2247 5167
rect 10713 5153 10727 5167
rect 10773 5153 10787 5167
rect 6533 5133 6547 5147
rect 6693 5113 6707 5127
rect 9913 5113 9927 5127
rect 9953 5113 9967 5127
rect 513 5093 527 5107
rect 733 5093 747 5107
rect 1633 5093 1647 5107
rect 1733 5093 1747 5107
rect 1973 5093 1987 5107
rect 2053 5093 2067 5107
rect 2553 5093 2567 5107
rect 2713 5093 2727 5107
rect 2973 5093 2987 5107
rect 3053 5093 3067 5107
rect 3193 5093 3207 5107
rect 5073 5093 5087 5107
rect 5153 5093 5167 5107
rect 6293 5093 6307 5107
rect 6413 5093 6427 5107
rect 6573 5093 6587 5107
rect 6693 5092 6707 5106
rect 8813 5093 8827 5107
rect 8913 5093 8927 5107
rect 10893 5093 10907 5107
rect 11013 5093 11027 5107
rect 11133 5093 11147 5107
rect 11233 5093 11247 5107
rect 2473 5073 2487 5087
rect 2573 5073 2587 5087
rect 2673 5073 2687 5087
rect 6533 5073 6547 5087
rect 6653 5073 6667 5087
rect 2773 5033 2787 5047
rect 2813 5033 2827 5047
rect 4553 5033 4567 5047
rect 5033 5033 5047 5047
rect 5113 5033 5127 5047
rect 5653 5033 5667 5047
rect 5813 5033 5827 5047
rect 8633 5033 8647 5047
rect 8733 5033 8747 5047
rect 8853 5033 8867 5047
rect 1893 5013 1907 5027
rect 2053 5013 2067 5027
rect 2453 5013 2467 5027
rect 2833 5013 2847 5027
rect 2933 5013 2947 5027
rect 4533 5013 4547 5027
rect 4573 5013 4587 5027
rect 4653 5013 4667 5027
rect 4953 5013 4967 5027
rect 5033 5012 5047 5026
rect 8973 5013 8987 5027
rect 10813 5013 10827 5027
rect 10973 5013 10987 5027
rect 2333 4993 2347 5007
rect 6113 4993 6127 5007
rect 2393 4973 2407 4987
rect 4113 4972 4127 4986
rect 4153 4973 4167 4987
rect 6233 4973 6247 4987
rect 2673 4913 2687 4927
rect 2773 4913 2787 4927
rect 7233 4913 7247 4927
rect 7313 4912 7327 4926
rect 5353 4893 5367 4907
rect 5473 4893 5487 4907
rect 1893 4873 1907 4887
rect 1993 4873 2007 4887
rect 2173 4873 2187 4887
rect 2273 4873 2287 4887
rect 6213 4873 6227 4887
rect 6313 4873 6327 4887
rect 6473 4874 6487 4888
rect 6613 4873 6627 4887
rect 2173 4852 2187 4866
rect 2293 4853 2307 4867
rect 4873 4853 4887 4867
rect 4993 4853 5007 4867
rect 6073 4853 6087 4867
rect 6173 4853 6187 4867
rect 7333 4873 7347 4887
rect 8133 4853 8147 4867
rect 7233 4833 7247 4847
rect 8873 4853 8887 4867
rect 8913 4853 8927 4867
rect 8273 4813 8287 4827
rect 2433 4793 2447 4807
rect 2573 4791 2587 4805
rect 2933 4793 2947 4807
rect 2973 4793 2987 4807
rect 6213 4793 6227 4807
rect 6273 4793 6287 4807
rect 11113 4793 11127 4807
rect 11313 4793 11327 4807
rect 1933 4773 1947 4787
rect 2073 4773 2087 4787
rect 3313 4773 3327 4787
rect 3393 4773 3407 4787
rect 11133 4773 11147 4787
rect 11173 4773 11187 4787
rect 1673 4753 1687 4767
rect 1773 4752 1787 4766
rect 4293 4673 4307 4687
rect 2073 4653 2087 4667
rect 2213 4653 2227 4667
rect 6833 4653 6847 4667
rect 8933 4673 8947 4687
rect 9333 4673 9347 4687
rect 11053 4673 11067 4687
rect 7273 4653 7287 4667
rect 7313 4653 7327 4667
rect 1873 4613 1887 4627
rect 1953 4613 1967 4627
rect 3053 4613 3067 4627
rect 3113 4613 3127 4627
rect 6753 4613 6767 4627
rect 6833 4613 6847 4627
rect 2053 4593 2067 4607
rect 2273 4593 2287 4607
rect 9593 4593 9607 4607
rect 9653 4593 9667 4607
rect 653 4573 667 4587
rect 753 4573 767 4587
rect 1593 4573 1607 4587
rect 1673 4573 1687 4587
rect 1773 4573 1787 4587
rect 1853 4573 1867 4587
rect 1933 4573 1947 4587
rect 2013 4573 2027 4587
rect 2953 4573 2967 4587
rect 3113 4573 3127 4587
rect 4853 4573 4867 4587
rect 4893 4573 4907 4587
rect 6073 4574 6087 4588
rect 6193 4573 6207 4587
rect 6553 4573 6567 4587
rect 6613 4573 6627 4587
rect 5853 4553 5867 4567
rect 5993 4553 6007 4567
rect 9313 4553 9327 4567
rect 9393 4553 9407 4567
rect 11233 4553 11247 4567
rect 11293 4553 11307 4567
rect 7253 4532 7267 4546
rect 7313 4533 7327 4547
rect 3613 4513 3627 4527
rect 3733 4513 3747 4527
rect 5693 4513 5707 4527
rect 5753 4513 5767 4527
rect 2953 4473 2967 4487
rect 3053 4473 3067 4487
rect 6613 4453 6627 4467
rect 6713 4453 6727 4467
rect 3773 4393 3787 4407
rect 3893 4393 3907 4407
rect 3853 4353 3867 4367
rect 3913 4353 3927 4367
rect 8393 4353 8407 4367
rect 8473 4353 8487 4367
rect 2953 4333 2967 4347
rect 3753 4333 3767 4347
rect 3873 4333 3887 4347
rect 4893 4333 4907 4347
rect 5013 4333 5027 4347
rect 2913 4312 2927 4326
rect 2393 4293 2407 4307
rect 3533 4293 3547 4307
rect 3633 4293 3647 4307
rect 7413 4293 7427 4307
rect 7453 4293 7467 4307
rect 2553 4273 2567 4287
rect 3033 4273 3047 4287
rect 3233 4273 3247 4287
rect 3513 4273 3527 4287
rect 3553 4273 3567 4287
rect 4413 4273 4427 4287
rect 4573 4273 4587 4287
rect 4773 4273 4787 4287
rect 4833 4273 4847 4287
rect 4973 4273 4987 4287
rect 5073 4273 5087 4287
rect 6133 4273 6147 4287
rect 6193 4273 6207 4287
rect 6613 4273 6627 4287
rect 6833 4273 6847 4287
rect 6873 4273 6887 4287
rect 7053 4273 7067 4287
rect 7153 4273 7167 4287
rect 7233 4273 7247 4287
rect 2393 4253 2407 4267
rect 2513 4253 2527 4267
rect 6073 4253 6087 4267
rect 6173 4253 6187 4267
rect 2213 4213 2227 4227
rect 2253 4212 2267 4226
rect 3193 4213 3207 4227
rect 3093 4193 3107 4207
rect 4473 4193 4487 4207
rect 4553 4193 4567 4207
rect 7193 4192 7207 4206
rect 7293 4193 7307 4207
rect 4553 4133 4567 4147
rect 4673 4133 4687 4147
rect 11233 4133 11247 4147
rect 1673 4093 1687 4107
rect 1713 4093 1727 4107
rect 3093 4073 3107 4087
rect 3133 4073 3147 4087
rect 1073 4053 1087 4067
rect 1333 4053 1347 4067
rect 2673 4053 2687 4067
rect 2753 4053 2767 4067
rect 3233 4053 3247 4067
rect 3393 4053 3407 4067
rect 3693 4053 3707 4067
rect 3833 4053 3847 4067
rect 4213 4053 4227 4067
rect 4293 4053 4307 4067
rect 5713 4053 5727 4067
rect 5893 4054 5907 4068
rect 6913 4053 6927 4067
rect 7093 4053 7107 4067
rect 8073 4053 8087 4067
rect 8213 4053 8227 4067
rect 3013 4033 3027 4047
rect 3133 4033 3147 4047
rect 3373 4033 3387 4047
rect 7673 4032 7687 4046
rect 7713 4033 7727 4047
rect 3573 4013 3587 4027
rect 2793 3993 2807 4007
rect 3373 3993 3387 4007
rect 3453 3993 3467 4007
rect 4333 3993 4347 4007
rect 4453 3993 4467 4007
rect 6933 3993 6947 4007
rect 7033 3993 7047 4007
rect 8873 3993 8887 4007
rect 8913 3993 8927 4007
rect 8993 3993 9007 4007
rect 9053 3993 9067 4007
rect 1233 3973 1247 3987
rect 1273 3973 1287 3987
rect 1633 3973 1647 3987
rect 1713 3973 1727 3987
rect 2933 3973 2947 3987
rect 4893 3973 4907 3987
rect 4953 3971 4967 3985
rect 9853 3971 9867 3985
rect 9953 3973 9967 3987
rect 3873 3953 3887 3967
rect 4033 3953 4047 3967
rect 6653 3953 6667 3967
rect 6793 3933 6807 3947
rect 2773 3873 2787 3887
rect 2873 3873 2887 3887
rect 3893 3873 3907 3887
rect 5773 3873 5787 3887
rect 1213 3853 1227 3867
rect 2733 3853 2747 3867
rect 2853 3853 2867 3867
rect 3153 3853 3167 3867
rect 3273 3853 3287 3867
rect 5853 3872 5867 3886
rect 4013 3853 4027 3867
rect 1313 3833 1327 3847
rect 2573 3833 2587 3847
rect 2693 3833 2707 3847
rect 3413 3833 3427 3847
rect 3533 3833 3547 3847
rect 4093 3833 4107 3847
rect 4133 3833 4147 3847
rect 553 3813 567 3827
rect 633 3813 647 3827
rect 3433 3813 3447 3827
rect 3553 3813 3567 3827
rect 3693 3813 3707 3827
rect 3793 3813 3807 3827
rect 7453 3813 7467 3827
rect 2293 3773 2307 3787
rect 2373 3773 2387 3787
rect 2573 3773 2587 3787
rect 2753 3773 2767 3787
rect 2853 3773 2867 3787
rect 3173 3773 3187 3787
rect 3253 3773 3267 3787
rect 7453 3773 7467 3787
rect 1213 3752 1227 3766
rect 1293 3753 1307 3767
rect 2173 3753 2187 3767
rect 2233 3753 2247 3767
rect 2333 3753 2347 3767
rect 2373 3752 2387 3766
rect 2513 3753 2527 3767
rect 2553 3753 2567 3767
rect 2693 3753 2707 3767
rect 4093 3753 4107 3767
rect 4213 3753 4227 3767
rect 7073 3753 7087 3767
rect 7153 3753 7167 3767
rect 7253 3753 7267 3767
rect 7693 3834 7707 3848
rect 8413 3833 8427 3847
rect 8573 3833 8587 3847
rect 10453 3833 10467 3847
rect 10573 3833 10587 3847
rect 7673 3813 7687 3827
rect 7673 3773 7687 3787
rect 9193 3773 9207 3787
rect 9313 3773 9327 3787
rect 9353 3773 9367 3787
rect 10893 3773 10907 3787
rect 11013 3773 11027 3787
rect 7693 3753 7707 3767
rect 9093 3753 9107 3767
rect 9293 3753 9307 3767
rect 10873 3751 10887 3765
rect 10993 3753 11007 3767
rect 11073 3753 11087 3767
rect 7133 3733 7147 3747
rect 7193 3733 7207 3747
rect 3013 3713 3027 3727
rect 3053 3713 3067 3727
rect 2953 3673 2967 3687
rect 2993 3673 3007 3687
rect 6353 3633 6367 3647
rect 7033 3633 7047 3647
rect 8113 3633 8127 3647
rect 9053 3633 9067 3647
rect 10173 3633 10187 3647
rect 10233 3633 10247 3647
rect 2933 3612 2947 3626
rect 3013 3613 3027 3627
rect 4513 3613 4527 3627
rect 4573 3613 4587 3627
rect 1873 3573 1887 3587
rect 1913 3573 1927 3587
rect 3333 3573 3347 3587
rect 3473 3572 3487 3586
rect 2253 3553 2267 3567
rect 2453 3553 2467 3567
rect 4893 3553 4907 3567
rect 5033 3553 5047 3567
rect 9913 3553 9927 3567
rect 10033 3553 10047 3567
rect 1893 3533 1907 3547
rect 1973 3533 1987 3547
rect 2493 3533 2507 3547
rect 2633 3533 2647 3547
rect 3073 3533 3087 3547
rect 3113 3533 3127 3547
rect 3533 3534 3547 3548
rect 3673 3533 3687 3547
rect 3793 3533 3807 3547
rect 3913 3533 3927 3547
rect 3953 3533 3967 3547
rect 4093 3533 4107 3547
rect 4773 3533 4787 3547
rect 4833 3533 4847 3547
rect 7693 3533 7707 3547
rect 7753 3533 7767 3547
rect 9093 3533 9107 3547
rect 1393 3513 1407 3527
rect 1473 3513 1487 3527
rect 1513 3513 1527 3527
rect 3473 3513 3487 3527
rect 5573 3513 5587 3527
rect 5653 3513 5667 3527
rect 8973 3513 8987 3527
rect 9633 3513 9647 3527
rect 9773 3513 9787 3527
rect 1153 3473 1167 3487
rect 1293 3473 1307 3487
rect 2973 3473 2987 3487
rect 3013 3473 3027 3487
rect 3333 3473 3347 3487
rect 3373 3473 3387 3487
rect 3473 3473 3487 3487
rect 4333 3473 4347 3487
rect 4393 3473 4407 3487
rect 4673 3473 4687 3487
rect 4753 3473 4767 3487
rect 1053 3453 1067 3467
rect 1093 3451 1107 3465
rect 1213 3453 1227 3467
rect 1293 3452 1307 3466
rect 3533 3453 3547 3467
rect 3593 3453 3607 3467
rect 1813 3433 1827 3447
rect 1933 3432 1947 3446
rect 2853 3433 2867 3447
rect 3033 3432 3047 3446
rect 3773 3432 3787 3446
rect 3813 3433 3827 3447
rect 8973 3433 8987 3447
rect 9113 3433 9127 3447
rect 10173 3433 10187 3447
rect 10233 3433 10247 3447
rect 3433 3413 3447 3427
rect 3473 3413 3487 3427
rect 9633 3413 9647 3427
rect 9773 3413 9787 3427
rect 1813 3353 1827 3367
rect 1913 3353 1927 3367
rect 2713 3353 2727 3367
rect 2773 3353 2787 3367
rect 3013 3353 3027 3367
rect 3093 3353 3107 3367
rect 4393 3353 4407 3367
rect 4533 3353 4547 3367
rect 10673 3353 10687 3367
rect 10713 3353 10727 3367
rect 4133 3333 4147 3347
rect 4173 3333 4187 3347
rect 1033 3313 1047 3327
rect 1213 3313 1227 3327
rect 1573 3313 1587 3327
rect 1673 3313 1687 3327
rect 3653 3314 3667 3328
rect 3733 3313 3747 3327
rect 4593 3313 4607 3327
rect 4733 3313 4747 3327
rect 6673 3313 6687 3327
rect 6833 3313 6847 3327
rect 9213 3313 9227 3327
rect 9313 3313 9327 3327
rect 1033 3292 1047 3306
rect 1093 3293 1107 3307
rect 1593 3293 1607 3307
rect 1653 3293 1667 3307
rect 9673 3293 9687 3307
rect 1913 3253 1927 3267
rect 1953 3253 1967 3267
rect 2973 3252 2987 3266
rect 3053 3253 3067 3267
rect 7573 3253 7587 3267
rect 7673 3253 7687 3267
rect 9673 3253 9687 3267
rect 10033 3293 10047 3307
rect 11093 3293 11107 3307
rect 11153 3293 11167 3307
rect 11293 3273 11307 3287
rect 1913 3232 1927 3246
rect 1973 3233 1987 3247
rect 2593 3233 2607 3247
rect 2653 3231 2667 3245
rect 2753 3233 2767 3247
rect 2893 3233 2907 3247
rect 3093 3233 3107 3247
rect 3153 3233 3167 3247
rect 3673 3231 3687 3245
rect 3733 3233 3747 3247
rect 3953 3233 3967 3247
rect 4093 3233 4107 3247
rect 4833 3233 4847 3247
rect 4933 3233 4947 3247
rect 8313 3233 8327 3247
rect 8413 3233 8427 3247
rect 9053 3233 9067 3247
rect 9113 3233 9127 3247
rect 9153 3233 9167 3247
rect 9293 3233 9307 3247
rect 9393 3233 9407 3247
rect 9553 3233 9567 3247
rect 9773 3233 9787 3247
rect 9813 3233 9827 3247
rect 9973 3233 9987 3247
rect 10013 3232 10027 3246
rect 10053 3233 10067 3247
rect 11233 3233 11247 3247
rect 11293 3233 11307 3247
rect 1593 3213 1607 3227
rect 1633 3213 1647 3227
rect 3833 3213 3847 3227
rect 3573 3193 3587 3207
rect 3713 3193 3727 3207
rect 3913 3212 3927 3226
rect 4033 3213 4047 3227
rect 3473 3173 3487 3187
rect 2273 3153 2287 3167
rect 2333 3153 2347 3167
rect 8953 3153 8967 3167
rect 9073 3153 9087 3167
rect 9493 3153 9507 3167
rect 9553 3153 9567 3167
rect 7813 3113 7827 3127
rect 8053 3113 8067 3127
rect 8853 3113 8867 3127
rect 9813 3113 9827 3127
rect 10073 3113 10087 3127
rect 9953 3093 9967 3107
rect 9993 3092 10007 3106
rect 4133 3073 4147 3087
rect 4193 3073 4207 3087
rect 2293 3053 2307 3067
rect 2373 3052 2387 3066
rect 2493 3053 2507 3067
rect 2633 3053 2647 3067
rect 2753 3053 2767 3067
rect 2893 3053 2907 3067
rect 1793 3032 1807 3046
rect 1913 3033 1927 3047
rect 1053 3013 1067 3027
rect 1113 3013 1127 3027
rect 1973 3013 1987 3027
rect 2153 3033 2167 3047
rect 2333 3033 2347 3047
rect 2393 3033 2407 3047
rect 9753 3033 9767 3047
rect 9793 3033 9807 3047
rect 1553 2993 1567 3007
rect 1673 2993 1687 3007
rect 2193 3013 2207 3027
rect 2253 3013 2267 3027
rect 2333 3012 2347 3026
rect 3673 3013 3687 3027
rect 3713 3013 3727 3027
rect 4973 3013 4987 3027
rect 5113 3013 5127 3027
rect 5413 3013 5427 3027
rect 5453 3013 5467 3027
rect 6093 3013 6107 3027
rect 6233 3013 6247 3027
rect 9773 3013 9787 3027
rect 9833 3013 9847 3027
rect 2253 2992 2267 3006
rect 2393 2993 2407 3007
rect 3953 2993 3967 3007
rect 4013 2993 4027 3007
rect 5233 2993 5247 3007
rect 5353 2993 5367 3007
rect 913 2953 927 2967
rect 993 2953 1007 2967
rect 1073 2953 1087 2967
rect 1213 2953 1227 2967
rect 1813 2953 1827 2967
rect 1913 2953 1927 2967
rect 2153 2953 2167 2967
rect 2293 2953 2307 2967
rect 2353 2953 2367 2967
rect 2493 2953 2507 2967
rect 2613 2953 2627 2967
rect 3213 2953 3227 2967
rect 3273 2953 3287 2967
rect 5213 2953 5227 2967
rect 5253 2953 5267 2967
rect 5913 2953 5927 2967
rect 6033 2953 6047 2967
rect 433 2933 447 2947
rect 593 2933 607 2947
rect 3393 2933 3407 2947
rect 3493 2933 3507 2947
rect 3653 2932 3667 2946
rect 3773 2933 3787 2947
rect 413 2913 427 2927
rect 493 2913 507 2927
rect 1553 2893 1567 2907
rect 1673 2893 1687 2907
rect 2973 2893 2987 2907
rect 3113 2893 3127 2907
rect 3873 2893 3887 2907
rect 4013 2893 4027 2907
rect 4153 2893 4167 2907
rect 4253 2893 4267 2907
rect 4413 2893 4427 2907
rect 4473 2893 4487 2907
rect 4793 2893 4807 2907
rect 4893 2893 4907 2907
rect 5293 2893 5307 2907
rect 5353 2893 5367 2907
rect 4733 2833 4747 2847
rect 4793 2833 4807 2847
rect 4033 2793 4047 2807
rect 4173 2793 4187 2807
rect 6393 2793 6407 2807
rect 6453 2793 6467 2807
rect 8193 2792 8207 2806
rect 8293 2793 8307 2807
rect 10473 2793 10487 2807
rect 10533 2793 10547 2807
rect 4693 2773 4707 2787
rect 4813 2773 4827 2787
rect 9733 2773 9747 2787
rect 9753 2752 9767 2766
rect 11213 2773 11227 2787
rect 6833 2733 6847 2747
rect 6893 2733 6907 2747
rect 11073 2733 11087 2747
rect 113 2713 127 2727
rect 193 2713 207 2727
rect 3613 2713 3627 2727
rect 3693 2713 3707 2727
rect 3833 2713 3847 2727
rect 3953 2713 3967 2727
rect 4733 2713 4747 2727
rect 4833 2713 4847 2727
rect 9713 2713 9727 2727
rect 9833 2713 9847 2727
rect 9993 2713 10007 2727
rect 10093 2712 10107 2726
rect 4273 2633 4287 2647
rect 4353 2633 4367 2647
rect 8553 2593 8567 2607
rect 8753 2593 8767 2607
rect 4833 2573 4847 2587
rect 4913 2573 4927 2587
rect 10653 2573 10667 2587
rect 10993 2573 11007 2587
rect 11073 2573 11087 2587
rect 2133 2553 2147 2567
rect 2213 2553 2227 2567
rect 8313 2553 8327 2567
rect 8433 2553 8447 2567
rect 733 2533 747 2547
rect 793 2533 807 2547
rect 1613 2533 1627 2547
rect 1673 2533 1687 2547
rect 2093 2533 2107 2547
rect 2253 2533 2267 2547
rect 8313 2532 8327 2546
rect 8473 2533 8487 2547
rect 2513 2513 2527 2527
rect 2553 2513 2567 2527
rect 2673 2513 2687 2527
rect 713 2493 727 2507
rect 813 2493 827 2507
rect 1573 2494 1587 2508
rect 1713 2493 1727 2507
rect 1953 2493 1967 2507
rect 1993 2493 2007 2507
rect 4073 2493 4087 2507
rect 4233 2513 4247 2527
rect 4573 2493 4587 2507
rect 4613 2493 4627 2507
rect 8733 2493 8747 2507
rect 8793 2493 8807 2507
rect 8953 2494 8967 2508
rect 9013 2493 9027 2507
rect 9633 2493 9647 2507
rect 9753 2493 9767 2507
rect 4593 2473 4607 2487
rect 4713 2473 4727 2487
rect 7493 2473 7507 2487
rect 7553 2473 7567 2487
rect 8533 2473 8547 2487
rect 8573 2473 8587 2487
rect 11033 2473 11047 2487
rect 11133 2473 11147 2487
rect 1873 2433 1887 2447
rect 1933 2433 1947 2447
rect 2973 2433 2987 2447
rect 3093 2433 3107 2447
rect 8573 2433 8587 2447
rect 8673 2433 8687 2447
rect 10633 2433 10647 2447
rect 10693 2433 10707 2447
rect 1873 2412 1887 2426
rect 2013 2413 2027 2427
rect 4773 2413 4787 2427
rect 4893 2413 4907 2427
rect 4873 2393 4887 2407
rect 4933 2393 4947 2407
rect 2093 2373 2107 2387
rect 2213 2373 2227 2387
rect 5213 2373 5227 2387
rect 5333 2373 5347 2387
rect 7933 2313 7947 2327
rect 7993 2313 8007 2327
rect 1093 2293 1107 2307
rect 1253 2293 1267 2307
rect 2533 2293 2547 2307
rect 2613 2293 2627 2307
rect 5033 2293 5047 2307
rect 5093 2293 5107 2307
rect 5773 2293 5787 2307
rect 5853 2293 5867 2307
rect 7873 2293 7887 2307
rect 7993 2292 8007 2306
rect 9553 2293 9567 2307
rect 9613 2293 9627 2307
rect 10873 2293 10887 2307
rect 10913 2292 10927 2306
rect 253 2273 267 2287
rect 393 2273 407 2287
rect 433 2273 447 2287
rect 553 2273 567 2287
rect 5273 2273 5287 2287
rect 5333 2272 5347 2286
rect 6473 2273 6487 2287
rect 6533 2274 6547 2288
rect 10193 2273 10207 2287
rect 10293 2273 10307 2287
rect 10713 2273 10727 2287
rect 10813 2273 10827 2287
rect 1813 2253 1827 2267
rect 4573 2253 4587 2267
rect 4693 2253 4707 2267
rect 6233 2253 6247 2267
rect 6333 2253 6347 2267
rect 7993 2253 8007 2267
rect 8033 2253 8047 2267
rect 9553 2253 9567 2267
rect 9713 2253 9727 2267
rect 753 2192 767 2206
rect 793 2193 807 2207
rect 853 2193 867 2207
rect 1013 2193 1027 2207
rect 1793 2193 1807 2207
rect 2033 2213 2047 2227
rect 2113 2213 2127 2227
rect 3053 2213 3067 2227
rect 8873 2213 8887 2227
rect 8993 2213 9007 2227
rect 2253 2193 2267 2207
rect 2453 2193 2467 2207
rect 2933 2193 2947 2207
rect 3033 2193 3047 2207
rect 2953 2173 2967 2187
rect 3933 2193 3947 2207
rect 4013 2193 4027 2207
rect 5213 2193 5227 2207
rect 5313 2193 5327 2207
rect 5453 2193 5467 2207
rect 5513 2193 5527 2207
rect 5633 2193 5647 2207
rect 8833 2193 8847 2207
rect 9033 2193 9047 2207
rect 9973 2193 9987 2207
rect 10013 2193 10027 2207
rect 10433 2193 10447 2207
rect 10513 2193 10527 2207
rect 10713 2193 10727 2207
rect 10813 2193 10827 2207
rect 10853 2193 10867 2207
rect 10973 2193 10987 2207
rect 9993 2173 10007 2187
rect 10033 2173 10047 2187
rect 1833 2153 1847 2167
rect 1933 2153 1947 2167
rect 2733 2153 2747 2167
rect 2853 2153 2867 2167
rect 953 2133 967 2147
rect 993 2133 1007 2147
rect 5233 2113 5247 2127
rect 5293 2113 5307 2127
rect 5633 2073 5647 2087
rect 6893 2073 6907 2087
rect 9213 2073 9227 2087
rect 3133 2053 3147 2067
rect 3273 2053 3287 2067
rect 6553 2033 6567 2047
rect 6673 2033 6687 2047
rect 1533 2013 1547 2027
rect 1693 2013 1707 2027
rect 11013 1993 11027 2007
rect 11173 1993 11187 2007
rect 1393 1973 1407 1987
rect 2553 1973 2567 1987
rect 2633 1973 2647 1987
rect 3353 1973 3367 1987
rect 3393 1973 3407 1987
rect 3493 1973 3507 1987
rect 1113 1953 1127 1967
rect 1233 1953 1247 1967
rect 1333 1953 1347 1967
rect 3573 1972 3587 1986
rect 7273 1973 7287 1987
rect 7373 1973 7387 1987
rect 8793 1973 8807 1987
rect 8853 1973 8867 1987
rect 9753 1973 9767 1987
rect 9793 1974 9807 1988
rect 10293 1973 10307 1987
rect 10333 1972 10347 1986
rect 3613 1953 3627 1967
rect 3733 1953 3747 1967
rect 4073 1953 4087 1967
rect 4193 1953 4207 1967
rect 4733 1953 4747 1967
rect 4813 1953 4827 1967
rect 6133 1953 6147 1967
rect 6233 1953 6247 1967
rect 9653 1953 9667 1967
rect 9733 1953 9747 1967
rect 9993 1953 10007 1967
rect 10553 1953 10567 1967
rect 3133 1913 3147 1927
rect 3253 1913 3267 1927
rect 8973 1913 8987 1927
rect 9073 1913 9087 1927
rect 9653 1913 9667 1927
rect 9713 1913 9727 1927
rect 9853 1913 9867 1927
rect 10553 1913 10567 1927
rect 5633 1873 5647 1887
rect 5753 1873 5767 1887
rect 5893 1853 5907 1867
rect 5933 1853 5947 1867
rect 7433 1853 7447 1867
rect 7573 1853 7587 1867
rect 3293 1753 3307 1767
rect 3453 1753 3467 1767
rect 9333 1753 9347 1767
rect 9913 1753 9927 1767
rect 10073 1753 10087 1767
rect 6953 1733 6967 1747
rect 7073 1733 7087 1747
rect 9193 1733 9207 1747
rect 10333 1732 10347 1746
rect 2013 1693 2027 1707
rect 2093 1693 2107 1707
rect 9193 1693 9207 1707
rect 9233 1693 9247 1707
rect 9513 1693 9527 1707
rect 9573 1693 9587 1707
rect 1093 1673 1107 1687
rect 1233 1673 1247 1687
rect 2053 1673 2067 1687
rect 2153 1673 2167 1687
rect 2653 1673 2667 1687
rect 2793 1671 2807 1685
rect 3073 1673 3087 1687
rect 3193 1673 3207 1687
rect 5753 1673 5767 1687
rect 5973 1673 5987 1687
rect 7013 1673 7027 1687
rect 7093 1673 7107 1687
rect 10113 1673 10127 1687
rect 10273 1673 10287 1687
rect 10313 1673 10327 1687
rect 1053 1633 1067 1647
rect 1213 1633 1227 1647
rect 1273 1633 1287 1647
rect 1333 1633 1347 1647
rect 3793 1593 3807 1607
rect 3913 1593 3927 1607
rect 4833 1552 4847 1566
rect 6393 1553 6407 1567
rect 7713 1553 7727 1567
rect 9113 1533 9127 1547
rect 9233 1533 9247 1547
rect 4933 1513 4947 1527
rect 8433 1513 8447 1527
rect 8473 1513 8487 1527
rect 4833 1493 4847 1507
rect 8833 1493 8847 1507
rect 8953 1493 8967 1507
rect 3773 1473 3787 1487
rect 3933 1473 3947 1487
rect 3273 1453 3287 1467
rect 3393 1453 3407 1467
rect 5033 1454 5047 1468
rect 5093 1453 5107 1467
rect 5933 1453 5947 1467
rect 5993 1453 6007 1467
rect 8033 1453 8047 1467
rect 8073 1454 8087 1468
rect 9073 1453 9087 1467
rect 9213 1453 9227 1467
rect 9693 1454 9707 1468
rect 9833 1453 9847 1467
rect 10173 1453 10187 1467
rect 10333 1453 10347 1467
rect 10833 1453 10847 1467
rect 10953 1453 10967 1467
rect 8993 1393 9007 1407
rect 10653 1393 10667 1407
rect 10733 1393 10747 1407
rect 1813 1373 1827 1387
rect 1853 1373 1867 1387
rect 5053 1373 5067 1387
rect 5093 1373 5107 1387
rect 8853 1373 8867 1387
rect 10173 1373 10187 1387
rect 10333 1373 10347 1387
rect 1293 1353 1307 1367
rect 1453 1353 1467 1367
rect 7173 1353 7187 1367
rect 7053 1333 7067 1347
rect 1993 1273 2007 1287
rect 2133 1273 2147 1287
rect 10373 1273 10387 1287
rect 10473 1273 10487 1287
rect 3633 1233 3647 1247
rect 3793 1234 3807 1248
rect 3833 1233 3847 1247
rect 3953 1233 3967 1247
rect 6153 1233 6167 1247
rect 6273 1233 6287 1247
rect 8793 1233 8807 1247
rect 8873 1233 8887 1247
rect 9013 1233 9027 1247
rect 9113 1233 9127 1247
rect 4753 1213 4767 1227
rect 4873 1213 4887 1227
rect 10133 1213 10147 1227
rect 10213 1213 10227 1227
rect 3693 1173 3707 1187
rect 11073 1173 11087 1187
rect 11133 1173 11147 1187
rect 2333 1153 2347 1167
rect 2373 1153 2387 1167
rect 3613 1153 3627 1167
rect 6133 1153 6147 1167
rect 6233 1153 6247 1167
rect 8393 1153 8407 1167
rect 8473 1153 8487 1167
rect 8613 1153 8627 1167
rect 8713 1153 8727 1167
rect 11053 1152 11067 1166
rect 11213 1153 11227 1167
rect 10093 1133 10107 1147
rect 10253 1133 10267 1147
rect 5733 1113 5747 1127
rect 5853 1113 5867 1127
rect 9233 1113 9247 1127
rect 9373 1113 9387 1127
rect 3373 953 3387 967
rect 3533 953 3547 967
rect 8893 953 8907 967
rect 9013 953 9027 967
rect 1473 933 1487 947
rect 1573 933 1587 947
rect 2673 933 2687 947
rect 2813 934 2827 948
rect 3313 933 3327 947
rect 3413 933 3427 947
rect 3493 933 3507 947
rect 4213 932 4227 946
rect 4313 933 4327 947
rect 4593 933 4607 947
rect 4633 933 4647 947
rect 7253 933 7267 947
rect 7313 933 7327 947
rect 10973 933 10987 947
rect 11053 933 11067 947
rect 4293 913 4307 927
rect 4413 913 4427 927
rect 10993 873 11007 887
rect 11033 873 11047 887
rect 4993 713 5007 727
rect 5533 713 5547 727
rect 5613 713 5627 727
rect 6473 713 6487 727
rect 6613 713 6627 727
rect 7853 713 7867 727
rect 7953 713 7967 727
rect 9073 713 9087 727
rect 9213 713 9227 727
rect 9393 713 9407 727
rect 9433 713 9447 727
rect 9473 713 9487 727
rect 9653 713 9667 727
rect 4933 693 4947 707
rect 8433 673 8447 687
rect 8493 673 8507 687
rect 833 633 847 647
rect 913 633 927 647
rect 4353 633 4367 647
rect 4413 633 4427 647
rect 4853 633 4867 647
rect 4953 633 4967 647
rect 5013 633 5027 647
rect 6213 633 6227 647
rect 6393 633 6407 647
rect 7853 633 7867 647
rect 7933 633 7947 647
rect 5773 613 5787 627
rect 5933 613 5947 627
rect 10633 593 10647 607
rect 10733 593 10747 607
rect 7933 553 7947 567
rect 8073 553 8087 567
rect 1133 513 1147 527
rect 1813 513 1827 527
rect 2293 513 2307 527
rect 10533 513 10547 527
rect 2193 413 2207 427
rect 2393 413 2407 427
rect 2633 413 2647 427
rect 2753 413 2767 427
rect 3433 413 3447 427
rect 3673 413 3687 427
rect 3733 413 3747 427
rect 3913 413 3927 427
rect 8453 413 8467 427
rect 8573 413 8587 427
rect 10293 413 10307 427
rect 10353 413 10367 427
rect 213 393 227 407
rect 333 393 347 407
rect 10493 393 10507 407
rect 10533 393 10547 407
rect 6193 353 6207 367
rect 6233 353 6247 367
rect 453 333 467 347
rect 573 333 587 347
rect 3233 333 3247 347
rect 3313 333 3327 347
rect 4173 333 4187 347
rect 4213 333 4227 347
rect 5513 333 5527 347
rect 5553 333 5567 347
rect 9993 333 10007 347
rect 10073 332 10087 346
rect 10193 293 10207 307
rect 10273 293 10287 307
rect 8113 193 8127 207
rect 8293 193 8307 207
rect 8333 133 8347 147
rect 8473 133 8487 147
rect 9233 133 9247 147
rect 9333 133 9347 147
rect 2713 113 2727 127
rect 2833 113 2847 127
rect 9233 112 9247 126
rect 9333 112 9347 126
rect 9693 113 9707 127
rect 9833 113 9847 127
<< metal2 >>
rect 16 10907 23 11094
rect 136 11056 153 11063
rect 16 5807 23 10893
rect 36 10687 43 10783
rect 96 10780 103 10783
rect 93 10767 107 10780
rect 136 10588 143 11056
rect 336 10947 343 11073
rect 376 11057 383 11243
rect 380 11056 383 11057
rect 397 11028 404 11104
rect 1353 11100 1367 11113
rect 1356 11096 1363 11100
rect 376 11021 404 11028
rect 376 10687 383 11021
rect 456 10827 463 11043
rect 616 11007 623 11083
rect 853 11080 867 11093
rect 856 11076 863 11080
rect 176 10576 183 10673
rect 136 9847 143 10574
rect 256 10246 263 10273
rect 196 10240 203 10243
rect 193 10227 207 10240
rect 216 10056 223 10093
rect 256 10068 263 10232
rect 196 9867 203 10023
rect 236 9756 243 9793
rect 256 9767 263 10054
rect 136 9548 143 9754
rect 76 5583 83 5993
rect 96 5747 103 9433
rect 116 8987 123 9213
rect 136 9027 143 9534
rect 256 9503 263 9534
rect 196 9487 203 9503
rect 236 9496 263 9503
rect 196 9476 213 9487
rect 200 9473 213 9476
rect 173 9240 187 9253
rect 176 9236 183 9240
rect 216 9167 223 9203
rect 213 9000 227 9013
rect 236 9007 243 9496
rect 276 9023 283 10633
rect 396 10607 403 10783
rect 416 10647 423 10774
rect 296 9567 303 9853
rect 316 9707 323 10113
rect 336 9867 343 10593
rect 416 10576 423 10633
rect 476 10546 483 10673
rect 536 10407 543 10783
rect 556 10687 563 10774
rect 576 10546 583 10613
rect 636 10576 643 10673
rect 796 10623 803 10993
rect 836 10767 843 10783
rect 836 10667 843 10753
rect 776 10616 803 10623
rect 676 10576 723 10583
rect 716 10547 723 10576
rect 656 10483 663 10543
rect 656 10476 683 10483
rect 647 10393 653 10407
rect 396 10276 403 10313
rect 636 10276 643 10313
rect 356 10023 363 10213
rect 416 10068 423 10243
rect 456 10056 463 10113
rect 496 10107 503 10274
rect 676 10207 683 10476
rect 716 10247 723 10274
rect 496 10026 503 10093
rect 356 10016 403 10023
rect 356 9727 363 9773
rect 376 9547 383 10016
rect 516 10007 523 10054
rect 416 9756 423 9833
rect 453 9760 467 9773
rect 456 9756 463 9760
rect 436 9720 443 9723
rect 433 9707 447 9720
rect 393 9540 407 9553
rect 396 9536 403 9540
rect 416 9500 423 9503
rect 336 9206 343 9493
rect 413 9487 427 9500
rect 496 9248 503 9533
rect 516 9506 523 9833
rect 436 9107 443 9203
rect 256 9016 283 9023
rect 216 8996 223 9000
rect 116 7827 123 8433
rect 136 8087 143 8973
rect 176 8767 183 8972
rect 216 8727 223 8913
rect 196 8587 203 8683
rect 176 8576 193 8583
rect 176 8496 183 8576
rect 216 8527 223 8713
rect 216 8496 223 8513
rect 236 8507 243 8953
rect 196 8196 203 8463
rect 236 8196 243 8333
rect 256 8203 263 9016
rect 316 9006 323 9093
rect 296 8647 303 8953
rect 556 8847 563 9873
rect 576 9807 583 10054
rect 636 10020 643 10023
rect 633 10007 647 10020
rect 776 9827 783 10616
rect 856 10576 863 10613
rect 896 10587 903 10783
rect 916 10667 923 11074
rect 1056 11060 1063 11063
rect 1053 11047 1067 11060
rect 1036 10707 1043 10814
rect 1056 10787 1063 10913
rect 1096 10796 1103 10993
rect 1216 10887 1223 11093
rect 1396 11067 1403 11243
rect 1116 10760 1123 10763
rect 1113 10747 1127 10760
rect 1216 10747 1223 10873
rect 1516 10786 1523 11093
rect 1536 11060 1543 11063
rect 1533 11047 1547 11060
rect 1536 10867 1543 11033
rect 1736 11007 1743 11243
rect 1796 11096 1803 11133
rect 1833 11100 1847 11113
rect 1836 11096 1843 11100
rect 1816 11007 1823 11063
rect 1736 10907 1743 10953
rect 956 10556 983 10563
rect 836 10347 843 10532
rect 876 10447 883 10532
rect 916 10487 923 10523
rect 816 10056 823 10113
rect 836 9887 843 10023
rect 576 9627 583 9793
rect 916 9787 923 10473
rect 976 10407 983 10556
rect 1076 10367 1083 10563
rect 1216 10487 1223 10693
rect 1496 10667 1503 10783
rect 1736 10763 1743 10893
rect 1793 10800 1807 10813
rect 1796 10796 1803 10800
rect 1736 10756 1763 10763
rect 1276 10563 1283 10653
rect 1256 10556 1283 10563
rect 1316 10556 1343 10563
rect 1416 10556 1443 10563
rect 1076 10276 1083 10313
rect 1196 10247 1203 10274
rect 1096 10223 1103 10232
rect 1076 10216 1103 10223
rect 1036 10023 1043 10093
rect 1076 10087 1083 10216
rect 1096 10056 1103 10113
rect 1116 10107 1123 10213
rect 1216 10187 1223 10433
rect 1236 10127 1243 10413
rect 1176 10096 1193 10103
rect 1156 10056 1163 10093
rect 1176 10068 1183 10096
rect 1036 10016 1063 10023
rect 1116 10020 1123 10023
rect 1113 10007 1127 10020
rect 1196 10007 1203 10093
rect 576 8996 583 9353
rect 596 9147 603 9774
rect 636 9756 663 9763
rect 636 9727 643 9756
rect 907 9763 920 9767
rect 907 9753 923 9763
rect 696 9720 703 9723
rect 693 9707 707 9720
rect 656 9536 663 9693
rect 636 9447 643 9503
rect 676 9407 683 9503
rect 776 9407 783 9534
rect 796 9363 803 9743
rect 916 9736 923 9753
rect 1096 9727 1103 9743
rect 876 9536 883 9613
rect 856 9467 863 9503
rect 956 9447 963 9633
rect 1096 9587 1103 9713
rect 796 9356 813 9363
rect 827 9353 833 9367
rect 856 9236 863 9273
rect 656 8967 663 9133
rect 676 9127 683 9203
rect 336 8547 343 8753
rect 453 8740 467 8753
rect 456 8736 463 8740
rect 416 8607 423 8683
rect 256 8196 283 8203
rect 176 8067 183 8163
rect 216 7976 223 8033
rect 116 5983 123 7813
rect 276 7787 283 8196
rect 296 8166 303 8513
rect 356 8327 363 8593
rect 456 8496 463 8533
rect 396 8443 403 8463
rect 436 8460 443 8463
rect 433 8447 447 8460
rect 396 8436 423 8443
rect 196 7676 203 7733
rect 256 7646 263 7673
rect 176 7468 183 7643
rect 176 6967 183 7123
rect 136 6648 143 6953
rect 233 6920 247 6933
rect 256 6927 263 7454
rect 276 7168 283 7273
rect 276 6967 283 7154
rect 236 6916 243 6920
rect 176 6663 183 6903
rect 216 6787 223 6893
rect 176 6656 203 6663
rect 196 6636 203 6656
rect 176 6567 183 6603
rect 276 6563 283 6953
rect 296 6916 303 6993
rect 316 6927 323 8313
rect 373 8287 387 8293
rect 416 8287 423 8436
rect 496 8307 503 8703
rect 416 8160 423 8163
rect 413 8147 427 8160
rect 396 7976 403 8073
rect 336 7427 343 7632
rect 356 7607 363 7974
rect 516 7967 523 8833
rect 616 8767 623 8952
rect 736 8927 743 9014
rect 756 8708 763 9053
rect 776 8747 783 9233
rect 876 9167 883 9203
rect 876 9023 883 9153
rect 856 9016 883 9023
rect 796 8647 803 8703
rect 636 8496 643 8533
rect 676 8496 683 8573
rect 776 8487 783 8533
rect 656 8427 663 8463
rect 696 8327 703 8463
rect 536 7956 543 8293
rect 556 8047 563 8152
rect 636 8067 643 8163
rect 676 8160 683 8163
rect 673 8147 687 8160
rect 416 7767 423 7932
rect 416 7703 423 7753
rect 456 7747 463 7943
rect 496 7920 503 7923
rect 493 7907 507 7920
rect 396 7696 423 7703
rect 396 7676 403 7696
rect 427 7493 433 7507
rect 396 7456 403 7493
rect 456 7468 463 7643
rect 476 7367 483 7593
rect 496 7426 503 7753
rect 556 7607 563 8033
rect 796 7927 803 8633
rect 816 8427 823 8733
rect 856 8700 863 8703
rect 853 8687 867 8700
rect 876 8496 883 8613
rect 976 8447 983 9453
rect 1016 9347 1023 9393
rect 996 8607 1003 9313
rect 1016 9206 1023 9333
rect 1076 9243 1083 9503
rect 1116 9487 1123 9813
rect 1136 9506 1143 9533
rect 1156 9407 1163 9743
rect 1056 9236 1083 9243
rect 1116 9236 1123 9273
rect 1056 9206 1063 9236
rect 1136 9107 1143 9203
rect 1096 9016 1103 9053
rect 1036 8947 1043 8983
rect 1136 8947 1143 9033
rect 1036 8727 1043 8833
rect 1076 8823 1083 8933
rect 1056 8816 1083 8823
rect 1056 8716 1063 8816
rect 1076 8567 1083 8672
rect 996 8467 1003 8494
rect 1156 8467 1163 9193
rect 1176 8647 1183 9573
rect 1196 9443 1203 9972
rect 1216 9767 1223 9993
rect 1216 9467 1223 9753
rect 1236 9687 1243 10073
rect 1276 9727 1283 10556
rect 1336 10447 1343 10556
rect 1376 10487 1383 10523
rect 1436 10407 1443 10556
rect 1396 10236 1423 10243
rect 1296 9987 1303 10093
rect 1356 10056 1363 10172
rect 1416 10147 1423 10236
rect 1476 10207 1483 10293
rect 1376 9788 1383 10023
rect 1316 9726 1323 9773
rect 1456 9727 1463 9754
rect 1296 9536 1303 9653
rect 1356 9627 1363 9712
rect 1396 9687 1403 9723
rect 1196 9436 1223 9443
rect 1216 8447 1223 9436
rect 1276 9427 1283 9503
rect 1313 9487 1327 9492
rect 1236 8847 1243 9413
rect 1276 9207 1283 9253
rect 1313 9240 1327 9253
rect 1356 9248 1363 9473
rect 1316 9236 1323 9240
rect 1416 9206 1423 9553
rect 1336 9127 1343 9203
rect 1273 9020 1287 9033
rect 1276 9016 1283 9020
rect 1316 9016 1323 9093
rect 1336 9067 1343 9113
rect 1413 9027 1427 9033
rect 1296 8787 1303 8983
rect 1336 8947 1343 8983
rect 1316 8748 1323 8853
rect 1376 8787 1383 8873
rect 1436 8867 1443 9254
rect 1456 9027 1463 9573
rect 1476 9567 1483 10013
rect 1516 9647 1523 10213
rect 1536 10207 1543 10353
rect 1593 10280 1607 10293
rect 1596 10276 1603 10280
rect 1676 10287 1683 10753
rect 1696 10566 1703 10613
rect 1716 10556 1723 10653
rect 1776 10556 1803 10563
rect 1796 10507 1803 10556
rect 1776 10307 1783 10433
rect 1876 10347 1883 11113
rect 1576 10240 1583 10243
rect 1573 10227 1587 10240
rect 1616 10207 1623 10243
rect 1556 10056 1563 10173
rect 1676 9763 1683 10273
rect 1776 10187 1783 10293
rect 1813 10280 1827 10293
rect 1876 10283 1883 10333
rect 1816 10276 1823 10280
rect 1856 10276 1883 10283
rect 1916 10246 1923 11133
rect 1996 11063 2003 11243
rect 1996 11056 2023 11063
rect 1936 10583 1943 10853
rect 1976 10796 1983 10853
rect 1996 10647 2003 10763
rect 1936 10576 1953 10583
rect 1996 10576 2003 10612
rect 2036 10576 2043 10613
rect 2076 10546 2083 10633
rect 2056 10167 2063 10232
rect 1796 10056 1803 10133
rect 1716 10027 1723 10054
rect 1856 10047 1863 10093
rect 1993 10068 2007 10073
rect 1776 10020 1783 10023
rect 1816 10020 1823 10023
rect 1716 9867 1723 10013
rect 1773 10007 1787 10020
rect 1813 10007 1827 10020
rect 1656 9756 1703 9763
rect 1636 9667 1643 9723
rect 1556 9536 1563 9573
rect 1636 9547 1643 9653
rect 1696 9506 1703 9756
rect 1756 9607 1763 9754
rect 1736 9536 1743 9573
rect 1776 9536 1783 9712
rect 1496 9500 1503 9503
rect 1493 9487 1507 9500
rect 1536 9467 1543 9503
rect 1756 9467 1763 9503
rect 1876 9487 1883 9933
rect 1476 9187 1483 9393
rect 1516 9227 1523 9353
rect 1556 9236 1563 9333
rect 1916 9327 1923 10053
rect 2056 10047 2063 10093
rect 1936 9726 1943 9753
rect 1976 9536 1983 9993
rect 2036 9807 2043 10023
rect 2096 9727 2103 11094
rect 2056 9687 2063 9723
rect 1996 9347 2003 9503
rect 2036 9287 2043 9503
rect 1916 9228 1923 9273
rect 1576 9187 1583 9203
rect 1576 9147 1583 9173
rect 1513 9020 1527 9033
rect 1516 9016 1523 9020
rect 1556 9016 1563 9053
rect 1233 8720 1247 8734
rect 1236 8716 1243 8720
rect 1276 8680 1283 8683
rect 1273 8667 1287 8680
rect 1376 8603 1383 8773
rect 1476 8696 1483 8733
rect 1676 8703 1683 9173
rect 1696 9016 1743 9023
rect 1776 9016 1783 9073
rect 1696 8747 1703 9016
rect 1796 8867 1803 8983
rect 1656 8696 1683 8703
rect 1376 8596 1403 8603
rect 1356 8496 1363 8573
rect 816 8247 823 8413
rect 1296 8407 1303 8463
rect 1336 8447 1343 8463
rect 1396 8447 1403 8596
rect 1436 8487 1443 8533
rect 1536 8496 1543 8573
rect 1336 8367 1343 8433
rect 876 8107 883 8163
rect 856 7987 863 8073
rect 836 7956 863 7963
rect 896 7956 903 8093
rect 936 7963 943 8193
rect 956 8127 963 8333
rect 1096 8196 1103 8313
rect 1296 8208 1303 8353
rect 1333 8200 1347 8213
rect 1336 8196 1343 8200
rect 1116 8127 1123 8163
rect 1276 8127 1283 8163
rect 1256 8007 1263 8113
rect 916 7956 943 7963
rect 996 7956 1023 7963
rect 856 7927 863 7956
rect 896 7767 903 7813
rect 916 7807 923 7956
rect 956 7907 963 7923
rect 636 7676 643 7753
rect 676 7676 683 7733
rect 656 7567 663 7643
rect 567 7493 573 7507
rect 336 6907 343 7313
rect 376 7156 383 7213
rect 416 7067 423 7123
rect 496 7047 503 7412
rect 596 7207 603 7393
rect 656 7287 663 7423
rect 656 7156 663 7193
rect 687 7154 693 7167
rect 680 7153 693 7154
rect 596 6967 603 7123
rect 476 6920 483 6923
rect 473 6907 487 6920
rect 576 6916 603 6923
rect 267 6556 283 6563
rect 213 6420 227 6433
rect 216 6416 223 6420
rect 256 6387 263 6553
rect 316 6447 323 6873
rect 336 6627 343 6893
rect 176 6327 183 6383
rect 236 6083 243 6253
rect 316 6227 323 6433
rect 336 6327 343 6453
rect 356 6128 363 6473
rect 376 6428 383 6633
rect 496 6607 503 6773
rect 576 6767 583 6916
rect 636 6747 643 6883
rect 676 6663 683 7033
rect 756 7027 763 7153
rect 696 6867 703 6993
rect 776 6948 783 7513
rect 816 7456 823 7493
rect 856 7468 863 7632
rect 896 7347 903 7454
rect 956 7427 963 7893
rect 1016 7807 1023 7956
rect 1296 7956 1323 7963
rect 1356 7956 1363 8073
rect 1316 7927 1323 7956
rect 1316 7847 1323 7913
rect 976 7647 983 7674
rect 976 7387 983 7553
rect 827 7163 840 7167
rect 827 7156 843 7163
rect 827 7153 840 7156
rect 796 7127 803 7153
rect 896 7140 903 7143
rect 893 7127 907 7140
rect 796 7007 803 7053
rect 676 6656 703 6663
rect 696 6648 703 6656
rect 416 6416 423 6473
rect 436 6380 443 6383
rect 433 6367 447 6380
rect 436 6116 443 6153
rect 216 6076 243 6083
rect 416 5987 423 6083
rect 456 6080 463 6083
rect 453 6067 467 6080
rect 516 6067 523 6372
rect 536 6367 543 6633
rect 776 6623 783 6934
rect 956 6867 963 7143
rect 976 6907 983 7033
rect 996 6867 1003 7693
rect 1073 7680 1087 7693
rect 1076 7676 1083 7680
rect 1276 7676 1283 7713
rect 1036 7487 1043 7513
rect 1056 7507 1063 7643
rect 1096 7587 1103 7643
rect 1296 7607 1303 7643
rect 1376 7587 1383 8433
rect 1036 7456 1043 7473
rect 1236 7456 1243 7493
rect 1056 7367 1063 7423
rect 1116 7407 1123 7454
rect 1256 7420 1263 7423
rect 1253 7407 1267 7420
rect 1133 7140 1147 7153
rect 1136 7136 1143 7140
rect 1236 7047 1243 7213
rect 1296 7188 1303 7413
rect 1356 7287 1363 7533
rect 1396 7503 1403 8412
rect 1456 8367 1463 8494
rect 1616 8407 1623 8493
rect 1636 8427 1643 8653
rect 1656 8647 1663 8696
rect 1716 8667 1723 8703
rect 1776 8496 1783 8733
rect 1796 8587 1803 8853
rect 1416 7887 1423 8194
rect 1436 7688 1443 8233
rect 1456 7927 1463 8353
rect 1796 8287 1803 8463
rect 1836 8407 1843 8933
rect 1856 8623 1863 9014
rect 1876 8647 1883 9033
rect 1916 8947 1923 9214
rect 1956 9187 1963 9223
rect 2016 9127 2023 9223
rect 2056 9047 2063 9133
rect 1993 9020 2007 9033
rect 1996 9016 2003 9020
rect 2076 8987 2083 9453
rect 1976 8947 1983 8983
rect 1916 8716 1923 8853
rect 1936 8680 1943 8683
rect 1933 8667 1947 8680
rect 1856 8616 1883 8623
rect 1473 8227 1487 8233
rect 1476 8127 1483 8192
rect 1656 8163 1663 8273
rect 1713 8200 1727 8213
rect 1716 8196 1723 8200
rect 1476 7988 1483 8113
rect 1536 8087 1543 8163
rect 1656 8156 1703 8163
rect 1736 8127 1743 8163
rect 1796 8147 1803 8194
rect 1516 7676 1523 8033
rect 1656 8007 1663 8113
rect 1593 7980 1607 7993
rect 1596 7976 1603 7980
rect 1576 7927 1583 7943
rect 1556 7676 1563 7753
rect 1576 7707 1583 7913
rect 1436 7547 1443 7674
rect 1536 7507 1543 7643
rect 1616 7643 1623 7693
rect 1596 7636 1623 7643
rect 1576 7527 1583 7632
rect 1376 7496 1403 7503
rect 1376 7307 1383 7496
rect 1456 7476 1513 7483
rect 1316 7247 1323 7273
rect 1033 6940 1047 6953
rect 1256 6948 1263 7073
rect 1036 6936 1043 6940
rect 1276 6936 1283 7033
rect 1316 6936 1323 7053
rect 836 6627 843 6853
rect 1016 6767 1023 6893
rect 1056 6883 1063 6903
rect 1096 6900 1103 6903
rect 1296 6900 1303 6903
rect 1093 6887 1107 6900
rect 1056 6876 1083 6883
rect 656 6583 663 6592
rect 656 6576 683 6583
rect 656 6467 663 6533
rect 676 6503 683 6576
rect 736 6527 743 6623
rect 756 6616 783 6623
rect 676 6496 703 6503
rect 656 6416 663 6453
rect 576 6327 583 6414
rect 576 6267 583 6313
rect 636 6116 643 6153
rect 696 6147 703 6496
rect 116 5976 143 5983
rect 36 5487 43 5583
rect 76 5576 103 5583
rect 136 4987 143 5976
rect 216 5896 223 5933
rect 293 5880 307 5893
rect 316 5886 323 5973
rect 296 5876 303 5880
rect 276 5576 283 5613
rect 176 5376 183 5473
rect 376 5383 383 5733
rect 416 5623 423 5833
rect 556 5727 563 5893
rect 596 5876 603 5993
rect 656 5888 663 6083
rect 416 5616 443 5623
rect 556 5587 563 5713
rect 367 5376 383 5383
rect 416 5376 423 5533
rect 596 5388 603 5793
rect 633 5600 647 5613
rect 636 5596 643 5600
rect 656 5560 663 5563
rect 653 5547 667 5560
rect 676 5388 683 5413
rect 156 5340 163 5343
rect 153 5327 167 5340
rect 196 5076 203 5173
rect 253 5080 267 5093
rect 256 5076 263 5080
rect 236 5023 243 5043
rect 216 5016 243 5023
rect 176 4856 183 4933
rect 216 4856 223 5016
rect 296 4826 303 4873
rect 236 4687 243 4823
rect 193 4560 207 4573
rect 196 4556 203 4560
rect 76 1287 83 3772
rect 136 3487 143 4512
rect 216 4427 223 4523
rect 213 4363 227 4373
rect 196 4360 227 4363
rect 196 4356 223 4360
rect 196 4336 203 4356
rect 156 4247 163 4303
rect 216 4267 223 4303
rect 196 4036 203 4233
rect 176 3983 183 4003
rect 176 3976 203 3983
rect 196 3816 203 3976
rect 216 3947 223 4003
rect 276 3787 283 4633
rect 176 3727 183 3783
rect 236 3516 243 3593
rect 216 3387 223 3483
rect 256 3267 263 3473
rect 276 3308 283 3633
rect 176 2996 183 3233
rect 196 2907 203 2963
rect 116 2447 123 2713
rect 136 2227 143 2833
rect 236 2807 243 3113
rect 173 2780 187 2793
rect 176 2776 183 2780
rect 196 2740 203 2743
rect 193 2727 207 2740
rect 196 2307 203 2432
rect 173 2260 187 2273
rect 253 2268 267 2273
rect 176 2256 183 2260
rect 256 2087 263 2254
rect 276 2107 283 2633
rect 196 1956 203 2073
rect 196 1736 203 1773
rect 176 1700 183 1703
rect 173 1687 187 1700
rect 256 1687 263 1912
rect 296 1787 303 4812
rect 316 2647 323 4713
rect 336 3987 343 5093
rect 356 4787 363 5374
rect 436 5307 443 5343
rect 456 4856 463 5113
rect 513 5088 527 5093
rect 496 4987 503 5043
rect 576 4826 583 4893
rect 416 4607 423 4773
rect 596 4727 603 5374
rect 636 5340 643 5343
rect 633 5327 647 5340
rect 696 5327 703 6053
rect 616 4967 623 5074
rect 636 4868 643 5273
rect 373 4560 387 4573
rect 376 4556 383 4560
rect 416 4556 423 4593
rect 653 4560 667 4573
rect 696 4567 703 5133
rect 716 5087 723 5613
rect 736 5147 743 6193
rect 756 5807 763 6616
rect 976 6616 983 6753
rect 776 5608 783 6513
rect 796 6467 803 6612
rect 796 6007 803 6453
rect 856 6416 863 6513
rect 836 6207 843 6383
rect 976 6207 983 6493
rect 996 6307 1003 6513
rect 1076 6507 1083 6876
rect 1293 6887 1307 6900
rect 1136 6668 1143 6733
rect 1096 6443 1103 6533
rect 1176 6527 1183 6853
rect 1033 6420 1047 6433
rect 1076 6436 1103 6443
rect 1036 6416 1043 6420
rect 1076 6416 1083 6436
rect 1096 6327 1103 6383
rect 1196 6366 1203 6653
rect 1276 6627 1283 6753
rect 1356 6663 1363 7174
rect 1376 7147 1383 7253
rect 1396 7126 1403 7473
rect 1456 7456 1463 7476
rect 1436 7420 1443 7423
rect 1433 7407 1447 7420
rect 1476 7387 1483 7423
rect 1347 6656 1363 6663
rect 1333 6640 1347 6654
rect 1336 6636 1343 6640
rect 1416 6606 1423 7293
rect 1436 6887 1443 7273
rect 1516 7207 1523 7373
rect 1536 7267 1543 7493
rect 1516 7156 1523 7193
rect 1556 7156 1563 7233
rect 1536 7087 1543 7123
rect 1456 6947 1463 6993
rect 1496 6936 1503 7013
rect 1276 6363 1283 6393
rect 1276 6356 1303 6363
rect 816 5987 823 6153
rect 833 6120 847 6133
rect 836 6116 843 6120
rect 856 5967 863 6083
rect 916 5896 923 5953
rect 756 5447 763 5533
rect 796 5483 803 5894
rect 896 5843 903 5863
rect 876 5836 903 5843
rect 876 5627 883 5836
rect 873 5600 887 5613
rect 876 5596 883 5600
rect 956 5567 963 5894
rect 856 5487 863 5563
rect 796 5476 813 5483
rect 816 5347 823 5473
rect 876 5376 883 5453
rect 747 5103 760 5107
rect 747 5093 763 5103
rect 756 5076 763 5093
rect 816 5046 823 5333
rect 736 4987 743 5043
rect 776 5007 783 5043
rect 656 4556 663 4560
rect 536 4527 543 4554
rect 396 4503 403 4523
rect 376 4496 403 4503
rect 376 4347 383 4496
rect 676 4467 683 4523
rect 396 4336 403 4413
rect 376 4047 383 4293
rect 416 4267 423 4303
rect 456 4247 463 4303
rect 516 4267 523 4313
rect 416 4036 423 4193
rect 356 3263 363 3513
rect 376 3307 383 3993
rect 396 3907 403 4003
rect 436 3987 443 4003
rect 436 3816 443 3973
rect 473 3820 487 3833
rect 476 3816 483 3820
rect 416 3727 423 3783
rect 456 3567 463 3783
rect 516 3647 523 3893
rect 536 3623 543 4453
rect 676 4348 683 4373
rect 636 4267 643 4303
rect 596 4036 603 4073
rect 556 4003 563 4034
rect 556 3996 583 4003
rect 556 3687 563 3813
rect 576 3747 583 3996
rect 616 3967 623 4003
rect 607 3936 633 3943
rect 516 3616 543 3623
rect 476 3516 483 3593
rect 356 3256 403 3263
rect 436 3260 443 3263
rect 433 3247 447 3260
rect 336 2488 343 3053
rect 396 2996 403 3233
rect 476 3107 483 3263
rect 516 3247 523 3616
rect 536 3267 543 3294
rect 576 3227 583 3553
rect 596 3528 603 3833
rect 616 3786 623 3873
rect 656 3847 663 3992
rect 696 3947 703 4013
rect 716 3887 723 4853
rect 736 4526 743 4553
rect 756 4507 763 4573
rect 736 4127 743 4334
rect 776 4107 783 4953
rect 856 4856 863 5213
rect 976 5187 983 5813
rect 996 5287 1003 5773
rect 1016 5347 1023 6114
rect 1036 6107 1043 6313
rect 1116 6116 1123 6293
rect 1196 6167 1203 6352
rect 1160 6123 1173 6127
rect 1156 6116 1173 6123
rect 1160 6113 1173 6116
rect 1096 5967 1103 6083
rect 1136 6063 1143 6083
rect 1116 6056 1143 6063
rect 1116 5908 1123 6056
rect 1096 5807 1103 5863
rect 1156 5747 1163 5863
rect 1056 5596 1063 5633
rect 1156 5627 1163 5673
rect 1093 5600 1107 5613
rect 1096 5596 1103 5600
rect 1116 5543 1123 5563
rect 1096 5536 1123 5543
rect 1133 5547 1147 5553
rect 1156 5547 1163 5613
rect 1036 5227 1043 5393
rect 896 4856 903 4893
rect 916 4867 923 5113
rect 956 5076 963 5113
rect 1036 4826 1043 5173
rect 796 4787 803 4812
rect 736 3847 743 3992
rect 647 3823 660 3827
rect 647 3816 663 3823
rect 647 3813 660 3816
rect 696 3516 743 3523
rect 416 2927 423 2963
rect 433 2947 447 2952
rect 436 2776 443 2933
rect 356 2746 363 2773
rect 456 2740 463 2743
rect 453 2727 467 2740
rect 396 2476 403 2693
rect 316 2163 323 2273
rect 376 2267 383 2432
rect 436 2287 443 2633
rect 456 2447 463 2553
rect 496 2447 503 2913
rect 516 2727 523 2833
rect 536 2707 543 3173
rect 556 2727 563 3093
rect 596 3067 603 3514
rect 616 2996 623 3294
rect 636 3127 643 3483
rect 596 2960 603 2963
rect 593 2947 607 2960
rect 656 2907 663 3053
rect 736 3007 743 3516
rect 756 3487 763 3713
rect 756 3266 763 3413
rect 776 3023 783 3773
rect 796 3103 803 4773
rect 836 4687 843 4823
rect 816 4207 823 4554
rect 836 4547 843 4673
rect 856 4607 863 4693
rect 916 4556 943 4563
rect 836 4307 843 4373
rect 876 4336 883 4493
rect 896 4467 903 4523
rect 916 4336 923 4373
rect 936 4367 943 4556
rect 956 4487 963 4533
rect 836 4036 843 4253
rect 936 4247 943 4292
rect 1056 4227 1063 5533
rect 1096 5407 1103 5536
rect 1116 5376 1123 5493
rect 1176 5376 1183 5893
rect 1196 5846 1203 6153
rect 1216 5747 1223 6113
rect 1276 5743 1283 6273
rect 1296 6247 1303 6356
rect 1436 6207 1443 6873
rect 1456 6606 1463 6933
rect 1516 6900 1523 6903
rect 1513 6887 1527 6900
rect 1556 6867 1563 6903
rect 1596 6827 1603 7636
rect 1633 7467 1647 7473
rect 1656 7467 1663 7993
rect 1676 7946 1683 7973
rect 1696 7627 1703 8053
rect 1756 7907 1763 8133
rect 1816 8127 1823 8213
rect 1856 8167 1863 8233
rect 1876 8063 1883 8616
rect 1867 8056 1883 8063
rect 1856 7976 1863 8053
rect 1796 7907 1803 7943
rect 1836 7940 1843 7943
rect 1833 7927 1847 7940
rect 1716 7487 1723 7753
rect 1776 7676 1783 7713
rect 1756 7607 1763 7643
rect 1736 7456 1743 7533
rect 1496 6487 1503 6813
rect 1596 6547 1603 6603
rect 1476 6396 1483 6453
rect 1296 6047 1303 6193
rect 1356 6116 1363 6193
rect 1393 6120 1407 6133
rect 1396 6116 1403 6120
rect 1336 6047 1343 6083
rect 1436 6047 1443 6193
rect 1336 5896 1343 5973
rect 1436 5907 1443 5933
rect 1456 5908 1463 6233
rect 1496 5866 1503 6473
rect 1533 6400 1547 6413
rect 1536 6396 1543 6400
rect 1616 6227 1623 6413
rect 1636 6287 1643 7432
rect 1656 6948 1663 7353
rect 1676 7247 1683 7423
rect 1716 7267 1723 7423
rect 1776 7367 1783 7613
rect 1796 7427 1803 7643
rect 1676 7067 1683 7154
rect 1696 7087 1703 7253
rect 1736 7156 1743 7213
rect 1816 7167 1823 7633
rect 1836 7327 1843 7892
rect 1856 7647 1863 7773
rect 1896 7567 1903 8593
rect 1936 8567 1943 8593
rect 1916 8467 1923 8494
rect 1936 8196 1943 8273
rect 2016 8067 2023 8972
rect 2096 8827 2103 9534
rect 2116 9187 2123 11243
rect 2276 11096 2283 11133
rect 2196 11047 2203 11094
rect 2356 11066 2363 11093
rect 2576 11086 2583 11133
rect 2596 11076 2623 11083
rect 2256 11027 2263 11063
rect 2476 11027 2483 11063
rect 2516 11043 2523 11052
rect 2516 11036 2543 11043
rect 2187 10796 2203 10803
rect 2176 10707 2183 10794
rect 2316 10787 2323 11013
rect 2296 10756 2323 10763
rect 2136 8907 2143 9593
rect 2156 9248 2163 10573
rect 2216 10507 2223 10543
rect 2216 10283 2223 10493
rect 2216 10276 2243 10283
rect 2256 10127 2263 10243
rect 2316 10227 2323 10756
rect 2416 10576 2423 10613
rect 2476 10607 2483 10763
rect 2453 10580 2467 10593
rect 2456 10576 2463 10580
rect 2236 10056 2243 10093
rect 2256 10020 2263 10023
rect 2253 10007 2267 10020
rect 2336 9967 2343 10274
rect 2196 9548 2203 9793
rect 2276 9756 2283 9933
rect 2256 9543 2263 9712
rect 2296 9703 2303 9723
rect 2276 9696 2303 9703
rect 2276 9627 2283 9696
rect 2236 9536 2263 9543
rect 2216 9287 2223 9503
rect 2256 9248 2263 9493
rect 2296 9387 2303 9633
rect 2316 9507 2323 9713
rect 2336 9507 2343 9953
rect 2356 9547 2363 10393
rect 2376 10187 2383 10573
rect 2536 10547 2543 11036
rect 2556 10987 2563 11043
rect 2556 10766 2563 10793
rect 2436 10467 2443 10543
rect 2476 10540 2483 10543
rect 2473 10527 2487 10540
rect 2376 10026 2383 10113
rect 2396 9983 2403 10093
rect 2416 10067 2423 10373
rect 2496 10327 2503 10533
rect 2556 10467 2563 10574
rect 2496 10276 2503 10313
rect 2476 10127 2483 10243
rect 2496 10056 2503 10093
rect 2536 10067 2543 10113
rect 2520 10023 2533 10027
rect 2476 10007 2483 10023
rect 2516 10016 2533 10023
rect 2520 10013 2533 10016
rect 2467 9996 2483 10007
rect 2467 9993 2480 9996
rect 2396 9976 2423 9983
rect 2376 9727 2383 9913
rect 2216 9127 2223 9203
rect 2276 9200 2283 9203
rect 2236 9016 2243 9193
rect 2273 9187 2287 9200
rect 2286 9180 2287 9187
rect 2216 8947 2223 8983
rect 1916 7927 1923 8053
rect 1916 7587 1923 7913
rect 1936 7646 1943 7793
rect 1996 7727 2003 7993
rect 2056 7988 2063 8813
rect 2176 8716 2183 8793
rect 2076 8467 2083 8714
rect 2116 8647 2123 8683
rect 2196 8567 2203 8613
rect 2216 8496 2223 8853
rect 2276 8787 2283 9173
rect 2276 8587 2283 8713
rect 2196 8407 2203 8463
rect 2236 8307 2243 8463
rect 2296 8367 2303 9173
rect 2316 8647 2323 9333
rect 2356 9206 2363 9533
rect 2336 9196 2353 9203
rect 2336 9087 2343 9196
rect 2376 9187 2383 9673
rect 2396 9627 2403 9773
rect 2416 9707 2423 9976
rect 2556 9887 2563 10054
rect 2436 9747 2443 9873
rect 2456 9767 2463 9873
rect 2493 9760 2507 9773
rect 2496 9756 2503 9760
rect 2536 9756 2543 9813
rect 2576 9788 2583 10973
rect 2616 10927 2623 11076
rect 2896 11076 2903 11153
rect 3136 11056 3163 11063
rect 2996 11027 3003 11053
rect 2756 10867 2763 10933
rect 2676 10796 2683 10853
rect 2713 10800 2727 10813
rect 2716 10796 2723 10800
rect 2596 10547 2603 10593
rect 2716 10576 2723 10693
rect 2756 10587 2763 10853
rect 3016 10816 3023 10973
rect 3136 10947 3143 11056
rect 2836 10707 2843 10813
rect 2953 10800 2967 10813
rect 2956 10796 2963 10800
rect 2976 10707 2983 10763
rect 2596 10067 2603 10453
rect 2656 10387 2663 10532
rect 2693 10527 2707 10532
rect 2756 10427 2763 10573
rect 2956 10367 2963 10574
rect 2636 10107 2643 10274
rect 2776 10246 2783 10273
rect 2696 10240 2703 10243
rect 2693 10227 2707 10240
rect 2756 10127 2763 10173
rect 2776 10147 2783 10232
rect 2756 10056 2763 10113
rect 2696 9887 2703 10023
rect 2736 10020 2743 10023
rect 2733 10007 2747 10020
rect 2796 10007 2803 10253
rect 2816 10247 2823 10313
rect 2976 10187 2983 10693
rect 3056 10387 3063 10783
rect 3076 10687 3083 10794
rect 3156 10576 3163 10673
rect 3136 10367 3143 10543
rect 2907 10093 2913 10107
rect 2853 10087 2867 10093
rect 2936 10056 2943 10173
rect 2876 9907 2883 9993
rect 2467 9723 2480 9727
rect 2636 9723 2643 9813
rect 2736 9736 2743 9793
rect 2467 9716 2483 9723
rect 2467 9713 2480 9716
rect 2436 9536 2443 9633
rect 2476 9536 2483 9693
rect 2516 9647 2523 9723
rect 2616 9716 2643 9723
rect 2396 9496 2423 9503
rect 2396 9107 2403 9496
rect 2456 9467 2463 9503
rect 2496 9236 2503 9273
rect 2416 9147 2423 9234
rect 2356 8747 2363 9093
rect 2416 9016 2423 9133
rect 2456 9016 2463 9173
rect 2436 8887 2443 8983
rect 2516 8927 2523 9203
rect 2576 9087 2583 9173
rect 2616 9127 2623 9716
rect 2876 9567 2883 9893
rect 2896 9807 2903 10053
rect 2956 9887 2963 10023
rect 2916 9707 2923 9743
rect 2880 9543 2893 9547
rect 2876 9536 2893 9543
rect 2880 9533 2893 9536
rect 2656 9187 2663 9492
rect 2696 9147 2703 9203
rect 2736 9200 2743 9203
rect 2733 9187 2747 9200
rect 2536 8867 2543 9033
rect 2556 8986 2563 9013
rect 2356 8716 2363 8733
rect 2433 8720 2447 8733
rect 2436 8716 2443 8720
rect 2316 8466 2323 8593
rect 2376 8567 2383 8683
rect 2416 8680 2423 8683
rect 2413 8667 2427 8680
rect 2376 8387 2383 8473
rect 2193 8200 2207 8213
rect 2196 8196 2203 8200
rect 2076 8007 2083 8194
rect 2236 8163 2243 8293
rect 2096 7976 2103 8033
rect 2136 7946 2143 8033
rect 2176 7988 2183 8163
rect 2216 8156 2243 8163
rect 2036 7787 2043 7943
rect 2033 7680 2047 7693
rect 2076 7688 2083 7873
rect 2096 7707 2103 7773
rect 2196 7747 2203 7893
rect 2036 7676 2043 7680
rect 2216 7687 2223 8156
rect 2316 8147 2323 8213
rect 2376 8208 2383 8373
rect 2396 8287 2403 8413
rect 2456 8347 2463 8494
rect 2276 7976 2283 8113
rect 2316 8087 2323 8133
rect 2336 8087 2343 8194
rect 2396 8027 2403 8163
rect 2413 8127 2427 8133
rect 2436 8107 2443 8153
rect 2236 7907 2243 7973
rect 2296 7940 2303 7943
rect 2336 7940 2343 7943
rect 2293 7927 2307 7940
rect 2333 7927 2347 7940
rect 2376 7927 2383 7993
rect 2396 7947 2403 7973
rect 2236 7896 2253 7907
rect 2240 7893 2253 7896
rect 2376 7867 2383 7913
rect 2016 7607 2023 7643
rect 1836 7127 1843 7253
rect 1856 7247 1863 7473
rect 1956 7423 1963 7454
rect 1936 7416 1963 7423
rect 1756 7087 1763 7123
rect 1776 6936 1783 6993
rect 1656 6687 1663 6934
rect 1756 6827 1763 6903
rect 1796 6900 1803 6903
rect 1793 6887 1807 6900
rect 1856 6887 1863 7153
rect 1876 7067 1883 7153
rect 1896 7126 1903 7193
rect 1516 6007 1523 6193
rect 1587 6143 1600 6147
rect 1587 6133 1603 6143
rect 1596 6116 1603 6133
rect 1513 5907 1527 5913
rect 1256 5736 1283 5743
rect 1236 5407 1243 5653
rect 1076 4687 1083 5074
rect 1116 5047 1123 5313
rect 1136 5267 1143 5343
rect 1176 5076 1183 5173
rect 1213 5080 1227 5093
rect 1216 5076 1223 5080
rect 1156 4947 1163 5043
rect 1256 5027 1263 5736
rect 1316 5596 1323 5833
rect 1356 5727 1363 5863
rect 1356 5563 1363 5713
rect 1296 5560 1303 5563
rect 1293 5547 1307 5560
rect 1336 5556 1363 5563
rect 1176 4967 1183 4993
rect 1276 4987 1283 5513
rect 1316 5287 1323 5413
rect 1336 5107 1343 5556
rect 1356 5447 1363 5473
rect 1396 5376 1403 5852
rect 1496 5596 1503 5793
rect 1536 5727 1543 6114
rect 1556 6076 1583 6083
rect 1556 5847 1563 6076
rect 1616 6027 1623 6083
rect 1596 5896 1603 5993
rect 1656 5967 1663 6673
rect 1836 6636 1843 6693
rect 1916 6607 1923 7033
rect 1936 7007 1943 7416
rect 1976 7387 1983 7573
rect 2076 7547 2083 7674
rect 2236 7676 2243 7833
rect 2316 7647 2323 7713
rect 2336 7676 2363 7683
rect 2336 7607 2343 7676
rect 2416 7627 2423 8073
rect 2436 7707 2443 8093
rect 2456 7827 2463 8333
rect 2476 7847 2483 8773
rect 2496 8687 2503 8833
rect 2496 8367 2503 8553
rect 2496 7987 2503 8353
rect 2516 8127 2523 8733
rect 2536 8728 2543 8793
rect 2536 8467 2543 8714
rect 2536 8008 2543 8453
rect 2556 8307 2563 8933
rect 2576 8427 2583 9073
rect 2696 9028 2703 9112
rect 2676 8980 2683 8983
rect 2673 8967 2687 8980
rect 2716 8947 2723 8983
rect 2636 8527 2643 8683
rect 2676 8567 2683 8613
rect 2696 8607 2703 8653
rect 2716 8647 2723 8853
rect 2636 8496 2643 8513
rect 2696 8467 2703 8593
rect 2616 8387 2623 8463
rect 2696 8163 2703 8413
rect 2736 8227 2743 8973
rect 2756 8847 2763 9014
rect 2776 8966 2783 9333
rect 2856 9303 2863 9503
rect 2836 9296 2863 9303
rect 2836 9247 2843 9296
rect 2916 9267 2923 9653
rect 2936 9347 2943 9773
rect 2996 9587 3003 10023
rect 3056 9987 3063 10352
rect 3076 10247 3083 10353
rect 3116 10276 3123 10313
rect 3176 10240 3183 10243
rect 3173 10227 3187 10240
rect 3216 10207 3223 10574
rect 3236 10247 3243 10313
rect 3296 10227 3303 10613
rect 3316 10587 3323 11094
rect 3376 11047 3383 11133
rect 3476 11096 3483 11133
rect 3396 11067 3403 11094
rect 3456 11060 3463 11063
rect 3496 11060 3503 11063
rect 3453 11047 3467 11060
rect 3493 11047 3507 11060
rect 3356 10727 3363 10783
rect 3376 10767 3383 10813
rect 3433 10783 3447 10793
rect 3416 10780 3447 10783
rect 3416 10776 3443 10780
rect 3376 10627 3383 10753
rect 3316 10536 3343 10543
rect 3316 10507 3323 10536
rect 3416 10527 3423 10776
rect 3136 10007 3143 10173
rect 2956 9467 2963 9573
rect 3056 9567 3063 9873
rect 3116 9827 3123 9853
rect 3056 9536 3063 9553
rect 2976 9267 2983 9533
rect 2996 9487 3003 9533
rect 3116 9507 3123 9754
rect 3136 9667 3143 9993
rect 3156 9847 3163 10133
rect 3196 10020 3203 10023
rect 3193 10007 3207 10020
rect 3236 9987 3243 10023
rect 3176 9867 3183 9933
rect 3216 9756 3223 9953
rect 2796 8987 2803 9053
rect 2816 8967 2823 9013
rect 2856 8907 2863 9253
rect 2907 9243 2920 9247
rect 2907 9236 2923 9243
rect 2907 9233 2920 9236
rect 2996 9247 3003 9452
rect 3136 9367 3143 9553
rect 2876 9063 2883 9233
rect 3016 9207 3023 9234
rect 2980 9203 2993 9207
rect 2936 9167 2943 9203
rect 2976 9196 2993 9203
rect 2980 9193 2993 9196
rect 3096 9127 3103 9253
rect 3136 9243 3143 9353
rect 3196 9307 3203 9723
rect 3216 9287 3223 9693
rect 3256 9536 3263 9953
rect 3296 9587 3303 10053
rect 3316 9947 3323 10493
rect 3356 10276 3363 10513
rect 3396 10276 3403 10373
rect 3436 10276 3443 10573
rect 3456 10387 3463 10973
rect 3476 10547 3483 11013
rect 3336 9727 3343 10232
rect 3376 9967 3383 10243
rect 3436 10056 3443 10193
rect 3476 10068 3483 10273
rect 3516 10027 3523 11052
rect 3536 11047 3543 11093
rect 3796 11083 3803 11153
rect 3856 11086 3863 11133
rect 3796 11076 3823 11083
rect 3716 11027 3723 11052
rect 3796 11043 3803 11076
rect 4096 11076 4123 11083
rect 3776 11036 3803 11043
rect 3676 10547 3683 10783
rect 3716 10767 3723 10853
rect 3736 10747 3743 10783
rect 3776 10747 3783 11036
rect 4096 10927 4103 11076
rect 4356 11056 4363 11243
rect 4396 11096 4423 11103
rect 4416 11065 4423 11096
rect 4416 11058 4584 11065
rect 4156 10987 4163 11043
rect 4597 11022 4604 11104
rect 4236 11015 4604 11022
rect 4036 10780 4043 10783
rect 3556 10540 3563 10543
rect 3536 10247 3543 10532
rect 3553 10527 3567 10540
rect 3596 10507 3603 10543
rect 3576 10267 3583 10393
rect 3676 10296 3683 10373
rect 3613 10287 3627 10293
rect 3607 10280 3627 10287
rect 3607 10276 3623 10280
rect 3607 10273 3620 10276
rect 3716 10167 3723 10213
rect 3416 9967 3423 10023
rect 3456 9907 3463 10023
rect 3536 9947 3543 10153
rect 3636 9987 3643 10073
rect 3736 10027 3743 10733
rect 4016 10576 4023 10774
rect 4033 10767 4047 10780
rect 3936 10546 3943 10573
rect 3776 10407 3783 10543
rect 3827 10536 3843 10543
rect 3836 10323 3843 10536
rect 4096 10407 4103 10574
rect 4116 10347 4123 10873
rect 4156 10827 4163 10973
rect 4136 10627 4143 10783
rect 4176 10767 4183 10913
rect 4196 10747 4203 10783
rect 4236 10707 4243 11015
rect 4567 10913 4573 10927
rect 4476 10783 4483 10913
rect 4716 10844 4723 11243
rect 4776 11096 4783 11133
rect 4796 11063 4803 11243
rect 4796 11056 4824 11063
rect 4716 10837 4783 10844
rect 4776 10796 4783 10837
rect 4476 10776 4503 10783
rect 4736 10743 4743 10763
rect 4736 10736 4763 10743
rect 4196 10546 4203 10693
rect 4236 10576 4243 10613
rect 4296 10546 4303 10613
rect 4576 10546 4583 10573
rect 3816 10316 3843 10323
rect 3816 10267 3823 10316
rect 3876 10056 3883 10153
rect 3393 9760 3407 9773
rect 3396 9756 3403 9760
rect 3476 9723 3483 9754
rect 3496 9727 3503 9773
rect 3416 9647 3423 9723
rect 3456 9716 3483 9723
rect 3293 9540 3307 9552
rect 3296 9536 3303 9540
rect 3316 9496 3343 9503
rect 3116 9236 3143 9243
rect 3173 9240 3187 9253
rect 3176 9236 3183 9240
rect 3116 9187 3123 9236
rect 3156 9200 3163 9203
rect 3153 9187 3167 9200
rect 3276 9167 3283 9192
rect 2876 9056 2903 9063
rect 2896 9028 2903 9056
rect 2996 8996 3023 9003
rect 2776 8867 2783 8893
rect 2856 8716 2863 8872
rect 2916 8827 2923 8983
rect 2933 8747 2947 8753
rect 2936 8716 2943 8733
rect 2816 8667 2823 8693
rect 2876 8680 2883 8683
rect 2916 8680 2923 8683
rect 2873 8667 2887 8680
rect 2913 8667 2927 8680
rect 2756 8587 2763 8613
rect 2776 8367 2783 8653
rect 2836 8607 2843 8633
rect 2796 8527 2803 8573
rect 2916 8466 2923 8533
rect 2836 8460 2843 8463
rect 2833 8447 2847 8460
rect 2976 8447 2983 8893
rect 3016 8847 3023 8996
rect 3116 8927 3123 9003
rect 2996 8747 3003 8773
rect 3036 8687 3043 8853
rect 3136 8827 3143 8853
rect 3136 8716 3143 8813
rect 3176 8716 3183 8793
rect 3216 8767 3223 8813
rect 3256 8807 3263 9093
rect 3276 9007 3283 9153
rect 3296 9067 3303 9273
rect 3316 9248 3323 9473
rect 3296 8996 3303 9053
rect 3193 8607 3207 8613
rect 3076 8496 3083 8533
rect 3100 8463 3113 8467
rect 3056 8407 3063 8463
rect 3096 8456 3113 8463
rect 3100 8453 3113 8456
rect 3096 8247 3103 8433
rect 2716 8176 2733 8183
rect 2576 7976 2583 8133
rect 2596 8067 2603 8163
rect 2696 8156 2723 8163
rect 2556 7927 2563 7943
rect 2547 7916 2563 7927
rect 2547 7913 2560 7916
rect 2596 7807 2603 7943
rect 2636 7807 2643 8113
rect 2676 7847 2683 7993
rect 2016 7407 2023 7533
rect 2036 7267 2043 7533
rect 2056 7367 2063 7473
rect 2116 7456 2123 7573
rect 2216 7487 2223 7513
rect 2153 7460 2167 7473
rect 2156 7456 2163 7460
rect 2216 7447 2223 7473
rect 2236 7436 2243 7533
rect 2256 7446 2263 7573
rect 2096 7420 2103 7423
rect 2093 7407 2107 7420
rect 2016 6936 2023 6973
rect 1996 6867 2003 6903
rect 2016 6636 2023 6873
rect 2076 6827 2083 7373
rect 2096 7147 2103 7333
rect 2116 7107 2123 7273
rect 2076 6648 2083 6813
rect 1816 6547 1823 6603
rect 2036 6600 2043 6603
rect 2033 6587 2047 6600
rect 2076 6587 2083 6634
rect 1676 6383 1683 6513
rect 1676 6376 1703 6383
rect 1676 6067 1683 6173
rect 1656 5767 1663 5863
rect 1476 5507 1483 5563
rect 1433 5380 1447 5393
rect 1516 5388 1523 5563
rect 1536 5487 1543 5533
rect 1436 5376 1443 5380
rect 1376 5340 1383 5343
rect 1373 5327 1387 5340
rect 1373 5307 1387 5313
rect 1136 4827 1143 4893
rect 1356 4887 1363 5213
rect 1416 5076 1423 5153
rect 1096 4727 1103 4823
rect 1216 4767 1223 4823
rect 1296 4587 1303 4853
rect 1296 4556 1303 4573
rect 1096 4487 1103 4523
rect 1116 4336 1123 4493
rect 856 3967 863 4003
rect 936 3816 943 4212
rect 1073 4040 1087 4053
rect 1076 4036 1083 4040
rect 996 4003 1003 4034
rect 1136 4006 1143 4153
rect 1196 4147 1203 4334
rect 1216 4087 1223 4353
rect 996 3996 1023 4003
rect 816 3187 823 3753
rect 856 3627 863 3813
rect 916 3780 923 3783
rect 913 3767 927 3780
rect 876 3567 883 3713
rect 956 3667 963 3783
rect 996 3687 1003 3814
rect 916 3516 923 3553
rect 936 3547 943 3593
rect 836 3127 843 3514
rect 956 3427 963 3513
rect 976 3486 983 3613
rect 916 3296 923 3373
rect 956 3296 963 3333
rect 796 3096 813 3103
rect 756 3016 783 3023
rect 633 2780 647 2793
rect 636 2776 643 2780
rect 393 2260 407 2273
rect 433 2260 447 2273
rect 396 2256 403 2260
rect 436 2256 443 2260
rect 316 2156 343 2163
rect 196 1436 203 1493
rect 96 367 103 1392
rect 176 1383 183 1403
rect 176 1376 203 1383
rect 196 1367 203 1376
rect 336 1367 343 2156
rect 396 1956 403 2053
rect 376 1887 383 1923
rect 416 1436 423 1593
rect 196 1216 203 1353
rect 396 1327 403 1403
rect 416 1216 423 1353
rect 176 947 183 1183
rect 216 1163 223 1172
rect 196 1156 223 1163
rect 136 708 143 933
rect 196 916 203 1156
rect 436 927 443 1183
rect 236 887 243 914
rect 247 876 263 883
rect 256 767 263 876
rect 196 696 203 733
rect 136 666 143 694
rect 176 627 183 663
rect 216 467 223 652
rect 256 627 263 753
rect 456 708 463 914
rect 456 667 463 694
rect 476 666 483 1673
rect 496 1367 503 1912
rect 516 1748 523 2613
rect 536 2587 543 2693
rect 656 2627 663 2743
rect 536 2287 543 2533
rect 593 2480 607 2493
rect 596 2476 603 2480
rect 616 2327 623 2443
rect 676 2427 683 2713
rect 696 2687 703 2743
rect 696 2367 703 2673
rect 516 1327 523 1734
rect 516 887 523 1313
rect 200 403 213 407
rect 196 396 213 403
rect 116 227 123 394
rect 200 393 213 396
rect 376 396 383 433
rect 176 176 183 213
rect 336 187 343 393
rect 456 347 463 433
rect 416 227 423 273
rect 416 176 423 213
rect 456 147 463 333
rect 196 140 203 143
rect 193 127 207 140
rect 476 127 483 652
rect 536 367 543 1873
rect 556 1227 563 2273
rect 576 2226 583 2293
rect 636 2256 643 2353
rect 716 2307 723 2493
rect 616 1956 623 2033
rect 656 1967 663 2223
rect 696 1926 703 2113
rect 616 1736 623 1793
rect 596 1667 603 1703
rect 636 1436 643 1633
rect 656 1227 663 1403
rect 616 880 623 883
rect 613 867 627 880
rect 616 696 623 753
rect 676 747 683 1214
rect 696 867 703 1912
rect 716 1607 723 1954
rect 736 1887 743 2533
rect 756 2488 763 3016
rect 816 2996 823 3093
rect 796 2887 803 2963
rect 836 2943 843 2963
rect 816 2940 843 2943
rect 816 2936 847 2940
rect 796 2547 803 2873
rect 816 2627 823 2936
rect 833 2927 847 2936
rect 876 2827 883 3113
rect 896 2947 903 3263
rect 916 3187 923 3213
rect 916 2967 923 3173
rect 936 3007 943 3263
rect 996 3247 1003 3652
rect 936 2867 943 2993
rect 836 2746 843 2813
rect 896 2776 903 2853
rect 956 2843 963 3233
rect 1016 3227 1023 3996
rect 1216 3927 1223 4033
rect 1236 4003 1243 4513
rect 1276 4347 1283 4523
rect 1296 4047 1303 4493
rect 1316 4487 1323 4523
rect 1376 4507 1383 4554
rect 1353 4340 1367 4353
rect 1356 4336 1363 4340
rect 1436 4306 1443 4573
rect 1336 4267 1343 4303
rect 1316 4048 1323 4233
rect 1347 4053 1353 4067
rect 1376 4036 1383 4093
rect 1236 3996 1263 4003
rect 1276 4000 1283 4003
rect 1036 3327 1043 3673
rect 1056 3467 1063 3913
rect 1076 3786 1083 3893
rect 1136 3816 1143 3893
rect 1216 3787 1223 3853
rect 1140 3483 1153 3487
rect 1136 3476 1153 3483
rect 1140 3473 1153 3476
rect 1216 3467 1223 3752
rect 1236 3467 1243 3973
rect 1096 3307 1103 3451
rect 1256 3347 1263 3996
rect 1273 3987 1287 4000
rect 1036 2996 1043 3292
rect 1056 3027 1063 3294
rect 1213 3300 1227 3313
rect 1216 3296 1223 3300
rect 1176 3256 1203 3263
rect 1060 2963 1073 2967
rect 936 2836 963 2843
rect 936 2776 943 2836
rect 896 2547 903 2573
rect 776 2347 783 2493
rect 813 2480 827 2493
rect 816 2476 823 2480
rect 836 2440 843 2443
rect 833 2427 847 2440
rect 916 2423 923 2743
rect 936 2446 943 2513
rect 916 2416 943 2423
rect 756 2227 763 2253
rect 796 2207 803 2373
rect 836 2256 843 2293
rect 876 2287 883 2313
rect 873 2260 887 2273
rect 876 2256 883 2260
rect 856 2220 863 2223
rect 896 2220 923 2223
rect 853 2207 867 2220
rect 896 2216 927 2220
rect 913 2207 927 2216
rect 756 1927 763 2192
rect 936 1987 943 2416
rect 956 2227 963 2273
rect 736 1467 743 1793
rect 816 1787 823 1833
rect 833 1740 847 1753
rect 836 1736 843 1740
rect 776 1527 783 1733
rect 876 1707 883 1954
rect 816 1607 823 1703
rect 936 1627 943 1973
rect 596 607 603 663
rect 736 547 743 1453
rect 853 1440 867 1453
rect 856 1436 863 1440
rect 776 1187 783 1434
rect 836 1327 843 1403
rect 956 1367 963 2133
rect 976 2127 983 2793
rect 996 2147 1003 2953
rect 1016 2907 1023 2963
rect 1056 2956 1073 2963
rect 1060 2953 1073 2956
rect 1116 2947 1123 3013
rect 1036 2387 1043 2873
rect 1056 2727 1063 2933
rect 1076 2807 1083 2932
rect 1116 2776 1123 2893
rect 1136 2863 1143 3133
rect 1156 2887 1163 3213
rect 1176 2927 1183 3256
rect 1276 3243 1283 3873
rect 1296 3767 1303 3993
rect 1313 3847 1327 3853
rect 1376 3816 1383 3893
rect 1396 3887 1403 4253
rect 1456 4247 1463 4613
rect 1476 4527 1483 5074
rect 1496 4767 1503 5373
rect 1516 5307 1523 5374
rect 1536 5327 1543 5473
rect 1576 5347 1583 5594
rect 1596 5387 1603 5693
rect 1676 5376 1683 5552
rect 1696 5547 1703 6376
rect 1736 6367 1743 6383
rect 1736 6327 1743 6353
rect 1716 5407 1723 6253
rect 1736 6086 1743 6313
rect 1816 6147 1823 6533
rect 1836 6116 1843 6473
rect 1956 6416 1963 6473
rect 1876 6367 1883 6414
rect 1936 6367 1943 6383
rect 1936 6356 1953 6367
rect 1940 6353 1953 6356
rect 1776 6080 1783 6083
rect 1773 6067 1787 6080
rect 1736 5866 1743 6033
rect 1736 5596 1743 5733
rect 1776 5667 1783 5953
rect 1816 5903 1823 6083
rect 1896 5987 1903 6133
rect 1796 5896 1823 5903
rect 1796 5643 1803 5896
rect 1896 5903 1903 5973
rect 1876 5896 1903 5903
rect 1856 5847 1863 5863
rect 1916 5847 1923 6213
rect 1936 6107 1943 6233
rect 1956 6187 1963 6313
rect 1956 6083 1963 6113
rect 1936 6076 1963 6083
rect 1856 5836 1873 5847
rect 1860 5833 1873 5836
rect 1796 5636 1823 5643
rect 1793 5600 1807 5613
rect 1816 5607 1823 5636
rect 1796 5596 1803 5600
rect 1876 5567 1883 5613
rect 1896 5507 1903 5573
rect 1936 5507 1943 6076
rect 1996 5923 2003 6573
rect 2096 6527 2103 7053
rect 2116 7047 2123 7072
rect 2136 6867 2143 7253
rect 2156 7167 2163 7233
rect 2196 7188 2203 7403
rect 2236 7156 2243 7313
rect 2496 7307 2503 7613
rect 2516 7547 2523 7793
rect 2656 7787 2663 7833
rect 2553 7680 2567 7693
rect 2556 7676 2563 7680
rect 2596 7676 2603 7772
rect 2647 7674 2653 7687
rect 2640 7673 2653 7674
rect 2576 7640 2583 7643
rect 2536 7507 2543 7633
rect 2573 7627 2587 7640
rect 2576 7527 2583 7613
rect 2596 7547 2603 7593
rect 2613 7463 2627 7473
rect 2596 7460 2627 7463
rect 2596 7456 2623 7460
rect 2536 7436 2563 7443
rect 2596 7436 2603 7456
rect 2556 7387 2563 7436
rect 2336 7147 2343 7293
rect 2176 7027 2183 7123
rect 2296 7083 2303 7133
rect 2316 7107 2323 7143
rect 2296 7076 2323 7083
rect 2236 6936 2243 6973
rect 2113 6567 2127 6573
rect 2136 6507 2143 6853
rect 2156 6707 2163 6934
rect 2216 6867 2223 6903
rect 2256 6900 2263 6903
rect 2253 6887 2267 6900
rect 2216 6636 2223 6693
rect 2276 6606 2283 6653
rect 2036 6207 2043 6273
rect 2056 6116 2063 6493
rect 2096 6116 2103 6413
rect 2153 6367 2167 6372
rect 2196 6307 2203 6383
rect 2276 6347 2283 6513
rect 2296 6428 2303 6953
rect 2316 6948 2323 7076
rect 2156 6187 2163 6293
rect 2133 6140 2147 6153
rect 2156 6147 2163 6173
rect 2136 6136 2143 6140
rect 2076 6027 2083 6083
rect 1996 5916 2013 5923
rect 1956 5707 1963 5873
rect 2016 5687 2023 5913
rect 2076 5896 2083 5992
rect 2056 5860 2063 5863
rect 2053 5847 2067 5860
rect 2066 5840 2067 5847
rect 2096 5843 2103 5863
rect 2096 5836 2123 5843
rect 2073 5827 2087 5833
rect 2116 5727 2123 5836
rect 2156 5627 2163 5893
rect 2176 5627 2183 5933
rect 2196 5866 2203 6233
rect 2296 6127 2303 6414
rect 2316 6227 2323 6934
rect 2396 6906 2403 6973
rect 2493 6940 2507 6953
rect 2496 6936 2503 6940
rect 2476 6900 2483 6903
rect 2516 6900 2543 6903
rect 2396 6767 2403 6892
rect 2473 6887 2487 6900
rect 2516 6896 2547 6900
rect 2533 6887 2547 6896
rect 2356 6606 2363 6673
rect 2396 6667 2403 6753
rect 2456 6707 2463 6813
rect 2456 6636 2463 6693
rect 2436 6567 2443 6603
rect 2396 6416 2403 6493
rect 2376 6380 2383 6383
rect 2416 6380 2443 6383
rect 2373 6367 2387 6380
rect 2416 6376 2447 6380
rect 2433 6367 2447 6376
rect 2426 6353 2427 6360
rect 2413 6347 2427 6353
rect 2456 6147 2463 6473
rect 2476 6387 2483 6513
rect 2287 6103 2300 6107
rect 2287 6096 2303 6103
rect 2287 6093 2300 6096
rect 2216 5747 2223 5993
rect 2316 5896 2323 5973
rect 2356 5896 2363 5993
rect 2396 5887 2403 5993
rect 2336 5860 2343 5863
rect 2333 5847 2347 5860
rect 2053 5600 2067 5613
rect 2093 5600 2107 5613
rect 2056 5596 2063 5600
rect 2096 5596 2103 5600
rect 1816 5346 1823 5393
rect 1836 5387 1843 5453
rect 1876 5376 1883 5413
rect 1587 5336 1623 5343
rect 1656 5340 1663 5343
rect 1536 4627 1543 5233
rect 1556 4787 1563 5113
rect 1596 5088 1603 5336
rect 1653 5327 1667 5340
rect 1636 5107 1643 5173
rect 1633 5080 1647 5093
rect 1636 5076 1643 5080
rect 1616 5040 1623 5043
rect 1613 5027 1627 5040
rect 1656 4927 1663 5043
rect 1696 4967 1703 5173
rect 1856 5167 1863 5343
rect 1576 4607 1583 4854
rect 1596 4827 1603 4913
rect 1716 4826 1723 5074
rect 1596 4587 1603 4813
rect 1636 4687 1643 4823
rect 1676 4707 1683 4753
rect 1696 4647 1703 4713
rect 1533 4560 1547 4573
rect 1536 4556 1543 4560
rect 1516 4348 1523 4523
rect 1596 4520 1603 4523
rect 1593 4507 1607 4520
rect 1576 4336 1603 4343
rect 1416 3828 1423 4093
rect 1436 4006 1443 4173
rect 1396 3707 1403 3783
rect 1456 3747 1463 3992
rect 1476 3767 1483 4053
rect 1496 3807 1503 4293
rect 1516 4107 1523 4334
rect 1576 4207 1583 4336
rect 1636 4300 1643 4303
rect 1633 4287 1647 4300
rect 1676 4247 1683 4573
rect 1696 4467 1703 4593
rect 1696 4287 1703 4334
rect 1576 4167 1583 4193
rect 1616 4036 1623 4173
rect 1676 4107 1683 4233
rect 1673 4043 1687 4053
rect 1656 4040 1687 4043
rect 1656 4036 1683 4040
rect 1336 3516 1343 3573
rect 1380 3523 1393 3527
rect 1376 3516 1393 3523
rect 1380 3513 1393 3516
rect 1307 3484 1320 3487
rect 1307 3477 1323 3484
rect 1307 3473 1320 3477
rect 1296 3267 1303 3452
rect 1356 3447 1363 3483
rect 1256 3236 1283 3243
rect 1136 2856 1163 2863
rect 1156 2788 1163 2856
rect 1076 2647 1083 2772
rect 1196 2747 1203 3193
rect 1256 2996 1263 3236
rect 1296 3067 1303 3253
rect 1316 3227 1323 3433
rect 1316 3087 1323 3213
rect 1316 2967 1323 3033
rect 1336 3007 1343 3333
rect 1227 2963 1240 2967
rect 1227 2953 1243 2963
rect 1276 2960 1283 2963
rect 1116 2647 1123 2713
rect 1127 2636 1143 2643
rect 1116 2476 1123 2533
rect 1096 2387 1103 2432
rect 1016 2207 1023 2333
rect 1036 2267 1043 2293
rect 1056 2256 1063 2373
rect 1096 2307 1103 2333
rect 1113 2263 1127 2273
rect 1096 2260 1127 2263
rect 1096 2256 1123 2260
rect 996 1827 1003 2093
rect 1076 1956 1083 2073
rect 1116 1887 1123 1953
rect 976 1547 983 1753
rect 1033 1740 1047 1753
rect 1036 1736 1043 1740
rect 1056 1647 1063 1703
rect 1096 1687 1103 1853
rect 1093 1667 1107 1673
rect 1033 1440 1047 1453
rect 1036 1436 1043 1440
rect 836 1228 843 1273
rect 1056 1216 1063 1353
rect 856 1143 863 1183
rect 1036 1163 1043 1183
rect 1036 1156 1053 1163
rect 856 1136 883 1143
rect 876 1007 883 1136
rect 816 823 823 883
rect 816 816 843 823
rect 816 696 823 793
rect 836 787 843 816
rect 836 647 843 663
rect 876 647 883 993
rect 916 647 923 953
rect 936 667 943 914
rect 976 666 983 853
rect 596 396 603 533
rect 576 360 583 363
rect 573 347 587 360
rect 616 343 623 363
rect 596 336 623 343
rect 596 307 603 336
rect 756 327 763 453
rect 816 396 823 633
rect 836 607 843 633
rect 876 366 883 612
rect 596 188 603 293
rect 796 267 803 363
rect 836 287 843 363
rect 756 147 763 253
rect 816 176 823 213
rect 876 156 883 352
rect 836 107 843 143
rect 916 107 923 273
rect 976 227 983 652
rect 996 627 1003 883
rect 1056 847 1063 1153
rect 1076 967 1083 1183
rect 1116 1167 1123 1873
rect 1136 1867 1143 2636
rect 1156 2187 1163 2213
rect 1176 2047 1183 2693
rect 1156 1926 1163 1954
rect 1196 1927 1203 2653
rect 1136 1706 1143 1793
rect 1156 1448 1163 1912
rect 1216 1903 1223 2893
rect 1236 2587 1243 2953
rect 1273 2947 1287 2960
rect 1356 2776 1363 3373
rect 1376 3247 1383 3293
rect 1376 2947 1383 2994
rect 1396 2907 1403 3453
rect 1416 3367 1423 3533
rect 1476 3527 1483 3753
rect 1516 3747 1523 4034
rect 1636 4000 1643 4003
rect 1633 3987 1647 4000
rect 1576 3687 1583 3783
rect 1576 3607 1583 3673
rect 1593 3520 1607 3533
rect 1596 3516 1603 3520
rect 1436 3296 1443 3393
rect 1516 3227 1523 3513
rect 1376 2647 1383 2743
rect 1236 2407 1243 2513
rect 1396 2488 1403 2733
rect 1256 2347 1263 2474
rect 1256 2223 1263 2293
rect 1256 2216 1283 2223
rect 1236 2067 1243 2212
rect 1336 2167 1343 2223
rect 1316 2047 1323 2073
rect 1296 1968 1303 2013
rect 1247 1963 1260 1967
rect 1247 1956 1263 1963
rect 1247 1953 1260 1956
rect 1196 1896 1223 1903
rect 1156 928 1163 1434
rect 1196 1147 1203 1896
rect 1336 1763 1343 1953
rect 1316 1756 1343 1763
rect 1236 1700 1243 1703
rect 1233 1687 1247 1700
rect 1276 1647 1283 1703
rect 1227 1633 1233 1647
rect 1276 1436 1283 1612
rect 1316 1447 1323 1756
rect 1216 1407 1223 1433
rect 1336 1406 1343 1633
rect 1356 1507 1363 2353
rect 1376 1963 1383 2313
rect 1396 2087 1403 2474
rect 1396 1987 1403 2073
rect 1376 1956 1403 1963
rect 1296 1367 1303 1403
rect 1276 1216 1283 1353
rect 1196 916 1203 953
rect 1236 916 1243 993
rect 1256 927 1263 1183
rect 1036 696 1043 733
rect 1096 696 1103 813
rect 1156 607 1163 914
rect 1036 396 1043 593
rect 1056 327 1063 363
rect 1136 347 1143 513
rect 1236 396 1243 833
rect 1276 667 1283 1133
rect 1296 1007 1303 1183
rect 1336 787 1343 914
rect 1356 887 1363 993
rect 1376 807 1383 1773
rect 1396 1367 1403 1956
rect 1416 1787 1423 3213
rect 1536 3207 1543 3473
rect 1636 3483 1643 3933
rect 1696 3827 1703 4273
rect 1716 4207 1723 4812
rect 1736 4727 1743 5093
rect 1876 5076 1883 5113
rect 1893 5027 1907 5032
rect 1756 4587 1763 4993
rect 1896 4887 1903 4933
rect 1893 4860 1907 4873
rect 1936 4868 1943 5053
rect 1896 4856 1903 4860
rect 1776 4787 1783 4853
rect 1936 4823 1943 4854
rect 1773 4747 1787 4752
rect 1876 4627 1883 4823
rect 1916 4816 1943 4823
rect 1896 4687 1903 4793
rect 1773 4560 1787 4573
rect 1813 4560 1827 4573
rect 1776 4556 1783 4560
rect 1816 4556 1823 4560
rect 1756 4487 1763 4523
rect 1796 4520 1803 4523
rect 1793 4507 1807 4520
rect 1856 4487 1863 4573
rect 1876 4527 1883 4592
rect 1716 3987 1723 4093
rect 1616 3476 1643 3483
rect 1576 3327 1583 3393
rect 1576 3147 1583 3313
rect 1596 3227 1603 3293
rect 1416 1567 1423 1733
rect 1436 1363 1443 2432
rect 1456 2367 1463 2933
rect 1556 2907 1563 2993
rect 1616 2907 1623 3476
rect 1656 3307 1663 3533
rect 1696 3487 1703 3613
rect 1716 3327 1723 3793
rect 1776 3707 1783 4253
rect 1896 4107 1903 4673
rect 1836 4036 1843 4093
rect 1673 3300 1687 3313
rect 1676 3296 1683 3300
rect 1736 3296 1743 3593
rect 1753 3520 1767 3533
rect 1756 3516 1763 3520
rect 1816 3447 1823 3733
rect 1807 3353 1813 3367
rect 1836 3363 1843 3693
rect 1856 3667 1863 3833
rect 1896 3607 1903 4053
rect 1916 3947 1923 4816
rect 1956 4807 1963 5433
rect 1976 5007 1983 5093
rect 1996 5047 2003 5493
rect 2176 5487 2183 5613
rect 2216 5587 2223 5733
rect 2436 5707 2443 6113
rect 2496 6103 2503 6453
rect 2516 6267 2523 6873
rect 2536 6567 2543 6852
rect 2556 6827 2563 7013
rect 2576 6887 2583 7233
rect 2596 7187 2603 7373
rect 2616 7367 2623 7433
rect 2636 7427 2643 7473
rect 2676 7387 2683 7812
rect 2696 7787 2703 8113
rect 2696 7646 2703 7673
rect 2616 6947 2623 7132
rect 2636 6967 2643 7333
rect 2676 7087 2683 7143
rect 2676 6987 2683 7073
rect 2696 6967 2703 7253
rect 2716 7127 2723 8156
rect 2736 8007 2743 8173
rect 2756 8027 2763 8233
rect 3016 8127 3023 8183
rect 2796 7976 2803 8013
rect 2836 7976 2843 8033
rect 2736 7627 2743 7972
rect 2756 7936 2783 7943
rect 2816 7940 2823 7943
rect 2756 7867 2763 7936
rect 2813 7927 2827 7940
rect 2796 7867 2803 7913
rect 2756 7607 2763 7832
rect 2816 7727 2823 7793
rect 2776 7646 2783 7713
rect 2816 7676 2823 7713
rect 2856 7676 2863 7913
rect 2896 7907 2903 8033
rect 2936 7946 2943 8033
rect 2876 7707 2883 7773
rect 2896 7688 2903 7872
rect 2916 7747 2923 7773
rect 2796 7587 2803 7633
rect 2876 7627 2883 7643
rect 2887 7616 2903 7623
rect 2756 7126 2763 7493
rect 2793 7460 2807 7473
rect 2796 7456 2803 7460
rect 2856 7427 2863 7533
rect 2776 7027 2783 7154
rect 2647 6956 2663 6963
rect 2556 6606 2563 6753
rect 2536 6207 2543 6453
rect 2556 6367 2563 6533
rect 2576 6467 2583 6852
rect 2636 6767 2643 6892
rect 2656 6847 2663 6956
rect 2716 6936 2723 6973
rect 2796 6903 2803 7353
rect 2613 6640 2627 6653
rect 2616 6636 2623 6640
rect 2656 6636 2663 6812
rect 2696 6636 2703 6833
rect 2736 6827 2743 6903
rect 2776 6896 2803 6903
rect 2636 6447 2643 6553
rect 2676 6547 2683 6603
rect 2653 6420 2667 6433
rect 2656 6416 2663 6420
rect 2716 6387 2723 6473
rect 2736 6407 2743 6792
rect 2756 6443 2763 6753
rect 2776 6547 2783 6896
rect 2796 6587 2803 6653
rect 2816 6547 2823 7373
rect 2836 6807 2843 7393
rect 2876 7307 2883 7573
rect 2896 7367 2903 7616
rect 2936 7267 2943 7793
rect 2956 7247 2963 8053
rect 2973 8027 2987 8033
rect 3016 8003 3023 8073
rect 2996 7996 3023 8003
rect 2996 7976 3003 7996
rect 3036 7976 3043 8153
rect 3096 8127 3103 8212
rect 3116 8087 3123 8213
rect 3136 8087 3143 8393
rect 3056 7940 3063 7943
rect 3016 7847 3023 7932
rect 3053 7927 3067 7940
rect 2976 7467 2983 7713
rect 3016 7587 3023 7833
rect 3073 7680 3087 7693
rect 3116 7688 3123 8073
rect 3136 7947 3143 7974
rect 3156 7927 3163 8493
rect 3216 8467 3223 8714
rect 3256 8686 3263 8753
rect 3196 8167 3203 8293
rect 3196 7847 3203 8073
rect 3216 7988 3223 8453
rect 3236 8407 3243 8613
rect 3276 8527 3283 8773
rect 3296 8667 3303 8933
rect 3316 8643 3323 9234
rect 3336 9107 3343 9496
rect 3356 9047 3363 9573
rect 3416 9567 3423 9633
rect 3376 9506 3383 9553
rect 3396 9467 3403 9533
rect 3416 9487 3423 9553
rect 3456 9447 3463 9716
rect 3556 9536 3563 9873
rect 3576 9723 3583 9973
rect 3653 9760 3667 9773
rect 3656 9756 3663 9760
rect 3576 9716 3603 9723
rect 3496 9407 3503 9503
rect 3516 9187 3523 9473
rect 3536 9467 3543 9503
rect 3536 9207 3543 9432
rect 3556 9147 3563 9393
rect 3596 9363 3603 9716
rect 3680 9723 3693 9727
rect 3676 9716 3693 9723
rect 3680 9713 3693 9716
rect 3716 9687 3723 10013
rect 3736 9727 3743 9773
rect 3756 9727 3763 9893
rect 3896 9807 3903 10023
rect 3756 9587 3763 9713
rect 3733 9540 3747 9553
rect 3776 9548 3783 9793
rect 3936 9787 3943 10054
rect 3976 9783 3983 10333
rect 3996 10207 4003 10254
rect 3996 9807 4003 10113
rect 4016 10087 4023 10263
rect 4016 10027 4023 10073
rect 4036 9907 4043 10313
rect 4093 10263 4107 10274
rect 4076 10260 4107 10263
rect 4076 10256 4103 10260
rect 4076 10203 4083 10256
rect 4076 10196 4103 10203
rect 4096 10056 4103 10196
rect 3956 9776 3983 9783
rect 3736 9536 3743 9540
rect 3816 9507 3823 9754
rect 3716 9407 3723 9492
rect 3756 9467 3763 9503
rect 3756 9407 3763 9453
rect 3576 9356 3603 9363
rect 3373 9003 3387 9013
rect 3356 9000 3387 9003
rect 3356 8996 3383 9000
rect 3376 8747 3383 8973
rect 3396 8947 3403 9093
rect 3396 8716 3403 8893
rect 3416 8787 3423 9113
rect 3436 8987 3443 9132
rect 3436 8727 3443 8753
rect 3296 8636 3323 8643
rect 3296 8547 3303 8636
rect 3316 8547 3323 8613
rect 3256 8496 3283 8503
rect 3256 8347 3263 8496
rect 3336 8463 3343 8513
rect 3316 8456 3343 8463
rect 3276 8287 3283 8313
rect 3336 8307 3343 8353
rect 3256 8196 3263 8233
rect 3293 8200 3307 8213
rect 3296 8196 3303 8200
rect 3296 7976 3303 8073
rect 3076 7676 3083 7680
rect 2856 6923 2863 7113
rect 2887 7076 2953 7083
rect 2907 7057 2933 7064
rect 2916 6947 2923 6993
rect 2936 6987 2943 7032
rect 2976 7007 2983 7154
rect 2996 7127 3003 7313
rect 3016 7083 3023 7412
rect 3056 7187 3063 7493
rect 3056 7087 3063 7152
rect 3016 7076 3043 7083
rect 3036 6987 3043 7076
rect 3027 6963 3040 6967
rect 3027 6953 3043 6963
rect 2856 6916 2883 6923
rect 2836 6507 2843 6673
rect 2876 6648 2883 6916
rect 3036 6923 3043 6953
rect 3076 6923 3083 7613
rect 3096 7227 3103 7643
rect 3156 7627 3163 7673
rect 3176 7627 3183 7693
rect 3156 7423 3163 7592
rect 3136 7416 3163 7423
rect 3176 7163 3183 7513
rect 3196 7287 3203 7693
rect 3216 7407 3223 7974
rect 3336 7847 3343 7993
rect 3356 7867 3363 8653
rect 3376 8627 3383 8683
rect 3456 8543 3463 9033
rect 3436 8536 3463 8543
rect 3416 8447 3423 8513
rect 3376 7847 3383 8433
rect 3396 8166 3403 8233
rect 3436 8166 3443 8536
rect 3476 8527 3483 9133
rect 3576 9127 3583 9356
rect 3736 9347 3743 9373
rect 3596 9023 3603 9293
rect 3616 9167 3623 9273
rect 3656 9236 3663 9313
rect 3756 9207 3763 9234
rect 3596 9016 3623 9023
rect 3496 8787 3503 8853
rect 3496 8643 3503 8733
rect 3516 8667 3523 9013
rect 3616 8986 3623 9016
rect 3536 8687 3543 8733
rect 3496 8636 3523 8643
rect 3456 8466 3463 8513
rect 3516 8496 3523 8636
rect 3556 8527 3563 8933
rect 3576 8827 3583 8913
rect 3636 8887 3643 9193
rect 3676 9187 3683 9203
rect 3716 9183 3723 9192
rect 3716 9176 3743 9183
rect 3673 9167 3687 9173
rect 3596 8767 3603 8833
rect 3596 8716 3603 8753
rect 3656 8747 3663 9113
rect 3676 8967 3683 9073
rect 3696 8947 3703 9033
rect 3676 8867 3683 8913
rect 3676 8716 3683 8853
rect 3656 8680 3663 8683
rect 3653 8667 3667 8680
rect 3716 8647 3723 9153
rect 3736 9028 3743 9176
rect 3776 9127 3783 9333
rect 3796 9187 3803 9313
rect 3816 9247 3823 9493
rect 3836 9407 3843 9713
rect 3876 9647 3883 9723
rect 3916 9720 3923 9723
rect 3913 9707 3927 9720
rect 3956 9647 3963 9776
rect 3976 9707 3983 9753
rect 3976 9587 3983 9693
rect 3836 9347 3843 9393
rect 3836 9047 3843 9333
rect 3773 9020 3787 9033
rect 3776 9016 3783 9020
rect 3856 9023 3863 9533
rect 3876 9347 3883 9473
rect 3916 9387 3923 9573
rect 3956 9500 3963 9503
rect 3996 9500 4003 9503
rect 3953 9487 3967 9500
rect 3993 9487 4007 9500
rect 3916 9236 3923 9273
rect 3976 9243 3983 9473
rect 3956 9236 3983 9243
rect 3896 9127 3903 9203
rect 3856 9016 3883 9023
rect 3756 8947 3763 8983
rect 3796 8907 3803 8983
rect 3560 8503 3573 8507
rect 3556 8496 3573 8503
rect 3560 8493 3573 8496
rect 3536 8460 3543 8463
rect 3236 7647 3243 7833
rect 3256 7667 3263 7793
rect 3316 7707 3323 7833
rect 3416 7703 3423 8113
rect 3456 8027 3463 8452
rect 3533 8447 3547 8460
rect 3553 8200 3567 8213
rect 3556 8196 3563 8200
rect 3496 8127 3503 8152
rect 3496 7976 3503 8053
rect 3536 7976 3543 8013
rect 3476 7847 3483 7943
rect 3596 7907 3603 8473
rect 3616 8167 3623 8373
rect 3636 8067 3643 8633
rect 3736 8627 3743 8873
rect 3733 8500 3747 8513
rect 3776 8508 3783 8873
rect 3876 8827 3883 9016
rect 3896 8947 3903 9013
rect 3916 8887 3923 9173
rect 3936 9147 3943 9203
rect 4016 9107 4023 9313
rect 4036 9107 4043 9853
rect 4056 9287 4063 10013
rect 4076 9767 4083 10023
rect 4136 9987 4143 10054
rect 4156 9967 4163 10333
rect 4116 9756 4123 9873
rect 4176 9727 4183 10153
rect 4196 9647 4203 10532
rect 4256 10327 4263 10543
rect 4476 10527 4483 10543
rect 4596 10527 4603 10553
rect 4316 10276 4323 10373
rect 4356 10247 4363 10274
rect 4376 10147 4383 10313
rect 4436 10207 4443 10393
rect 4456 10307 4463 10373
rect 4476 10327 4483 10513
rect 4516 10276 4523 10333
rect 4496 10240 4503 10243
rect 4493 10227 4507 10240
rect 4256 10027 4263 10133
rect 4396 10036 4403 10193
rect 3796 8687 3803 8733
rect 3736 8496 3743 8500
rect 3816 8507 3823 8813
rect 3956 8803 3963 9093
rect 4056 9027 4063 9252
rect 4036 8980 4043 8983
rect 4033 8967 4047 8980
rect 3936 8796 3963 8803
rect 3856 8716 3863 8773
rect 3936 8727 3943 8796
rect 4076 8748 4083 9533
rect 4096 8967 4103 9473
rect 4116 9247 4123 9473
rect 4136 9268 4143 9633
rect 4176 9536 4183 9573
rect 4216 9536 4223 9573
rect 4236 9563 4243 9933
rect 4256 9707 4263 9793
rect 4336 9756 4343 9853
rect 4276 9567 4283 9713
rect 4356 9720 4363 9723
rect 4353 9707 4367 9720
rect 4396 9687 4403 9953
rect 4416 9647 4423 10193
rect 4536 10147 4543 10243
rect 4616 10207 4623 10613
rect 4676 10576 4683 10733
rect 4756 10543 4763 10736
rect 4696 10540 4703 10543
rect 4693 10527 4707 10540
rect 4736 10536 4763 10543
rect 4516 9947 4523 10043
rect 4236 9556 4263 9563
rect 4256 9548 4263 9556
rect 4196 9500 4203 9503
rect 4193 9487 4207 9500
rect 4196 9447 4203 9473
rect 4276 9407 4283 9492
rect 4176 9236 4183 9333
rect 4236 9206 4243 9253
rect 4116 8987 4123 9193
rect 3696 8267 3703 8493
rect 3836 8467 3843 8533
rect 3756 8367 3763 8463
rect 3796 8327 3803 8463
rect 3813 8287 3827 8293
rect 3676 8143 3683 8213
rect 3696 8166 3703 8253
rect 3836 8247 3843 8333
rect 3800 8203 3813 8207
rect 3796 8196 3813 8203
rect 3800 8193 3813 8196
rect 3676 8136 3703 8143
rect 3696 7983 3703 8136
rect 3716 8047 3723 8073
rect 3727 7993 3733 8007
rect 3696 7976 3723 7983
rect 3756 7976 3763 8033
rect 3776 8007 3783 8163
rect 3856 8067 3863 8493
rect 3876 8487 3883 8613
rect 3896 8287 3903 8653
rect 3916 8627 3923 8683
rect 3956 8667 3963 8714
rect 3976 8547 3983 8593
rect 3996 8587 4003 8713
rect 4016 8627 4023 8733
rect 4156 8727 4163 8972
rect 4016 8528 4023 8613
rect 4036 8567 4043 8713
rect 4096 8680 4103 8683
rect 4093 8667 4107 8680
rect 4036 8556 4053 8567
rect 4040 8553 4053 8556
rect 3916 8427 3923 8494
rect 3947 8463 3960 8467
rect 3947 8456 3963 8463
rect 3947 8453 3960 8456
rect 3927 8293 3933 8307
rect 3896 8227 3903 8273
rect 3996 8228 4003 8463
rect 3776 7936 3803 7943
rect 3476 7807 3483 7833
rect 3407 7696 3423 7703
rect 3316 7676 3323 7693
rect 3353 7680 3367 7693
rect 3356 7676 3363 7680
rect 3156 7156 3203 7163
rect 3196 7126 3203 7156
rect 3136 7087 3143 7123
rect 3136 7047 3143 7073
rect 3216 7067 3223 7193
rect 3236 7067 3243 7453
rect 3276 7426 3283 7613
rect 3296 7587 3303 7643
rect 3436 7527 3443 7613
rect 3456 7503 3463 7694
rect 3696 7663 3703 7932
rect 3756 7867 3763 7913
rect 3796 7827 3803 7936
rect 3816 7927 3823 8033
rect 3696 7656 3723 7663
rect 3436 7496 3463 7503
rect 3296 7407 3303 7454
rect 3356 7387 3363 7423
rect 3396 7267 3403 7333
rect 3396 7156 3403 7253
rect 3196 7027 3203 7053
rect 3313 7047 3327 7053
rect 3336 6947 3343 6993
rect 3376 6947 3383 6973
rect 3036 6916 3063 6923
rect 3076 6916 3103 6923
rect 2936 6887 2943 6903
rect 2916 6707 2923 6753
rect 2936 6643 2943 6873
rect 2916 6636 2943 6643
rect 2756 6436 2783 6443
rect 2596 6347 2603 6383
rect 2756 6367 2763 6414
rect 2776 6367 2783 6436
rect 2796 6407 2803 6433
rect 2876 6416 2883 6493
rect 2896 6487 2903 6603
rect 2916 6416 2923 6573
rect 2956 6427 2963 6634
rect 2976 6606 2983 6893
rect 2560 6346 2580 6347
rect 2567 6343 2580 6346
rect 2567 6336 2593 6343
rect 2567 6333 2580 6336
rect 2476 6096 2503 6103
rect 2536 6100 2543 6103
rect 2533 6087 2547 6100
rect 2536 6027 2543 6073
rect 2336 5596 2343 5693
rect 2456 5687 2463 5733
rect 2056 5346 2063 5473
rect 2113 5327 2127 5332
rect 2116 5187 2123 5273
rect 2136 5167 2143 5293
rect 2156 5187 2163 5332
rect 2196 5307 2203 5374
rect 1936 4747 1943 4773
rect 1976 4667 1983 4773
rect 1936 4587 1943 4653
rect 1956 3947 1963 4613
rect 1996 4607 2003 4873
rect 2016 4767 2023 5093
rect 2053 5080 2067 5093
rect 2056 5076 2063 5080
rect 2096 5076 2103 5113
rect 2196 5047 2203 5272
rect 2216 5247 2223 5453
rect 2236 5447 2243 5594
rect 2316 5560 2323 5563
rect 2313 5547 2327 5560
rect 2247 5436 2263 5443
rect 2256 5307 2263 5436
rect 2276 5307 2283 5473
rect 2236 5267 2243 5293
rect 2296 5287 2303 5393
rect 2313 5387 2327 5393
rect 2356 5376 2363 5413
rect 2396 5376 2403 5473
rect 2413 5387 2427 5393
rect 2336 5307 2343 5343
rect 2376 5340 2383 5343
rect 2373 5327 2387 5340
rect 2216 5067 2223 5193
rect 2256 5187 2263 5233
rect 2036 4703 2043 5033
rect 2176 5036 2193 5043
rect 2067 5023 2080 5027
rect 2067 5020 2083 5023
rect 2067 5013 2087 5020
rect 2073 5007 2087 5013
rect 2136 4856 2143 4913
rect 2176 4887 2183 5036
rect 2076 4787 2083 4823
rect 2036 4696 2063 4703
rect 2033 4603 2047 4613
rect 2056 4607 2063 4696
rect 2076 4667 2083 4773
rect 2016 4600 2047 4603
rect 2016 4596 2043 4600
rect 2016 4587 2023 4596
rect 2013 4560 2027 4573
rect 2016 4556 2023 4560
rect 1996 4327 2003 4512
rect 2036 4487 2043 4523
rect 2076 4348 2083 4393
rect 2096 4367 2103 4593
rect 2116 4336 2123 4753
rect 2136 4727 2143 4793
rect 2136 4487 2143 4692
rect 2016 4267 2023 4334
rect 2056 4207 2063 4303
rect 1867 3573 1873 3587
rect 1913 3567 1927 3573
rect 1856 3387 1863 3433
rect 1836 3356 1863 3363
rect 1636 3267 1643 3293
rect 1716 3260 1723 3263
rect 1776 3260 1783 3263
rect 1713 3247 1727 3260
rect 1773 3247 1787 3260
rect 1636 3047 1643 3213
rect 1636 2966 1643 3033
rect 1476 2447 1483 2533
rect 1496 2487 1503 2893
rect 1556 2776 1563 2893
rect 1636 2747 1643 2774
rect 1536 2476 1543 2513
rect 1576 2508 1583 2743
rect 1616 2487 1623 2533
rect 1496 2327 1503 2473
rect 1636 2443 1643 2513
rect 1616 2436 1643 2443
rect 1556 2256 1563 2293
rect 1476 1987 1483 2093
rect 1536 2027 1543 2223
rect 1616 2167 1623 2436
rect 1496 1956 1503 2013
rect 1516 1887 1523 1923
rect 1456 1748 1463 1813
rect 1496 1700 1503 1703
rect 1493 1687 1507 1700
rect 1496 1436 1503 1473
rect 1536 1427 1543 1692
rect 1436 1356 1453 1363
rect 1456 1267 1463 1353
rect 1456 1183 1463 1253
rect 1516 1216 1523 1273
rect 1456 1176 1483 1183
rect 1413 920 1427 933
rect 1456 928 1463 1013
rect 1476 947 1483 1176
rect 1416 916 1423 920
rect 1436 723 1443 883
rect 1476 847 1483 872
rect 1436 716 1463 723
rect 1333 700 1347 713
rect 1336 696 1343 700
rect 1436 567 1443 693
rect 1456 666 1463 716
rect 1476 667 1483 713
rect 1536 627 1543 1413
rect 1556 1406 1563 1553
rect 1576 1327 1583 1573
rect 1596 1487 1603 1993
rect 1596 1167 1603 1313
rect 1616 1127 1623 2153
rect 1636 1627 1643 2273
rect 1656 2227 1663 3193
rect 1676 3007 1683 3173
rect 1716 3008 1723 3133
rect 1756 2996 1763 3093
rect 1796 3067 1803 3273
rect 1816 3147 1823 3313
rect 1836 3187 1843 3253
rect 1676 2547 1683 2893
rect 1736 2847 1743 2963
rect 1736 2767 1743 2833
rect 1796 2776 1803 3032
rect 1816 2967 1823 3093
rect 1836 2947 1843 3053
rect 1816 2723 1823 2743
rect 1796 2716 1823 2723
rect 1796 2627 1803 2716
rect 1796 2567 1803 2613
rect 1716 2268 1723 2493
rect 1776 2476 1783 2533
rect 1856 2507 1863 3356
rect 1876 3307 1883 3552
rect 1896 3283 1903 3533
rect 1916 3487 1923 3514
rect 1936 3467 1943 3633
rect 1976 3547 1983 4073
rect 2056 4036 2063 4193
rect 1996 3907 2003 3992
rect 1996 3528 2003 3893
rect 2056 3727 2063 3783
rect 1913 3367 1927 3373
rect 1876 3276 1903 3283
rect 1876 3207 1883 3276
rect 1916 3267 1923 3332
rect 1876 2746 1883 2993
rect 1756 2407 1763 2443
rect 1796 2423 1803 2443
rect 1796 2416 1823 2423
rect 1816 2267 1823 2416
rect 1836 2268 1843 2313
rect 1836 2223 1843 2254
rect 1776 2207 1783 2223
rect 1816 2216 1843 2223
rect 1776 2196 1793 2207
rect 1780 2193 1793 2196
rect 1696 1907 1703 2013
rect 1796 1968 1803 2153
rect 1816 2027 1823 2216
rect 1756 1956 1783 1963
rect 1696 1736 1703 1893
rect 1716 1748 1723 1923
rect 1776 1787 1783 1956
rect 1816 1847 1823 1954
rect 1836 1807 1843 2153
rect 1856 2047 1863 2493
rect 1876 2447 1883 2732
rect 1876 2307 1883 2412
rect 1856 1783 1863 2012
rect 1876 1947 1883 2133
rect 1896 2107 1903 3213
rect 1916 3047 1923 3232
rect 1936 3107 1943 3432
rect 1956 3307 1963 3353
rect 1976 3347 1983 3483
rect 1996 3296 2003 3453
rect 2016 3327 2023 3483
rect 2036 3296 2043 3333
rect 2056 3327 2063 3653
rect 2076 3627 2083 3693
rect 2076 3267 2083 3333
rect 1976 3260 1983 3263
rect 1956 3127 1963 3253
rect 1973 3247 1987 3260
rect 1976 3107 1983 3233
rect 2016 3227 2023 3263
rect 2016 3067 2023 3133
rect 1933 3000 1947 3013
rect 1973 3000 1987 3013
rect 1936 2996 1943 3000
rect 1976 2996 1983 3000
rect 1916 2587 1923 2953
rect 1936 2647 1943 2933
rect 1956 2907 1963 2963
rect 2036 2907 2043 3053
rect 1956 2807 1963 2853
rect 2056 2847 2063 2973
rect 2076 2967 2083 3193
rect 2096 2927 2103 3953
rect 1916 2207 1923 2293
rect 1936 2167 1943 2433
rect 1956 2367 1963 2493
rect 1976 2488 1983 2813
rect 2076 2747 2083 2853
rect 1996 2507 2003 2693
rect 2016 2503 2023 2533
rect 2036 2527 2043 2743
rect 2096 2707 2103 2892
rect 2096 2547 2103 2633
rect 2016 2496 2043 2503
rect 1993 2480 2007 2493
rect 1996 2476 2003 2480
rect 2036 2476 2043 2496
rect 2076 2476 2083 2513
rect 2016 2440 2023 2443
rect 2013 2427 2027 2440
rect 1996 2256 2003 2293
rect 2016 2287 2023 2413
rect 1976 2167 1983 2223
rect 1896 2007 1903 2093
rect 1996 2007 2003 2053
rect 1936 1887 1943 1923
rect 1996 1907 2003 1993
rect 2016 1887 2023 2212
rect 2016 1827 2023 1873
rect 1836 1776 1863 1783
rect 1696 1436 1703 1473
rect 1756 1467 1763 1673
rect 1776 1647 1783 1733
rect 1636 1267 1643 1333
rect 1676 1267 1683 1392
rect 1736 1347 1743 1392
rect 1716 1216 1723 1293
rect 1756 1228 1763 1453
rect 1796 1347 1803 1753
rect 1836 1667 1843 1776
rect 1916 1736 1923 1793
rect 2016 1707 2023 1773
rect 1896 1700 1903 1703
rect 1893 1687 1907 1700
rect 1936 1683 1943 1703
rect 1916 1676 1943 1683
rect 1816 1387 1823 1433
rect 1656 1183 1663 1213
rect 1656 1176 1683 1183
rect 1696 1180 1703 1183
rect 1676 1067 1683 1176
rect 1693 1167 1707 1180
rect 1576 886 1583 933
rect 1676 916 1683 1053
rect 1713 928 1727 933
rect 1796 928 1803 1213
rect 1836 1186 1843 1473
rect 1896 1436 1903 1652
rect 1916 1507 1923 1676
rect 1936 1527 1943 1593
rect 2036 1567 2043 2213
rect 2056 2067 2063 2443
rect 2076 2227 2083 2353
rect 2056 1787 2063 1954
rect 2096 1907 2103 2373
rect 2116 2227 2123 4153
rect 2136 4027 2143 4133
rect 2156 4067 2163 4453
rect 2176 4043 2183 4852
rect 2196 4826 2203 4853
rect 2216 4667 2223 4973
rect 2236 4667 2243 5153
rect 2276 4967 2283 5043
rect 2333 4987 2347 4993
rect 2356 4967 2363 5073
rect 2276 4927 2283 4953
rect 2156 4036 2183 4043
rect 2136 3787 2143 3833
rect 2136 2567 2143 3773
rect 2156 3247 2163 4036
rect 2176 3767 2183 3793
rect 2196 3627 2203 4573
rect 2236 4556 2243 4653
rect 2256 4587 2263 4853
rect 2276 4687 2283 4873
rect 2296 4867 2303 4893
rect 2316 4887 2323 4953
rect 2376 4907 2383 5273
rect 2396 4987 2403 5153
rect 2396 4863 2403 4973
rect 2376 4856 2403 4863
rect 2287 4603 2300 4607
rect 2287 4600 2303 4603
rect 2287 4593 2307 4600
rect 2293 4587 2307 4593
rect 2216 4227 2223 4512
rect 2296 4487 2303 4523
rect 2316 4336 2323 4513
rect 2336 4487 2343 4573
rect 2356 4336 2363 4393
rect 2376 4347 2383 4773
rect 2396 4627 2403 4713
rect 2256 4247 2263 4334
rect 2396 4307 2403 4613
rect 2416 4307 2423 5332
rect 2436 5207 2443 5593
rect 2456 5388 2463 5533
rect 2476 5503 2483 5893
rect 2496 5627 2503 6013
rect 2536 5896 2543 5953
rect 2556 5947 2563 6073
rect 2576 5967 2583 5993
rect 2573 5900 2587 5913
rect 2596 5907 2603 6312
rect 2576 5896 2583 5900
rect 2556 5747 2563 5863
rect 2536 5596 2543 5713
rect 2573 5600 2587 5613
rect 2593 5607 2607 5613
rect 2576 5596 2583 5600
rect 2476 5496 2503 5503
rect 2436 5027 2443 5074
rect 2456 5043 2463 5374
rect 2476 5347 2483 5473
rect 2496 5346 2503 5496
rect 2516 5387 2523 5563
rect 2616 5527 2623 6353
rect 2636 5827 2643 6333
rect 2716 6303 2723 6352
rect 2696 6296 2723 6303
rect 2656 6007 2663 6073
rect 2676 6047 2683 6213
rect 2696 6107 2703 6296
rect 2836 6207 2843 6273
rect 2856 6267 2863 6383
rect 2736 6167 2743 6193
rect 2736 6116 2743 6153
rect 2656 5707 2663 5893
rect 2636 5647 2643 5673
rect 2636 5566 2643 5633
rect 2656 5543 2663 5613
rect 2636 5536 2663 5543
rect 2536 5287 2543 5513
rect 2556 5427 2563 5493
rect 2616 5403 2623 5492
rect 2636 5427 2643 5536
rect 2656 5447 2663 5473
rect 2676 5467 2683 6033
rect 2696 5866 2703 6072
rect 2696 5767 2703 5813
rect 2716 5523 2723 6073
rect 2756 5927 2763 6072
rect 2796 6047 2803 6083
rect 2816 5896 2823 5973
rect 2856 5947 2863 6153
rect 2796 5747 2803 5863
rect 2796 5687 2803 5733
rect 2773 5600 2787 5613
rect 2816 5608 2823 5653
rect 2776 5596 2783 5600
rect 2716 5516 2743 5523
rect 2616 5396 2643 5403
rect 2636 5376 2643 5396
rect 2736 5388 2743 5516
rect 2756 5487 2763 5563
rect 2756 5347 2763 5473
rect 2793 5447 2807 5453
rect 2856 5447 2863 5473
rect 2656 5307 2663 5332
rect 2576 5187 2583 5233
rect 2553 5107 2567 5113
rect 2487 5083 2500 5087
rect 2487 5076 2503 5083
rect 2487 5073 2500 5076
rect 2576 5087 2583 5133
rect 2596 5127 2603 5213
rect 2456 5036 2483 5043
rect 2436 4826 2443 4953
rect 2433 4807 2447 4812
rect 2456 4667 2463 5013
rect 2476 4747 2483 5036
rect 2496 4727 2503 5013
rect 2556 4987 2563 5043
rect 2616 4987 2623 5133
rect 2656 5087 2663 5233
rect 2676 5187 2683 5233
rect 2716 5107 2723 5213
rect 2776 5087 2783 5233
rect 2676 4987 2683 5073
rect 2756 5023 2763 5032
rect 2736 5016 2763 5023
rect 2556 4888 2563 4973
rect 2596 4856 2603 4913
rect 2516 4787 2523 4853
rect 2496 4587 2503 4633
rect 2516 4556 2523 4733
rect 2296 4283 2303 4303
rect 2296 4276 2323 4283
rect 2236 3967 2243 4213
rect 2256 4187 2263 4212
rect 2256 3816 2263 4173
rect 2316 4147 2323 4276
rect 2316 4036 2323 4133
rect 2336 4087 2343 4303
rect 2376 4207 2383 4293
rect 2436 4287 2443 4554
rect 2456 4516 2483 4523
rect 2276 3907 2283 4003
rect 2236 3780 2243 3783
rect 2276 3780 2283 3783
rect 2233 3767 2247 3780
rect 2273 3767 2287 3780
rect 2216 3667 2223 3753
rect 2176 3347 2183 3593
rect 2253 3567 2267 3573
rect 2216 3296 2223 3453
rect 2196 3147 2203 3263
rect 2216 3167 2223 3213
rect 2236 3207 2243 3263
rect 2276 3167 2283 3513
rect 2153 3027 2167 3033
rect 2256 3027 2263 3093
rect 2193 3000 2207 3013
rect 2240 3006 2260 3007
rect 2240 3003 2253 3006
rect 2196 2996 2203 3000
rect 2236 2996 2253 3003
rect 2240 2993 2253 2996
rect 2156 2627 2163 2953
rect 2176 2727 2183 2952
rect 2216 2927 2223 2963
rect 2276 2788 2283 3132
rect 2296 3067 2303 3773
rect 2316 3767 2323 3873
rect 2336 3767 2343 4052
rect 2316 3467 2323 3732
rect 2316 3266 2323 3313
rect 2336 3263 2343 3633
rect 2356 3367 2363 4093
rect 2376 3787 2383 4193
rect 2396 3947 2403 4253
rect 2376 3483 2383 3752
rect 2396 3567 2403 3933
rect 2416 3807 2423 4073
rect 2436 3947 2443 4013
rect 2456 4007 2463 4516
rect 2476 4047 2483 4473
rect 2536 4427 2543 4793
rect 2573 4787 2587 4791
rect 2556 4487 2563 4653
rect 2596 4367 2603 4673
rect 2616 4627 2623 4823
rect 2636 4727 2643 4812
rect 2636 4527 2643 4554
rect 2636 4487 2643 4513
rect 2556 4300 2563 4303
rect 2516 4267 2523 4293
rect 2553 4287 2567 4300
rect 2496 4036 2503 4133
rect 2536 4036 2543 4093
rect 2456 3967 2463 3993
rect 2496 3867 2503 3893
rect 2513 3820 2527 3833
rect 2536 3827 2543 3853
rect 2516 3816 2523 3820
rect 2456 3747 2463 3783
rect 2416 3516 2423 3693
rect 2496 3667 2503 3783
rect 2556 3767 2563 3953
rect 2576 3787 2583 3833
rect 2516 3647 2523 3753
rect 2500 3646 2523 3647
rect 2507 3636 2523 3646
rect 2507 3633 2520 3636
rect 2456 3528 2463 3553
rect 2493 3528 2507 3533
rect 2376 3476 2403 3483
rect 2327 3256 2343 3263
rect 2316 3187 2323 3213
rect 2336 3047 2343 3153
rect 2316 2966 2323 2993
rect 2296 2907 2303 2953
rect 2136 2187 2143 2513
rect 2156 2226 2163 2613
rect 2176 2267 2183 2573
rect 2196 2327 2203 2533
rect 2216 2387 2223 2553
rect 2256 2547 2263 2733
rect 2253 2480 2267 2493
rect 2256 2476 2263 2480
rect 2296 2476 2303 2853
rect 2316 2483 2323 2952
rect 2336 2907 2343 3012
rect 2356 3007 2363 3294
rect 2376 3087 2383 3333
rect 2396 3327 2403 3476
rect 2436 3347 2443 3472
rect 2476 3427 2483 3483
rect 2433 3300 2447 3312
rect 2436 3296 2443 3300
rect 2416 3127 2423 3263
rect 2356 2967 2363 2993
rect 2356 2746 2363 2793
rect 2336 2587 2343 2653
rect 2316 2476 2333 2483
rect 2216 2256 2223 2352
rect 2236 2187 2243 2223
rect 2156 1956 2163 2033
rect 2256 1967 2263 2193
rect 2276 2047 2283 2253
rect 2136 1920 2143 1923
rect 2133 1907 2147 1920
rect 2136 1807 2143 1893
rect 2176 1887 2183 1923
rect 2276 1867 2283 2033
rect 2296 2027 2303 2173
rect 2176 1736 2183 1833
rect 2056 1687 2063 1733
rect 2107 1703 2120 1707
rect 2107 1696 2123 1703
rect 2156 1700 2163 1703
rect 2107 1693 2120 1696
rect 2153 1687 2167 1700
rect 1976 1427 1983 1493
rect 2116 1436 2123 1553
rect 2153 1440 2167 1453
rect 2156 1436 2163 1440
rect 2216 1406 2223 1793
rect 2236 1748 2243 1793
rect 2247 1736 2263 1743
rect 1856 1228 1863 1373
rect 1993 1287 2007 1293
rect 1896 1186 1903 1253
rect 1956 1147 1963 1183
rect 2056 1167 2063 1353
rect 2096 1228 2103 1392
rect 2136 1327 2143 1403
rect 2133 1287 2147 1292
rect 2116 1216 2163 1223
rect 1816 1027 1823 1073
rect 1576 696 1583 872
rect 1596 627 1603 663
rect 1596 587 1603 613
rect 1296 396 1323 403
rect 933 160 947 173
rect 1216 166 1223 253
rect 936 156 943 160
rect 1236 156 1243 333
rect 1256 287 1263 363
rect 1316 307 1323 396
rect 1336 327 1343 383
rect 1256 168 1263 273
rect 1396 168 1403 383
rect 1576 376 1583 453
rect 1736 428 1743 833
rect 1796 827 1803 914
rect 1836 887 1843 914
rect 1856 887 1863 1013
rect 1896 1007 1903 1033
rect 1956 827 1963 883
rect 1836 696 1843 733
rect 1873 700 1887 713
rect 1876 696 1883 700
rect 1776 627 1783 693
rect 1956 666 1963 813
rect 2016 666 2023 733
rect 2096 727 2103 1214
rect 2116 1147 2123 1216
rect 2116 1007 2123 1133
rect 2176 1127 2183 1183
rect 2216 1087 2223 1133
rect 2236 967 2243 1214
rect 2256 886 2263 1736
rect 2276 1047 2283 1853
rect 2316 1807 2323 2433
rect 2336 1987 2343 2474
rect 2356 2287 2363 2693
rect 2376 2667 2383 3052
rect 2393 3027 2407 3033
rect 2396 3007 2403 3013
rect 2416 2996 2423 3053
rect 2456 2996 2463 3073
rect 2496 3027 2503 3053
rect 2476 2827 2483 2952
rect 2496 2803 2503 2953
rect 2433 2780 2447 2793
rect 2476 2796 2503 2803
rect 2436 2776 2443 2780
rect 2476 2776 2483 2796
rect 2376 2347 2383 2653
rect 2416 2287 2423 2732
rect 2456 2547 2463 2743
rect 2516 2607 2523 3613
rect 2536 3087 2543 3553
rect 2556 3147 2563 3753
rect 2596 3707 2603 4303
rect 2616 3747 2623 4273
rect 2636 3743 2643 3793
rect 2656 3767 2663 4953
rect 2736 4927 2743 5016
rect 2676 4556 2683 4913
rect 2676 4067 2683 4353
rect 2696 4047 2703 4512
rect 2716 4307 2723 4393
rect 2756 4387 2763 4973
rect 2776 4927 2783 5033
rect 2796 4947 2803 5333
rect 2816 5047 2823 5293
rect 2836 5027 2843 5332
rect 2856 5047 2863 5193
rect 2836 4967 2843 5013
rect 2776 4823 2783 4873
rect 2776 4816 2803 4823
rect 2816 4547 2823 4773
rect 2776 4127 2783 4303
rect 2753 4040 2767 4053
rect 2756 4036 2763 4040
rect 2676 3987 2683 4032
rect 2780 4004 2793 4007
rect 2736 3867 2743 4003
rect 2776 3997 2793 4004
rect 2780 3993 2793 3997
rect 2693 3828 2707 3833
rect 2733 3820 2747 3832
rect 2736 3816 2743 3820
rect 2716 3767 2723 3783
rect 2707 3756 2723 3767
rect 2707 3753 2720 3756
rect 2636 3736 2663 3743
rect 2607 3696 2623 3703
rect 2576 3587 2583 3653
rect 2576 3487 2583 3533
rect 2596 3247 2603 3653
rect 2616 3527 2623 3696
rect 2636 3627 2643 3713
rect 2656 3707 2663 3736
rect 2647 3540 2683 3543
rect 2647 3536 2687 3540
rect 2673 3527 2687 3536
rect 2716 3427 2723 3453
rect 2676 3296 2683 3373
rect 2716 3307 2723 3353
rect 2736 3266 2743 3753
rect 2756 3447 2763 3773
rect 2576 3167 2583 3233
rect 2556 2807 2563 3053
rect 2576 3007 2583 3053
rect 2616 2967 2623 3193
rect 2633 3067 2647 3073
rect 2656 2996 2663 3231
rect 2696 3027 2703 3263
rect 2636 2967 2643 2994
rect 2676 2960 2683 2963
rect 2673 2947 2687 2960
rect 2536 2667 2543 2713
rect 2556 2527 2563 2793
rect 2596 2707 2603 2793
rect 2616 2767 2623 2932
rect 2653 2788 2667 2793
rect 2516 2476 2523 2513
rect 2376 2226 2383 2273
rect 2436 2256 2443 2313
rect 2496 2287 2503 2443
rect 2556 2327 2563 2513
rect 2456 2220 2463 2223
rect 2453 2207 2467 2220
rect 2373 1960 2387 1973
rect 2416 1968 2423 2013
rect 2376 1956 2383 1960
rect 2396 1920 2403 1923
rect 2393 1907 2407 1920
rect 2456 1867 2463 1993
rect 2296 1483 2303 1653
rect 2316 1507 2323 1734
rect 2456 1706 2463 1793
rect 2296 1476 2323 1483
rect 2316 1436 2323 1476
rect 2416 1447 2423 1703
rect 2336 1167 2343 1403
rect 2436 1267 2443 1434
rect 2436 1216 2443 1253
rect 2476 1187 2483 2133
rect 2376 1180 2383 1183
rect 2373 1167 2387 1180
rect 2356 916 2363 953
rect 2336 867 2343 883
rect 2336 856 2353 867
rect 2340 853 2353 856
rect 2116 696 2123 813
rect 2293 700 2307 713
rect 2296 696 2303 700
rect 2336 696 2343 793
rect 1856 587 1863 663
rect 1816 387 1823 513
rect 1276 87 1283 123
rect 1576 67 1583 163
rect 1696 156 1703 213
rect 1836 163 1843 413
rect 1936 396 1943 453
rect 2193 400 2207 413
rect 2196 396 2203 400
rect 2216 366 2223 693
rect 2376 627 2383 883
rect 2436 867 2443 913
rect 1956 327 1963 363
rect 1836 156 1863 163
rect 1736 87 1743 123
rect 1856 87 1863 156
rect 1956 87 1963 163
rect 2096 127 2103 213
rect 2196 156 2203 293
rect 2296 227 2303 513
rect 2336 366 2343 433
rect 2376 396 2383 613
rect 2396 587 2403 693
rect 2396 427 2403 573
rect 2456 507 2463 793
rect 2496 703 2503 1833
rect 2516 1547 2523 1633
rect 2536 1487 2543 2293
rect 2576 2087 2583 2474
rect 2616 2327 2623 2613
rect 2636 2447 2643 2493
rect 2613 2307 2627 2313
rect 2656 2287 2663 2533
rect 2676 2527 2683 2743
rect 2736 2567 2743 3252
rect 2756 3247 2763 3433
rect 2776 3367 2783 3873
rect 2753 3067 2767 3073
rect 2756 2747 2763 3013
rect 2776 2966 2783 3293
rect 2796 2707 2803 3972
rect 2816 3727 2823 3793
rect 2836 3747 2843 4793
rect 2856 4227 2863 4913
rect 2876 4247 2883 6353
rect 2896 6147 2903 6333
rect 2936 6187 2943 6383
rect 2896 6067 2903 6093
rect 2936 6086 2943 6113
rect 2896 6007 2903 6053
rect 2896 5567 2903 5873
rect 2916 5747 2923 5933
rect 2896 5007 2903 5473
rect 2936 5347 2943 5833
rect 2956 5427 2963 6373
rect 2976 6127 2983 6493
rect 2996 6407 3003 6473
rect 3036 6467 3043 6916
rect 3016 6387 3023 6413
rect 3016 6167 3023 6233
rect 3016 6116 3023 6153
rect 3036 6127 3043 6413
rect 3056 6407 3063 6833
rect 3096 6767 3103 6916
rect 3336 6916 3363 6923
rect 3336 6767 3343 6916
rect 3396 6827 3403 6883
rect 3436 6827 3443 7496
rect 3473 7483 3487 7493
rect 3456 7480 3487 7483
rect 3456 7476 3483 7480
rect 3456 7207 3463 7476
rect 3456 7107 3463 7154
rect 3307 6753 3313 6767
rect 3073 6707 3087 6713
rect 3156 6647 3163 6693
rect 3136 6567 3143 6603
rect 3153 6527 3167 6533
rect 3176 6507 3183 6693
rect 3236 6648 3243 6753
rect 3196 6487 3203 6633
rect 3276 6607 3283 6733
rect 3307 6643 3320 6647
rect 3307 6636 3323 6643
rect 3307 6633 3320 6636
rect 3416 6606 3423 6673
rect 3336 6567 3343 6603
rect 3326 6553 3327 6560
rect 3287 6533 3293 6547
rect 3313 6543 3327 6553
rect 3313 6540 3343 6543
rect 3316 6536 3343 6540
rect 3056 6227 3063 6293
rect 2996 6080 3003 6083
rect 2993 6067 3007 6080
rect 3076 5987 3083 6414
rect 3096 6167 3103 6373
rect 3136 6363 3143 6383
rect 3136 6356 3163 6363
rect 3156 6267 3163 6356
rect 3176 6347 3183 6383
rect 3136 6086 3143 6153
rect 3156 6083 3163 6253
rect 3236 6187 3243 6473
rect 3256 6116 3263 6153
rect 3156 6076 3183 6083
rect 2976 5807 2983 5973
rect 3116 5896 3123 5933
rect 2996 5866 3003 5893
rect 3016 5827 3023 5863
rect 3056 5596 3063 5673
rect 2996 5447 3003 5563
rect 3116 5407 3123 5833
rect 3136 5567 3143 5853
rect 3156 5847 3163 5894
rect 3013 5380 3027 5393
rect 3016 5376 3023 5380
rect 2976 5307 2983 5353
rect 3036 5323 3043 5343
rect 3036 5316 3063 5323
rect 3016 5167 3023 5273
rect 3036 5227 3043 5293
rect 3056 5107 3063 5316
rect 3076 5247 3083 5343
rect 3096 5223 3103 5333
rect 3156 5287 3163 5613
rect 3176 5347 3183 6076
rect 3236 5947 3243 6083
rect 3236 5867 3243 5894
rect 3256 5596 3263 5753
rect 3276 5627 3283 6072
rect 3296 5967 3303 6293
rect 3316 6067 3323 6333
rect 3336 6027 3343 6536
rect 3376 6167 3383 6383
rect 3336 5896 3343 5992
rect 3376 5987 3383 6132
rect 3316 5687 3323 5863
rect 3356 5767 3363 5863
rect 3396 5847 3403 6353
rect 3436 6147 3443 6792
rect 3456 6307 3463 6933
rect 3476 6267 3483 7393
rect 3496 7367 3503 7553
rect 3696 7547 3703 7633
rect 3456 6116 3463 6153
rect 3496 6123 3503 7213
rect 3516 7127 3523 7193
rect 3536 7107 3543 7412
rect 3576 7387 3583 7423
rect 3716 7423 3723 7656
rect 3736 7607 3743 7663
rect 3756 7587 3763 7773
rect 3776 7456 3783 7513
rect 3796 7487 3803 7553
rect 3816 7507 3823 7892
rect 3836 7867 3843 7993
rect 3856 7967 3863 8013
rect 3816 7456 3823 7493
rect 3716 7416 3743 7423
rect 3596 7156 3603 7413
rect 3516 6787 3523 7092
rect 3536 6863 3543 7013
rect 3556 7007 3563 7073
rect 3576 7027 3583 7123
rect 3616 6987 3623 7123
rect 3656 7120 3663 7123
rect 3653 7107 3667 7120
rect 3656 6936 3663 7013
rect 3556 6883 3563 6933
rect 3596 6887 3603 6903
rect 3556 6876 3583 6883
rect 3536 6856 3563 6863
rect 3516 6747 3523 6773
rect 3536 6767 3543 6813
rect 3556 6636 3563 6856
rect 3576 6707 3583 6876
rect 3596 6807 3603 6873
rect 3636 6847 3643 6903
rect 3536 6567 3543 6603
rect 3496 6116 3523 6123
rect 3196 5307 3203 5594
rect 3216 5327 3223 5513
rect 3236 5407 3243 5563
rect 3276 5556 3303 5563
rect 3276 5376 3283 5533
rect 3296 5527 3303 5556
rect 3316 5547 3323 5613
rect 3236 5336 3263 5343
rect 3193 5287 3207 5293
rect 3076 5216 3103 5223
rect 2960 5103 2973 5107
rect 2956 5093 2973 5103
rect 2956 5076 2963 5093
rect 2936 5040 2943 5043
rect 2933 5027 2947 5040
rect 2916 4868 2923 4893
rect 2933 4787 2947 4793
rect 2956 4747 2963 4854
rect 2976 4807 2983 5043
rect 3036 4987 3043 5073
rect 3076 4856 3083 5216
rect 3116 5103 3123 5233
rect 3096 5096 3123 5103
rect 3096 5046 3103 5096
rect 3193 5080 3207 5093
rect 3236 5087 3243 5336
rect 3296 5323 3303 5343
rect 3276 5316 3303 5323
rect 3196 5076 3203 5080
rect 2956 4667 2963 4733
rect 2976 4587 2983 4713
rect 3016 4587 3023 4823
rect 3056 4747 3063 4823
rect 3076 4687 3083 4793
rect 2940 4583 2953 4587
rect 2936 4573 2953 4583
rect 2936 4556 2943 4573
rect 2896 4227 2903 4413
rect 2916 4347 2923 4523
rect 3056 4487 3063 4613
rect 2916 4287 2923 4312
rect 2876 3887 2883 4013
rect 2916 3987 2923 4273
rect 2936 4267 2943 4373
rect 2956 4347 2963 4473
rect 3076 4407 3083 4673
rect 3116 4627 3123 5074
rect 3216 5040 3223 5043
rect 3213 5027 3227 5040
rect 3236 5003 3243 5033
rect 3216 4996 3243 5003
rect 3156 4807 3163 4833
rect 3176 4787 3183 4993
rect 3113 4560 3127 4573
rect 3116 4556 3123 4560
rect 2976 4300 2983 4303
rect 2973 4287 2987 4300
rect 3033 4267 3047 4273
rect 3056 4227 3063 4292
rect 3013 4047 3027 4053
rect 3036 4007 3043 4033
rect 2933 3987 2947 3992
rect 2956 3907 2963 4003
rect 2856 3787 2863 3853
rect 2876 3776 2903 3783
rect 2876 3707 2883 3776
rect 2856 3447 2863 3483
rect 2896 3407 2903 3733
rect 2936 3647 2943 3783
rect 2920 3626 2940 3627
rect 2927 3613 2933 3626
rect 2956 3463 2963 3673
rect 2976 3487 2983 3973
rect 2996 3687 3003 3893
rect 3013 3727 3027 3733
rect 3036 3727 3043 3813
rect 3056 3767 3063 4213
rect 3076 4087 3083 4334
rect 3096 4127 3103 4193
rect 3116 4127 3123 4473
rect 3136 4087 3143 4523
rect 3196 4507 3203 4953
rect 3216 4567 3223 4996
rect 3256 4967 3263 5313
rect 3276 5247 3283 5316
rect 3276 5127 3283 5233
rect 3296 5007 3303 5173
rect 3316 5027 3323 5313
rect 3256 4787 3263 4823
rect 3236 4543 3243 4573
rect 3216 4536 3243 4543
rect 3156 4287 3163 4493
rect 3176 4207 3183 4393
rect 3216 4348 3223 4536
rect 3256 4336 3263 4554
rect 3276 4547 3283 4673
rect 3296 4523 3303 4813
rect 3316 4787 3323 4873
rect 3336 4827 3343 5273
rect 3356 5147 3363 5374
rect 3356 4727 3363 4873
rect 3376 4807 3383 5773
rect 3396 5567 3403 5812
rect 3396 5487 3403 5553
rect 3416 5327 3423 5973
rect 3436 5263 3443 6051
rect 3456 5827 3463 6013
rect 3476 5947 3483 6083
rect 3476 5887 3483 5933
rect 3496 5596 3503 6073
rect 3516 5967 3523 6116
rect 3536 6087 3543 6433
rect 3573 6420 3587 6433
rect 3576 6416 3583 6420
rect 3616 6416 3623 6813
rect 3596 6263 3603 6383
rect 3636 6380 3643 6383
rect 3633 6367 3647 6380
rect 3676 6367 3683 6634
rect 3696 6367 3703 6953
rect 3716 6887 3723 7133
rect 3716 6603 3723 6852
rect 3736 6827 3743 7416
rect 3756 6907 3763 7423
rect 3796 7420 3803 7423
rect 3793 7407 3807 7420
rect 3856 7267 3863 7793
rect 3836 7156 3843 7193
rect 3876 7187 3883 8113
rect 3896 7407 3903 8213
rect 3916 8187 3923 8213
rect 4036 8196 4043 8373
rect 3936 8147 3943 8193
rect 3976 8160 3983 8163
rect 3956 8127 3963 8153
rect 3973 8147 3987 8160
rect 4076 8163 4083 8613
rect 4096 8227 4103 8593
rect 4136 8567 4143 8633
rect 4156 8507 4163 8673
rect 4176 8607 4183 9093
rect 4236 9087 4243 9192
rect 4213 9020 4227 9033
rect 4256 9028 4263 9373
rect 4216 9016 4223 9020
rect 4196 8587 4203 8793
rect 4216 8607 4223 8873
rect 4236 8867 4243 8983
rect 4276 8927 4283 9393
rect 4296 9327 4303 9513
rect 4296 9227 4303 9273
rect 4316 9183 4323 9633
rect 4436 9587 4443 9773
rect 4476 9727 4483 9754
rect 4376 9506 4383 9573
rect 4413 9540 4427 9553
rect 4453 9540 4467 9553
rect 4496 9548 4503 9913
rect 4596 9756 4603 9793
rect 4616 9787 4623 9853
rect 4536 9687 4543 9723
rect 4576 9667 4583 9723
rect 4416 9536 4423 9540
rect 4456 9536 4463 9540
rect 4476 9496 4503 9503
rect 4456 9267 4463 9473
rect 4387 9263 4400 9267
rect 4387 9253 4403 9263
rect 4336 9207 4343 9253
rect 4396 9236 4403 9253
rect 4316 9176 4343 9183
rect 4236 8686 4243 8733
rect 4236 8547 4243 8672
rect 4256 8547 4263 8713
rect 4276 8667 4283 8773
rect 4316 8748 4323 8993
rect 4336 8947 4343 9176
rect 4436 9167 4443 9223
rect 4356 8987 4363 9153
rect 4476 9107 4483 9453
rect 4496 9287 4503 9496
rect 4516 9467 4523 9553
rect 4536 9223 4543 9633
rect 4616 9487 4623 9553
rect 4636 9543 4643 9873
rect 4656 9707 4663 10453
rect 4676 10127 4683 10413
rect 4736 10276 4743 10536
rect 4796 10347 4803 10574
rect 4816 10487 4823 10814
rect 4696 10087 4703 10233
rect 4716 10127 4723 10243
rect 4776 10167 4783 10263
rect 4756 10083 4763 10133
rect 4776 10107 4783 10153
rect 4756 10080 4783 10083
rect 4756 10076 4787 10080
rect 4696 10036 4703 10073
rect 4773 10067 4787 10076
rect 4767 10036 4783 10043
rect 4696 9687 4703 9833
rect 4636 9536 4663 9543
rect 4696 9536 4703 9593
rect 4716 9567 4723 10034
rect 4776 10007 4783 10036
rect 4796 9967 4803 10033
rect 4816 10007 4823 10473
rect 4836 10467 4843 11133
rect 4856 10547 4863 11243
rect 4876 10527 4883 11094
rect 4976 10796 4983 11013
rect 4936 10576 4943 10613
rect 4956 10527 4963 10763
rect 5076 10543 5083 11133
rect 5096 10804 5103 11243
rect 5177 11063 5184 11243
rect 5176 11060 5184 11063
rect 5177 11057 5184 11060
rect 5356 11063 5363 11243
rect 5356 11056 5444 11063
rect 5096 10797 5164 10804
rect 5076 10536 5123 10543
rect 4856 10347 4863 10373
rect 4836 10260 4843 10263
rect 4833 10247 4847 10260
rect 4876 10207 4883 10513
rect 5116 10307 5123 10513
rect 5176 10296 5183 10473
rect 5196 10407 5203 10763
rect 5356 10627 5363 10853
rect 5458 10804 5465 11243
rect 5616 11096 5623 11133
rect 5656 11058 5663 11243
rect 5416 10797 5465 10804
rect 4836 9987 4843 10193
rect 4856 10027 4863 10053
rect 4736 9767 4743 9873
rect 4776 9787 4783 9833
rect 4773 9760 4787 9773
rect 4776 9756 4783 9760
rect 4756 9687 4763 9723
rect 4676 9447 4683 9503
rect 4696 9367 4703 9413
rect 4716 9407 4723 9503
rect 4753 9407 4767 9413
rect 4496 9220 4503 9223
rect 4493 9207 4507 9220
rect 4516 9216 4543 9223
rect 4436 9016 4443 9053
rect 4416 8967 4423 8983
rect 4456 8963 4463 8983
rect 4456 8956 4483 8963
rect 4396 8727 4403 8753
rect 4336 8623 4343 8683
rect 4376 8663 4383 8683
rect 4356 8660 4383 8663
rect 4353 8656 4383 8660
rect 4353 8647 4367 8656
rect 4366 8640 4367 8647
rect 4373 8623 4387 8633
rect 4336 8620 4387 8623
rect 4336 8616 4383 8620
rect 4396 8607 4403 8673
rect 4416 8627 4423 8953
rect 4436 8603 4443 8933
rect 4476 8927 4483 8956
rect 4416 8596 4443 8603
rect 4136 8467 4143 8493
rect 4096 8167 4103 8213
rect 4056 8156 4083 8163
rect 3933 8007 3947 8013
rect 3916 7946 3923 7993
rect 3996 7976 4003 8033
rect 4036 7988 4043 8053
rect 4056 8007 4063 8156
rect 4093 7967 4107 7974
rect 3896 7247 3903 7393
rect 3916 7323 3923 7932
rect 3976 7887 3983 7911
rect 4036 7907 4043 7933
rect 4013 7887 4027 7893
rect 3936 7666 3943 7733
rect 3976 7676 3983 7873
rect 4033 7847 4047 7853
rect 4056 7767 4063 7932
rect 4076 7807 4083 7953
rect 4016 7676 4023 7753
rect 4060 7683 4073 7687
rect 4056 7676 4073 7683
rect 4060 7673 4073 7676
rect 3996 7640 4003 7643
rect 3993 7627 4007 7640
rect 3956 7327 3963 7513
rect 3976 7507 3983 7573
rect 3996 7527 4003 7613
rect 4016 7547 4023 7593
rect 4036 7507 4043 7643
rect 4076 7507 4083 7553
rect 4096 7487 4103 7932
rect 4033 7460 4047 7472
rect 4036 7456 4043 7460
rect 3916 7316 3943 7323
rect 3916 7223 3923 7273
rect 3896 7216 3923 7223
rect 3896 7156 3903 7216
rect 3776 6863 3783 7112
rect 3796 6887 3803 7053
rect 3853 6940 3867 6953
rect 3856 6936 3863 6940
rect 3836 6867 3843 6903
rect 3876 6900 3883 6903
rect 3873 6887 3887 6900
rect 3916 6887 3923 7153
rect 3936 6867 3943 7316
rect 3976 7307 3983 7413
rect 4056 7420 4063 7423
rect 4053 7407 4067 7420
rect 3776 6856 3803 6863
rect 3756 6707 3763 6753
rect 3796 6636 3803 6856
rect 3916 6856 3933 6863
rect 3836 6636 3843 6793
rect 3716 6596 3733 6603
rect 3596 6256 3623 6263
rect 3533 6067 3547 6073
rect 3556 6047 3563 6114
rect 3596 6087 3603 6233
rect 3576 5896 3583 5973
rect 3616 5847 3623 6256
rect 3736 6247 3743 6592
rect 3776 6583 3783 6603
rect 3876 6603 3883 6852
rect 3856 6596 3883 6603
rect 3756 6576 3783 6583
rect 3673 6120 3687 6133
rect 3676 6116 3683 6120
rect 3716 6116 3723 6153
rect 3496 5376 3503 5453
rect 3536 5376 3543 5493
rect 3436 5256 3463 5263
rect 3433 5080 3447 5093
rect 3436 5076 3443 5080
rect 3396 4987 3403 5043
rect 3456 5007 3463 5256
rect 3536 5046 3543 5093
rect 3396 4827 3403 4952
rect 3476 4856 3483 4933
rect 3396 4727 3403 4773
rect 3336 4556 3343 4653
rect 3373 4560 3387 4573
rect 3376 4556 3383 4560
rect 3296 4516 3323 4523
rect 3236 4300 3243 4303
rect 3233 4287 3247 4300
rect 3193 4207 3207 4213
rect 3076 3947 3083 4052
rect 3096 3823 3103 4073
rect 3176 4036 3183 4133
rect 3236 4067 3243 4273
rect 3136 3987 3143 4033
rect 3136 3976 3153 3987
rect 3140 3973 3153 3976
rect 3196 3967 3203 4003
rect 3216 3947 3223 3973
rect 3156 3867 3163 3893
rect 3076 3816 3103 3823
rect 3116 3816 3123 3853
rect 3156 3816 3163 3853
rect 3053 3707 3067 3713
rect 3016 3627 3023 3673
rect 3076 3547 3083 3816
rect 2956 3456 2983 3463
rect 2836 3347 2843 3393
rect 2816 3227 2823 3273
rect 2816 2907 2823 3093
rect 2836 2863 2843 3333
rect 2896 3296 2903 3353
rect 2976 3287 2983 3456
rect 2960 3266 2980 3267
rect 2856 3256 2883 3263
rect 2856 3127 2863 3256
rect 2967 3253 2973 3266
rect 2896 3167 2903 3233
rect 2816 2856 2843 2863
rect 2693 2480 2707 2493
rect 2696 2476 2703 2480
rect 2756 2436 2783 2443
rect 2616 2256 2663 2263
rect 2693 2260 2707 2273
rect 2696 2256 2703 2260
rect 2616 2187 2623 2256
rect 2556 1887 2563 1973
rect 2633 1968 2647 1973
rect 2616 1827 2623 1923
rect 2656 1887 2663 1923
rect 2656 1687 2663 1713
rect 2656 1627 2663 1652
rect 2536 1347 2543 1403
rect 2676 1347 2683 1734
rect 2556 1167 2563 1214
rect 2596 943 2603 1033
rect 2616 967 2623 1183
rect 2596 936 2623 943
rect 2616 916 2623 936
rect 2476 696 2503 703
rect 2536 696 2543 773
rect 2676 767 2683 933
rect 2476 366 2483 696
rect 2516 660 2523 663
rect 2513 647 2527 660
rect 2636 427 2643 753
rect 2696 743 2703 2173
rect 2716 1787 2723 2223
rect 2736 1747 2743 2153
rect 2756 1567 2763 2413
rect 2776 2367 2783 2436
rect 2776 1807 2783 2353
rect 2796 2207 2803 2672
rect 2816 2427 2823 2856
rect 2856 2788 2863 3113
rect 2896 3067 2903 3113
rect 2996 3047 3003 3513
rect 3116 3486 3123 3533
rect 3136 3528 3143 3783
rect 3036 3480 3043 3483
rect 3016 3367 3023 3473
rect 3033 3467 3047 3480
rect 3156 3467 3163 3633
rect 3016 3107 3023 3294
rect 3036 3287 3043 3432
rect 3136 3387 3143 3433
rect 3107 3353 3113 3367
rect 3056 3267 3063 3333
rect 3176 3296 3183 3773
rect 3196 3427 3203 3753
rect 3156 3260 3163 3263
rect 3153 3247 3167 3260
rect 2896 2996 2903 3032
rect 2996 2967 3003 2994
rect 2956 2907 2963 2963
rect 2956 2896 2973 2907
rect 2960 2893 2973 2896
rect 2816 2187 2823 2254
rect 2836 2067 2843 2553
rect 2856 2167 2863 2693
rect 2876 2687 2883 2743
rect 2996 2607 3003 2913
rect 3036 2907 3043 3233
rect 3096 3207 3103 3233
rect 3076 3008 3083 3053
rect 3016 2747 3023 2853
rect 3056 2776 3063 2813
rect 3096 2787 3103 3153
rect 3116 3067 3123 3173
rect 3136 2996 3143 3113
rect 3216 3107 3223 3912
rect 3236 3807 3243 3893
rect 3256 3787 3263 4273
rect 3276 4147 3283 4303
rect 3276 3867 3283 4093
rect 3236 3567 3243 3753
rect 3256 3687 3263 3733
rect 3276 3647 3283 3814
rect 3296 3707 3303 4233
rect 3316 3987 3323 4516
rect 3356 4487 3363 4523
rect 3416 4467 3423 4854
rect 3556 4827 3563 5074
rect 3336 3828 3343 4453
rect 3436 4443 3443 4813
rect 3456 4787 3463 4823
rect 3496 4820 3503 4823
rect 3493 4807 3507 4820
rect 3476 4547 3483 4693
rect 3416 4436 3443 4443
rect 3356 3847 3363 4413
rect 3376 4047 3383 4334
rect 3416 4107 3423 4436
rect 3496 4427 3503 4793
rect 3516 4487 3523 4753
rect 3536 4583 3543 4653
rect 3556 4627 3563 4653
rect 3576 4607 3583 5493
rect 3636 5347 3643 6073
rect 3656 5987 3663 6083
rect 3696 6047 3703 6083
rect 3756 6067 3763 6576
rect 3836 6507 3843 6573
rect 3856 6567 3863 6596
rect 3776 6367 3783 6493
rect 3856 6416 3863 6493
rect 3896 6427 3903 6753
rect 3836 6363 3843 6383
rect 3836 6356 3863 6363
rect 3776 6187 3783 6293
rect 3656 5103 3663 5952
rect 3716 5747 3723 5973
rect 3776 5896 3783 6093
rect 3816 6086 3823 6353
rect 3816 5987 3823 6072
rect 3836 6007 3843 6273
rect 3796 5767 3803 5863
rect 3856 5847 3863 6356
rect 3916 6347 3923 6856
rect 3936 6587 3943 6813
rect 3936 6287 3943 6552
rect 3956 6428 3963 7173
rect 3976 7107 3983 7293
rect 3976 6447 3983 7053
rect 3996 6867 4003 7373
rect 4056 7167 4063 7393
rect 4096 7168 4103 7412
rect 4116 7383 4123 8452
rect 4136 7847 4143 8152
rect 4156 7927 4163 8413
rect 4176 8247 4183 8513
rect 4193 8447 4207 8453
rect 4196 8307 4203 8412
rect 4216 8267 4223 8463
rect 4236 8243 4243 8393
rect 4296 8287 4303 8593
rect 4216 8240 4243 8243
rect 4213 8236 4243 8240
rect 4213 8228 4227 8236
rect 4256 8196 4263 8273
rect 4176 8087 4183 8193
rect 4196 8067 4203 8153
rect 4236 8127 4243 8163
rect 4216 7976 4223 8093
rect 4256 7988 4263 8033
rect 4236 7940 4243 7943
rect 4233 7927 4247 7940
rect 4173 7887 4187 7893
rect 4167 7833 4173 7847
rect 4136 7823 4143 7833
rect 4136 7816 4163 7823
rect 4136 7707 4143 7733
rect 4136 7407 4143 7693
rect 4156 7507 4163 7816
rect 4116 7376 4143 7383
rect 4036 6943 4043 7093
rect 4076 6967 4083 7123
rect 4116 7007 4123 7073
rect 4036 6936 4063 6943
rect 4093 6940 4107 6953
rect 4096 6936 4103 6940
rect 4136 6903 4143 7376
rect 4156 7147 4163 7412
rect 4176 7387 4183 7793
rect 4173 7168 4187 7173
rect 4196 7163 4203 7911
rect 4296 7867 4303 7993
rect 4316 7747 4323 8313
rect 4336 7827 4343 8533
rect 4356 8387 4363 8593
rect 4416 8496 4423 8596
rect 4476 8527 4483 8913
rect 4496 8527 4503 8813
rect 4516 8547 4523 9216
rect 4696 9227 4703 9273
rect 4536 9147 4543 9193
rect 4556 8986 4563 9053
rect 4536 8727 4543 8893
rect 4576 8767 4583 9093
rect 4676 9047 4683 9073
rect 4616 8947 4623 9013
rect 4756 8983 4763 9113
rect 4716 8976 4763 8983
rect 4593 8720 4607 8733
rect 4596 8716 4603 8720
rect 4616 8667 4623 8683
rect 4616 8656 4633 8667
rect 4620 8653 4633 8656
rect 4656 8587 4663 8693
rect 4696 8627 4703 8714
rect 4716 8707 4723 8953
rect 4736 8907 4743 8976
rect 4776 8963 4783 9693
rect 4796 9506 4803 9593
rect 4796 9287 4803 9353
rect 4816 9267 4823 9393
rect 4836 9327 4843 9453
rect 4856 9283 4863 9992
rect 4876 9467 4883 10113
rect 4936 10020 4943 10023
rect 4933 10007 4947 10020
rect 5036 9987 5043 10053
rect 5076 10027 5083 10054
rect 5096 10047 5103 10153
rect 5116 10023 5123 10293
rect 5156 10068 5163 10233
rect 5216 10167 5223 10473
rect 5233 10247 5247 10253
rect 5240 10226 5260 10227
rect 5247 10213 5253 10226
rect 5116 10016 5143 10023
rect 4896 9647 4903 9973
rect 5016 9756 5023 9873
rect 4916 9536 4923 9754
rect 5036 9667 5043 9723
rect 4953 9540 4967 9553
rect 4956 9536 4963 9540
rect 4976 9500 4983 9503
rect 4973 9487 4987 9500
rect 4887 9393 4893 9407
rect 4847 9276 4863 9283
rect 4833 9260 4847 9273
rect 4836 9256 4843 9260
rect 4796 9220 4803 9223
rect 4793 9207 4807 9220
rect 4796 8967 4803 9093
rect 4756 8956 4783 8963
rect 4736 8687 4743 8872
rect 4356 7907 4363 8373
rect 4436 8367 4443 8463
rect 4456 8387 4463 8433
rect 4356 7727 4363 7773
rect 4376 7767 4383 8333
rect 4396 8007 4403 8273
rect 4496 8166 4503 8193
rect 4416 8156 4443 8163
rect 4233 7680 4247 7693
rect 4273 7680 4287 7693
rect 4236 7676 4243 7680
rect 4276 7676 4283 7680
rect 4256 7640 4263 7643
rect 4253 7627 4267 7640
rect 4316 7643 4323 7693
rect 4307 7636 4323 7643
rect 4216 7456 4243 7463
rect 4216 7367 4223 7456
rect 4296 7423 4303 7632
rect 4356 7627 4363 7692
rect 4376 7427 4383 7732
rect 4396 7527 4403 7972
rect 4416 7567 4423 8156
rect 4496 8107 4503 8152
rect 4436 7907 4443 7943
rect 4496 7807 4503 7943
rect 4516 7927 4523 8512
rect 4536 8466 4543 8493
rect 4513 7887 4527 7892
rect 4436 7687 4443 7733
rect 4453 7680 4467 7693
rect 4456 7676 4463 7680
rect 4536 7687 4543 8452
rect 4556 8427 4563 8513
rect 4676 8496 4683 8593
rect 4716 8496 4723 8672
rect 4756 8467 4763 8956
rect 4776 8727 4783 8873
rect 4816 8807 4823 8993
rect 4836 8887 4843 9053
rect 4856 9047 4863 9153
rect 4876 9023 4883 9333
rect 4916 9207 4923 9353
rect 4956 9347 4963 9453
rect 4936 9107 4943 9293
rect 4956 9127 4963 9293
rect 4856 9016 4883 9023
rect 4856 8927 4863 9016
rect 4976 9027 4983 9413
rect 4996 9087 5003 9493
rect 5016 9307 5023 9553
rect 5036 9527 5043 9653
rect 5056 9503 5063 9633
rect 5096 9603 5103 9853
rect 5036 9496 5063 9503
rect 5076 9596 5103 9603
rect 5036 9307 5043 9496
rect 5056 9367 5063 9473
rect 5056 9236 5063 9313
rect 5076 9307 5083 9596
rect 5116 9587 5123 9754
rect 5136 9727 5143 10016
rect 5176 9907 5183 10023
rect 5216 9987 5223 10023
rect 5236 9927 5243 10013
rect 5256 9947 5263 10053
rect 5276 9907 5283 10574
rect 5376 10547 5383 10763
rect 5096 9367 5103 9573
rect 5176 9536 5183 9712
rect 5216 9536 5223 9613
rect 5113 9527 5127 9534
rect 5296 9503 5303 10353
rect 5316 10267 5323 10393
rect 5396 10367 5403 10613
rect 5496 10583 5503 10873
rect 5496 10576 5523 10583
rect 5556 10576 5563 10853
rect 5699 10804 5706 11243
rect 5636 10797 5706 10804
rect 5596 10576 5603 10613
rect 5536 10523 5543 10543
rect 5516 10516 5543 10523
rect 5516 10367 5523 10516
rect 5393 10280 5407 10293
rect 5396 10276 5403 10280
rect 5367 10246 5380 10247
rect 5367 10233 5373 10246
rect 5416 10223 5423 10243
rect 5476 10227 5483 10274
rect 5496 10247 5503 10313
rect 5367 10216 5423 10223
rect 5316 9867 5323 10113
rect 5316 9647 5323 9793
rect 5156 9447 5163 9503
rect 5196 9483 5203 9503
rect 5276 9496 5303 9503
rect 5196 9476 5223 9483
rect 5093 9240 5107 9253
rect 5096 9236 5103 9240
rect 5036 9167 5043 9203
rect 5116 9187 5123 9203
rect 5096 9176 5113 9183
rect 5040 9143 5053 9147
rect 5036 9133 5053 9143
rect 4956 9016 4973 9023
rect 4996 8986 5003 9052
rect 4896 8947 4903 8983
rect 4920 8965 4940 8967
rect 4927 8953 4933 8965
rect 4876 8787 4883 8853
rect 4956 8827 4963 8933
rect 4907 8793 4913 8807
rect 4776 8487 4783 8673
rect 4820 8665 4833 8667
rect 4827 8653 4833 8665
rect 4876 8627 4883 8673
rect 4896 8647 4903 8714
rect 4916 8687 4923 8772
rect 4936 8747 4943 8773
rect 4556 7947 4563 8033
rect 4576 7867 4583 8233
rect 4636 8196 4643 8453
rect 4656 8407 4663 8463
rect 4696 8247 4703 8463
rect 4736 8347 4743 8453
rect 4596 8156 4623 8163
rect 4476 7607 4483 7643
rect 4416 7467 4423 7553
rect 4456 7547 4463 7573
rect 4476 7456 4483 7493
rect 4516 7456 4523 7573
rect 4276 7416 4303 7423
rect 4296 7207 4303 7416
rect 4196 7156 4223 7163
rect 4293 7160 4307 7172
rect 4333 7160 4347 7173
rect 4356 7167 4363 7353
rect 4496 7327 4503 7423
rect 4556 7327 4563 7813
rect 4596 7683 4603 8156
rect 4616 7827 4623 8053
rect 4776 8047 4783 8473
rect 4796 8387 4803 8573
rect 4816 8327 4823 8613
rect 4936 8587 4943 8693
rect 4956 8687 4963 8733
rect 4976 8667 4983 8793
rect 4916 8496 4923 8533
rect 4956 8496 4963 8553
rect 4973 8507 4987 8513
rect 4853 8467 4867 8473
rect 4876 8327 4883 8353
rect 4896 8347 4903 8463
rect 4836 8196 4843 8233
rect 4816 8007 4823 8163
rect 4916 8127 4923 8413
rect 4936 8407 4943 8463
rect 4996 8447 5003 8913
rect 5016 8887 5023 9013
rect 5036 8867 5043 9133
rect 5076 9067 5083 9153
rect 5076 8986 5083 9013
rect 5096 8927 5103 9176
rect 5156 9147 5163 9293
rect 5176 9187 5183 9233
rect 5116 9028 5123 9053
rect 5136 9016 5143 9113
rect 5196 9107 5203 9433
rect 5216 9387 5223 9476
rect 5276 9427 5283 9496
rect 5336 9487 5343 10193
rect 5436 10056 5443 10153
rect 5476 10056 5483 10113
rect 5356 10027 5363 10054
rect 5416 10020 5423 10023
rect 5356 9867 5363 10013
rect 5413 10007 5427 10020
rect 5456 10003 5463 10023
rect 5516 10007 5523 10353
rect 5536 10067 5543 10413
rect 5576 10363 5583 10532
rect 5656 10427 5663 10573
rect 5676 10487 5683 10574
rect 5556 10356 5583 10363
rect 5436 9996 5463 10003
rect 5436 9967 5443 9996
rect 5216 9187 5223 9333
rect 5236 9207 5243 9234
rect 5256 9187 5263 9273
rect 5276 9247 5283 9293
rect 5296 9236 5303 9473
rect 5356 9447 5363 9793
rect 5396 9536 5403 9893
rect 5436 9807 5443 9953
rect 5456 9687 5463 9723
rect 5116 8827 5123 8953
rect 5016 8727 5023 8793
rect 5033 8720 5047 8733
rect 5073 8720 5087 8733
rect 5036 8716 5043 8720
rect 5076 8716 5083 8720
rect 5100 8684 5113 8687
rect 5096 8677 5113 8684
rect 5100 8673 5113 8677
rect 5056 8647 5063 8672
rect 5016 8527 5023 8553
rect 5036 8487 5043 8533
rect 4936 8087 4943 8194
rect 4680 8003 4693 8007
rect 4676 7993 4693 8003
rect 4676 7976 4683 7993
rect 4647 7893 4653 7907
rect 4696 7887 4703 7943
rect 4736 7907 4743 7943
rect 4796 7927 4803 7993
rect 4816 7887 4823 7933
rect 4587 7676 4603 7683
rect 4576 7607 4583 7674
rect 4616 7247 4623 7673
rect 4636 7527 4643 7872
rect 4656 7587 4663 7773
rect 4716 7676 4723 7833
rect 4796 7707 4803 7733
rect 4696 7607 4703 7643
rect 4796 7627 4803 7693
rect 4816 7646 4823 7833
rect 4636 7347 4643 7453
rect 4656 7387 4663 7493
rect 4716 7456 4723 7513
rect 4756 7456 4763 7553
rect 4676 7287 4683 7413
rect 4696 7367 4703 7423
rect 4456 7187 4463 7233
rect 4296 7156 4303 7160
rect 4336 7156 4343 7160
rect 4036 6636 4043 6893
rect 4076 6867 4083 6903
rect 4116 6896 4143 6903
rect 4056 6647 4063 6733
rect 4116 6623 4123 6896
rect 4136 6767 4143 6873
rect 4156 6847 4163 7013
rect 4176 6967 4183 7154
rect 4096 6616 4123 6623
rect 4016 6547 4023 6603
rect 4076 6487 4083 6612
rect 4076 6447 4083 6473
rect 4096 6428 4103 6616
rect 4136 6587 4143 6623
rect 4136 6527 4143 6573
rect 4136 6467 4143 6513
rect 3907 6143 3920 6147
rect 3907 6133 3923 6143
rect 3916 6116 3923 6133
rect 3936 6067 3943 6083
rect 3713 5600 3727 5613
rect 3716 5596 3723 5600
rect 3676 5427 3683 5563
rect 3736 5247 3743 5343
rect 3656 5096 3683 5103
rect 3676 5076 3683 5096
rect 3616 4627 3623 5032
rect 3536 4576 3563 4583
rect 3556 4556 3563 4576
rect 3613 4507 3627 4513
rect 3636 4487 3643 4993
rect 3656 4787 3663 5043
rect 3756 4927 3763 5313
rect 3776 5187 3783 5273
rect 3753 4848 3767 4854
rect 3656 4607 3663 4693
rect 3393 4040 3407 4053
rect 3396 4036 3403 4040
rect 3436 4036 3443 4133
rect 3456 4087 3463 4273
rect 3476 4227 3483 4303
rect 3516 4300 3523 4303
rect 3513 4287 3527 4300
rect 3456 4043 3463 4073
rect 3476 4067 3483 4133
rect 3456 4036 3483 4043
rect 3376 3887 3383 3993
rect 3396 3867 3403 3973
rect 3413 3820 3427 3833
rect 3436 3827 3443 3933
rect 3456 3907 3463 3993
rect 3416 3816 3423 3820
rect 3456 3786 3463 3853
rect 3313 3763 3327 3773
rect 3313 3760 3343 3763
rect 3316 3756 3343 3760
rect 3336 3587 3343 3756
rect 3356 3716 3403 3723
rect 3356 3687 3363 3716
rect 3276 3516 3283 3573
rect 3256 3467 3263 3483
rect 3296 3480 3303 3483
rect 3293 3467 3307 3480
rect 3267 3456 3283 3463
rect 3236 3266 3243 3353
rect 3216 3007 3223 3093
rect 3116 2747 3123 2893
rect 2896 2467 2903 2513
rect 2996 2446 3003 2593
rect 2936 2256 2943 2413
rect 2956 2267 2963 2353
rect 2936 2167 2943 2193
rect 2796 1903 2803 2033
rect 2876 1956 2883 2053
rect 2956 2047 2963 2173
rect 2796 1896 2813 1903
rect 2816 1736 2823 1893
rect 2896 1787 2903 1923
rect 2796 1436 2803 1671
rect 2836 1647 2843 1703
rect 2876 1700 2883 1703
rect 2873 1687 2887 1700
rect 2716 1287 2723 1353
rect 2736 1267 2743 1403
rect 2836 1367 2843 1553
rect 2896 1407 2903 1493
rect 2716 886 2723 1213
rect 2736 927 2743 1253
rect 2836 1216 2843 1293
rect 2816 948 2823 1183
rect 2876 1007 2883 1183
rect 2916 1167 2923 1734
rect 2936 1687 2943 1773
rect 2956 1443 2963 1913
rect 2976 1607 2983 2433
rect 2996 2147 3003 2373
rect 3016 1847 3023 2553
rect 3036 2207 3043 2593
rect 3056 2227 3063 2474
rect 3036 2007 3043 2053
rect 3056 1956 3063 2133
rect 3076 2007 3083 2653
rect 3096 2447 3103 2693
rect 3136 2476 3143 2773
rect 3156 2627 3163 2893
rect 3196 2667 3203 2893
rect 3216 2767 3223 2953
rect 3156 2440 3163 2443
rect 3153 2427 3167 2440
rect 3196 2407 3203 2443
rect 3236 2387 3243 3252
rect 3256 2907 3263 3413
rect 3276 2967 3283 3456
rect 3296 3087 3303 3213
rect 3116 2256 3123 2313
rect 3256 2268 3263 2743
rect 3316 2687 3323 3313
rect 3336 3247 3343 3473
rect 3356 3327 3363 3633
rect 3376 3487 3383 3693
rect 3396 3687 3403 3716
rect 3456 3707 3463 3733
rect 3396 3467 3403 3633
rect 3476 3607 3483 4036
rect 3496 3747 3503 3813
rect 3516 3767 3523 4073
rect 3536 3927 3543 4293
rect 3556 4287 3563 4393
rect 3556 4007 3563 4093
rect 3596 4067 3603 4473
rect 3656 4463 3663 4554
rect 3676 4526 3683 4673
rect 3636 4456 3663 4463
rect 3636 4307 3643 4456
rect 3676 4347 3683 4393
rect 3696 4367 3703 4713
rect 3736 4707 3743 4813
rect 3796 4767 3803 5293
rect 3816 5087 3823 5373
rect 3836 5227 3843 5693
rect 3896 5608 3903 6051
rect 3916 5667 3923 5993
rect 3936 5827 3943 6053
rect 3976 6047 3983 6412
rect 3996 6386 4003 6413
rect 4016 5987 4023 6053
rect 4036 6007 4043 6313
rect 4076 6283 4083 6383
rect 4056 6276 4083 6283
rect 4056 6067 4063 6276
rect 4076 6067 4083 6233
rect 4136 6187 4143 6293
rect 4136 6116 4143 6173
rect 4053 5888 4067 5894
rect 4096 5883 4103 6113
rect 4116 5967 4123 6013
rect 4136 5887 4143 6033
rect 4096 5876 4123 5883
rect 3996 5860 4003 5863
rect 3936 5547 3943 5713
rect 3956 5707 3963 5853
rect 3993 5847 4007 5860
rect 3976 5687 3983 5833
rect 3976 5388 3983 5673
rect 3996 5487 4003 5812
rect 3856 5346 3863 5373
rect 3956 5207 3963 5343
rect 4016 5307 4023 5613
rect 4036 5567 4043 5853
rect 4096 5596 4103 5813
rect 4136 5627 4143 5833
rect 4120 5563 4133 5567
rect 4076 5560 4083 5563
rect 4073 5547 4087 5560
rect 4116 5556 4133 5563
rect 4120 5553 4133 5556
rect 4156 5547 4163 6414
rect 4176 6047 4183 6953
rect 4196 6827 4203 6953
rect 4216 6867 4223 7156
rect 4416 7146 4423 7173
rect 4276 7107 4283 7123
rect 4236 6807 4243 7013
rect 4276 6967 4283 7093
rect 4376 7027 4383 7132
rect 4376 6967 4383 7013
rect 4393 6967 4407 6973
rect 4333 6947 4347 6953
rect 4253 6847 4267 6853
rect 4276 6747 4283 6903
rect 4296 6727 4303 6793
rect 4356 6767 4363 6953
rect 4416 6906 4423 6933
rect 4316 6616 4323 6753
rect 4436 6723 4443 7143
rect 4476 6943 4483 7213
rect 4716 7027 4723 7353
rect 4796 7227 4803 7493
rect 4796 7183 4803 7213
rect 4776 7176 4803 7183
rect 4796 7027 4803 7073
rect 4816 7067 4823 7632
rect 4836 7627 4843 8073
rect 4956 8067 4963 8433
rect 4976 8127 4983 8233
rect 4996 8163 5003 8333
rect 5016 8307 5023 8353
rect 5056 8287 5063 8493
rect 5076 8447 5083 8613
rect 5116 8607 5123 8652
rect 5136 8547 5143 8913
rect 5156 8527 5163 8733
rect 5196 8687 5203 8951
rect 5176 8496 5183 8653
rect 5216 8627 5223 8873
rect 5236 8547 5243 9014
rect 5256 8967 5263 9073
rect 5276 9007 5283 9133
rect 5116 8367 5123 8463
rect 5096 8307 5103 8353
rect 5093 8200 5107 8213
rect 5136 8203 5143 8433
rect 5156 8427 5163 8463
rect 5156 8227 5163 8333
rect 5193 8207 5207 8213
rect 5096 8196 5103 8200
rect 5136 8196 5163 8203
rect 5156 8167 5163 8196
rect 4996 8156 5023 8163
rect 4976 7976 4983 8013
rect 4993 7987 5007 7993
rect 5016 7947 5023 8156
rect 5036 8027 5043 8163
rect 5116 8143 5123 8163
rect 5096 8136 5123 8143
rect 5056 8087 5063 8133
rect 4916 7940 4923 7943
rect 4856 7583 4863 7913
rect 4876 7647 4883 7753
rect 4847 7576 4863 7583
rect 4836 7426 4843 7573
rect 4836 7227 4843 7273
rect 4856 7267 4863 7513
rect 4876 7367 4883 7612
rect 4856 7183 4863 7232
rect 4836 7176 4863 7183
rect 4836 7067 4843 7176
rect 4416 6716 4443 6723
rect 4456 6936 4483 6943
rect 4516 6936 4523 6973
rect 4416 6587 4423 6716
rect 4456 6707 4463 6936
rect 4596 6906 4603 6953
rect 4456 6663 4463 6693
rect 4456 6656 4483 6663
rect 4516 6627 4523 6753
rect 4236 6467 4243 6493
rect 4196 6107 4203 6353
rect 4216 6087 4223 6433
rect 4256 6128 4263 6513
rect 4293 6420 4307 6433
rect 4333 6420 4347 6433
rect 4296 6416 4303 6420
rect 4336 6416 4343 6420
rect 4396 6386 4403 6513
rect 4316 6047 4323 6383
rect 4356 6287 4363 6383
rect 4436 6327 4443 6553
rect 4536 6447 4543 6653
rect 4496 6436 4513 6443
rect 4496 6407 4503 6436
rect 4527 6436 4543 6447
rect 4527 6433 4540 6436
rect 4556 6416 4563 6813
rect 4576 6447 4583 6713
rect 4656 6707 4663 7013
rect 4733 6967 4747 6973
rect 4816 6967 4823 7053
rect 4696 6906 4703 6953
rect 4696 6648 4703 6853
rect 4836 6827 4843 6993
rect 4856 6947 4863 7154
rect 4876 6847 4883 7233
rect 4536 6327 4543 6383
rect 4576 6327 4583 6351
rect 4296 5827 4303 5883
rect 4196 5647 4203 5713
rect 4176 5567 4183 5593
rect 4036 5407 4043 5513
rect 3856 5076 3863 5153
rect 4076 5076 4083 5293
rect 4096 5147 4103 5374
rect 3836 4967 3843 5043
rect 4056 4987 4063 5043
rect 4116 5007 4123 5533
rect 4196 5376 4203 5612
rect 4236 5427 4243 5733
rect 4296 5608 4303 5753
rect 4216 5340 4223 5343
rect 4213 5327 4227 5340
rect 4256 5307 4263 5594
rect 4316 5560 4323 5563
rect 4313 5547 4327 5560
rect 4326 5540 4327 5547
rect 4156 4987 4163 5193
rect 3816 4836 3823 4873
rect 3736 4527 3743 4653
rect 3756 4556 3763 4673
rect 3813 4560 3827 4573
rect 3816 4556 3823 4560
rect 3767 4393 3773 4407
rect 3733 4340 3747 4353
rect 3736 4336 3743 4340
rect 3576 4056 3593 4063
rect 3576 4027 3583 4056
rect 3636 4036 3643 4253
rect 3673 4040 3687 4053
rect 3693 4047 3707 4053
rect 3676 4036 3683 4040
rect 3616 3987 3623 4003
rect 3616 3976 3633 3987
rect 3620 3973 3633 3976
rect 3536 3687 3543 3833
rect 3616 3816 3623 3933
rect 3556 3786 3563 3813
rect 3676 3683 3683 3772
rect 3696 3707 3703 3813
rect 3676 3676 3703 3683
rect 3436 3467 3443 3573
rect 3476 3527 3483 3572
rect 3496 3516 3503 3553
rect 3536 3548 3543 3673
rect 3676 3607 3683 3653
rect 3476 3427 3483 3473
rect 3596 3467 3603 3513
rect 3616 3487 3623 3573
rect 3696 3567 3703 3676
rect 3716 3667 3723 4173
rect 3736 4147 3743 4273
rect 3736 4007 3743 4133
rect 3756 3927 3763 4333
rect 3776 4227 3783 4313
rect 3736 3787 3743 3814
rect 3376 3256 3403 3263
rect 3376 2996 3383 3233
rect 3396 3027 3403 3256
rect 3436 3003 3443 3413
rect 3456 3227 3463 3273
rect 3476 3187 3483 3294
rect 3516 3223 3523 3333
rect 3536 3267 3543 3453
rect 3636 3347 3643 3453
rect 3656 3328 3663 3553
rect 3676 3487 3683 3533
rect 3696 3516 3703 3553
rect 3736 3407 3743 3483
rect 3516 3216 3543 3223
rect 3476 3127 3483 3173
rect 3436 2996 3463 3003
rect 3276 2447 3283 2613
rect 3336 2607 3343 2773
rect 3356 2583 3363 2963
rect 3396 2960 3403 2963
rect 3393 2947 3407 2960
rect 3336 2576 3363 2583
rect 3336 2407 3343 2576
rect 3416 2527 3423 2833
rect 3436 2567 3443 2973
rect 3456 2703 3463 2996
rect 3496 2947 3503 3113
rect 3476 2740 3483 2743
rect 3473 2727 3487 2740
rect 3456 2696 3483 2703
rect 3096 2167 3103 2213
rect 3127 2053 3133 2067
rect 3076 1887 3083 1923
rect 3116 1827 3123 1923
rect 3076 1736 3083 1793
rect 2936 1436 2963 1443
rect 2996 1436 3003 1473
rect 3036 1448 3043 1673
rect 3056 1627 3063 1703
rect 3073 1667 3087 1673
rect 3096 1587 3103 1673
rect 2856 916 2863 993
rect 2676 736 2703 743
rect 2676 666 2683 736
rect 2736 727 2743 913
rect 2696 666 2703 713
rect 2756 696 2763 773
rect 2796 696 2803 873
rect 2676 547 2683 593
rect 2636 396 2643 413
rect 2676 396 2683 533
rect 2436 360 2443 363
rect 2433 347 2447 360
rect 2616 287 2623 363
rect 2396 176 2403 213
rect 2656 176 2663 293
rect 2556 147 2563 174
rect 2736 168 2743 533
rect 2776 507 2783 663
rect 2816 447 2823 653
rect 2596 140 2603 143
rect 2593 127 2607 140
rect 2713 127 2727 132
rect 2756 127 2763 413
rect 2796 307 2803 413
rect 2836 383 2843 713
rect 2936 708 2943 1436
rect 2976 1228 2983 1403
rect 2976 1127 2983 1214
rect 2996 1067 3003 1273
rect 3016 1207 3023 1313
rect 3136 1287 3143 1913
rect 3156 1687 3163 1993
rect 3176 1748 3183 2093
rect 3216 2047 3223 2113
rect 3196 1687 3203 1873
rect 3036 1067 3043 1172
rect 3036 916 3043 1013
rect 3073 920 3087 933
rect 3116 927 3123 1172
rect 3076 916 3083 920
rect 3056 863 3063 883
rect 3056 856 3083 863
rect 2973 700 2987 713
rect 2976 696 2983 700
rect 3036 627 3043 663
rect 3076 627 3083 856
rect 3096 727 3103 883
rect 3116 666 3123 773
rect 2856 396 2863 453
rect 2816 376 2843 383
rect 2816 227 2823 376
rect 2836 188 2843 352
rect 2856 307 2863 333
rect 2876 176 2883 213
rect 3056 176 3063 473
rect 3096 396 3103 473
rect 3156 403 3163 1573
rect 3216 1467 3223 2033
rect 3236 1927 3243 2053
rect 3256 2007 3263 2254
rect 3276 2187 3283 2293
rect 3296 2227 3303 2313
rect 3396 2307 3403 2443
rect 3413 2263 3427 2273
rect 3396 2260 3427 2263
rect 3396 2256 3423 2260
rect 3376 2187 3383 2223
rect 3276 2067 3283 2113
rect 3353 1960 3367 1973
rect 3356 1956 3363 1960
rect 3256 1927 3263 1954
rect 3296 1807 3303 1923
rect 3296 1767 3303 1793
rect 3293 1740 3307 1753
rect 3296 1736 3303 1740
rect 3376 1707 3383 1913
rect 3396 1787 3403 1973
rect 3416 1887 3423 2093
rect 3436 1927 3443 2433
rect 3456 1967 3463 2673
rect 3476 2567 3483 2696
rect 3476 2407 3483 2553
rect 3476 2227 3483 2253
rect 3496 2127 3503 2673
rect 3516 2287 3523 2453
rect 3536 2263 3543 3216
rect 3556 3147 3563 3294
rect 3573 3187 3587 3193
rect 3596 3147 3603 3252
rect 3616 3127 3623 3233
rect 3636 3023 3643 3263
rect 3676 3027 3683 3231
rect 3716 3207 3723 3293
rect 3736 3247 3743 3313
rect 3716 3087 3723 3193
rect 3636 3016 3663 3023
rect 3556 2767 3563 3013
rect 3656 2967 3663 3016
rect 3616 2727 3623 2873
rect 3616 2488 3623 2653
rect 3656 2587 3663 2932
rect 3676 2927 3683 2992
rect 3696 2827 3703 3013
rect 3716 2803 3723 3013
rect 3696 2796 3723 2803
rect 3696 2776 3703 2796
rect 3736 2776 3743 2893
rect 3756 2847 3763 3913
rect 3776 3467 3783 4033
rect 3796 3907 3803 4473
rect 3816 4247 3823 4353
rect 3836 4263 3843 4733
rect 3856 4467 3863 4873
rect 3996 4807 4003 4843
rect 4016 4787 4023 4833
rect 3893 4407 3907 4413
rect 3916 4407 3923 4693
rect 3936 4487 3943 4673
rect 3956 4526 3963 4613
rect 3996 4583 4003 4653
rect 4036 4587 4043 4693
rect 3996 4576 4023 4583
rect 4016 4556 4023 4576
rect 3856 4287 3863 4353
rect 3887 4334 3893 4347
rect 3913 4340 3927 4353
rect 3916 4336 3923 4340
rect 3887 4333 3900 4334
rect 3936 4300 3943 4303
rect 3933 4287 3947 4300
rect 3836 4256 3863 4263
rect 3836 4067 3843 4193
rect 3856 4187 3863 4256
rect 3816 3996 3843 4003
rect 3816 3987 3823 3996
rect 3816 3827 3823 3973
rect 3853 3967 3867 3973
rect 3853 3960 3873 3967
rect 3856 3956 3873 3960
rect 3860 3953 3873 3956
rect 3893 3867 3907 3873
rect 3807 3816 3823 3827
rect 3853 3820 3867 3833
rect 3856 3816 3863 3820
rect 3807 3813 3820 3816
rect 3836 3763 3843 3772
rect 3816 3756 3843 3763
rect 3776 2947 3783 3432
rect 3796 3187 3803 3533
rect 3816 3447 3823 3756
rect 3836 3243 3843 3693
rect 3876 3567 3883 3783
rect 3916 3707 3923 3992
rect 3956 3967 3963 4213
rect 3876 3467 3883 3553
rect 3936 3547 3943 3893
rect 3956 3547 3963 3873
rect 3976 3767 3983 4253
rect 3996 4227 4003 4334
rect 3996 4027 4003 4073
rect 3913 3520 3927 3533
rect 3916 3516 3923 3520
rect 3956 3516 3963 3533
rect 3936 3467 3943 3483
rect 3927 3456 3943 3467
rect 3927 3453 3940 3456
rect 3876 3296 3883 3393
rect 3916 3260 3923 3263
rect 3913 3247 3927 3260
rect 3836 3236 3863 3243
rect 3833 3207 3847 3213
rect 3796 3003 3803 3173
rect 3836 3023 3843 3093
rect 3856 3067 3863 3236
rect 3876 3147 3883 3173
rect 3836 3016 3863 3023
rect 3796 2996 3823 3003
rect 3856 2996 3863 3016
rect 3596 2347 3603 2443
rect 3516 2256 3543 2263
rect 3556 2256 3563 2333
rect 3593 2268 3607 2273
rect 3516 2127 3523 2256
rect 3476 1767 3483 1993
rect 3496 1867 3503 1973
rect 3536 1956 3543 2173
rect 3576 2007 3583 2223
rect 3573 1960 3587 1972
rect 3616 1967 3623 2213
rect 3576 1956 3583 1960
rect 3556 1827 3563 1873
rect 3596 1847 3603 1923
rect 3467 1753 3483 1767
rect 3476 1736 3483 1753
rect 3516 1796 3583 1803
rect 3516 1736 3523 1796
rect 3556 1747 3563 1773
rect 3276 1467 3283 1692
rect 3416 1567 3423 1733
rect 3576 1706 3583 1796
rect 3496 1700 3503 1703
rect 3493 1687 3507 1700
rect 3176 1436 3223 1443
rect 3253 1440 3267 1453
rect 3256 1436 3263 1440
rect 3176 1407 3183 1436
rect 3396 1427 3403 1453
rect 3176 687 3183 1333
rect 3196 1186 3203 1293
rect 3236 1067 3243 1403
rect 3356 1216 3363 1373
rect 3256 1186 3263 1213
rect 3336 1087 3343 1183
rect 3236 947 3243 1053
rect 3313 920 3327 933
rect 3316 916 3323 920
rect 3376 887 3383 953
rect 3396 928 3403 1213
rect 3416 947 3423 1473
rect 3476 1436 3483 1553
rect 3536 1443 3543 1653
rect 3556 1467 3563 1513
rect 3516 1436 3543 1443
rect 3456 1127 3463 1392
rect 3496 1243 3503 1403
rect 3576 1307 3583 1553
rect 3596 1407 3603 1433
rect 3476 1236 3503 1243
rect 3476 1186 3483 1236
rect 3596 1228 3603 1372
rect 3636 1347 3643 2393
rect 3656 2187 3663 2254
rect 3656 1667 3663 2173
rect 3676 2107 3683 2633
rect 3696 2307 3703 2713
rect 3696 2167 3703 2212
rect 3676 1787 3683 1953
rect 3696 1947 3703 2113
rect 3716 2087 3723 2743
rect 3756 2707 3763 2743
rect 3796 2607 3803 2733
rect 3816 2707 3823 2933
rect 3836 2727 3843 2963
rect 3856 2627 3863 2773
rect 3876 2767 3883 2893
rect 3756 2387 3763 2573
rect 3876 2487 3883 2513
rect 3836 2387 3843 2443
rect 3776 2256 3783 2333
rect 3736 2147 3743 2233
rect 3776 1956 3783 2053
rect 3876 1968 3883 2473
rect 3896 2407 3903 3153
rect 3916 2947 3923 3212
rect 3936 3127 3943 3433
rect 3956 3247 3963 3393
rect 3976 3327 3983 3393
rect 3996 3167 4003 3992
rect 4016 3947 4023 4473
rect 4036 4147 4043 4523
rect 4096 4087 4103 4913
rect 4116 4836 4123 4972
rect 4196 4847 4203 5074
rect 4216 4887 4223 5292
rect 4316 5207 4323 5413
rect 4256 5076 4263 5153
rect 4336 5047 4343 5533
rect 4356 5387 4363 5563
rect 4396 5547 4403 6253
rect 4636 6207 4643 6414
rect 4676 6386 4683 6592
rect 4696 6447 4703 6513
rect 4716 6367 4723 6413
rect 4556 6086 4563 6113
rect 4456 5727 4463 5843
rect 4516 5607 4523 5874
rect 4576 5867 4583 5973
rect 4576 5687 4583 5832
rect 4596 5647 4603 6173
rect 4656 6116 4663 6333
rect 4700 6143 4713 6147
rect 4696 6133 4713 6143
rect 4696 6116 4703 6133
rect 4676 6047 4683 6083
rect 4376 5376 4383 5413
rect 4416 5376 4423 5473
rect 4436 5407 4443 5513
rect 4396 5247 4403 5343
rect 4436 5307 4443 5343
rect 4476 5247 4483 5593
rect 4576 5560 4583 5563
rect 4536 5367 4543 5552
rect 4573 5547 4587 5560
rect 4536 5347 4543 5353
rect 4556 5347 4563 5413
rect 4520 5346 4543 5347
rect 4527 5333 4543 5346
rect 4376 5167 4383 5213
rect 4396 5127 4403 5233
rect 4536 5043 4543 5333
rect 4556 5047 4563 5073
rect 4516 5036 4543 5043
rect 4256 4836 4283 4843
rect 4116 4347 4123 4773
rect 4156 4727 4163 4803
rect 4216 4727 4223 4803
rect 4276 4687 4283 4836
rect 4276 4676 4293 4687
rect 4280 4673 4293 4676
rect 4276 4556 4283 4593
rect 4136 4527 4143 4554
rect 4196 4487 4203 4533
rect 4036 3907 4043 3953
rect 4013 3867 4027 3873
rect 4053 3820 4067 3833
rect 4093 3820 4107 3833
rect 4116 3827 4123 4133
rect 4136 4107 4143 4303
rect 4236 4107 4243 4393
rect 4336 4207 4343 4433
rect 4436 4407 4443 4593
rect 4496 4556 4503 4593
rect 4456 4383 4463 4523
rect 4456 4376 4483 4383
rect 4396 4287 4403 4303
rect 4396 4276 4413 4287
rect 4400 4273 4413 4276
rect 4436 4247 4443 4293
rect 4136 3947 4143 4093
rect 4056 3816 4063 3820
rect 4096 3816 4103 3820
rect 3936 2966 3943 3113
rect 3996 3067 4003 3093
rect 3956 2927 3963 2993
rect 3976 2867 3983 2994
rect 3996 2807 4003 3053
rect 4016 3007 4023 3813
rect 4076 3767 4083 3783
rect 4076 3756 4093 3767
rect 4080 3753 4093 3756
rect 4036 3308 4043 3533
rect 4036 3227 4043 3294
rect 4056 3147 4063 3493
rect 4096 3347 4103 3533
rect 4116 3483 4123 3773
rect 4136 3747 4143 3833
rect 4196 3787 4203 4093
rect 4216 3767 4223 4053
rect 4293 4040 4307 4053
rect 4296 4036 4303 4040
rect 4320 4003 4333 4007
rect 4316 3996 4333 4003
rect 4320 3993 4333 3996
rect 4356 3927 4363 4033
rect 4376 4006 4383 4033
rect 4416 4007 4423 4173
rect 4316 3816 4323 3913
rect 4416 3907 4423 3953
rect 4356 3787 4363 3814
rect 4116 3476 4143 3483
rect 4256 3463 4263 3753
rect 4296 3747 4303 3783
rect 4436 3707 4443 4233
rect 4456 4007 4463 4334
rect 4476 4307 4483 4376
rect 4476 4067 4483 4193
rect 4516 4167 4523 5036
rect 4576 5027 4583 5453
rect 4616 5427 4623 5993
rect 4647 5903 4660 5907
rect 4647 5896 4663 5903
rect 4696 5896 4703 6053
rect 4736 5947 4743 6634
rect 4756 6247 4763 6693
rect 4776 6367 4783 6634
rect 4796 6607 4803 6673
rect 4816 6567 4823 6653
rect 4836 6606 4843 6773
rect 4896 6767 4903 7933
rect 4913 7927 4927 7940
rect 4956 7827 4963 7943
rect 5036 7847 5043 7973
rect 4933 7680 4947 7693
rect 4936 7676 4943 7680
rect 4936 7456 4943 7613
rect 4956 7587 4963 7643
rect 4976 7487 4983 7593
rect 4996 7527 5003 7833
rect 5036 7647 5043 7812
rect 5056 7767 5063 7953
rect 5076 7946 5083 7973
rect 4973 7460 4987 7473
rect 4976 7456 4983 7460
rect 5056 7463 5063 7753
rect 5076 7527 5083 7773
rect 5096 7567 5103 8136
rect 5216 8123 5223 8513
rect 5207 8116 5223 8123
rect 5136 7988 5143 8053
rect 5176 7988 5183 8033
rect 5196 8007 5203 8113
rect 5176 7887 5183 7913
rect 5196 7887 5203 7943
rect 5116 7688 5123 7773
rect 5136 7727 5143 7793
rect 5136 7676 5143 7713
rect 5047 7456 5063 7463
rect 5036 7426 5043 7453
rect 4956 7420 4963 7423
rect 4953 7407 4967 7420
rect 5056 7343 5063 7432
rect 5056 7336 5083 7343
rect 4916 7107 4923 7193
rect 4936 7147 4943 7273
rect 5036 7267 5043 7333
rect 5056 7287 5063 7313
rect 4996 7156 5003 7253
rect 4976 7120 4983 7123
rect 4973 7107 4987 7120
rect 4916 6906 4923 7093
rect 4936 7007 4943 7073
rect 4953 6967 4967 6973
rect 5036 6967 5043 7073
rect 4953 6960 4973 6967
rect 4956 6953 4973 6960
rect 5056 6963 5063 7053
rect 5076 7007 5083 7336
rect 5096 7327 5103 7553
rect 5056 6956 5083 6963
rect 4956 6936 4963 6953
rect 5056 6903 5063 6933
rect 4896 6648 4903 6693
rect 4936 6636 4943 6713
rect 4976 6607 4983 6903
rect 5016 6900 5023 6903
rect 5013 6887 5027 6900
rect 5036 6896 5063 6903
rect 5016 6807 5023 6833
rect 5016 6607 5023 6753
rect 4776 6007 4783 6293
rect 4796 6107 4803 6383
rect 4647 5893 4660 5896
rect 4636 5467 4643 5853
rect 4776 5863 4783 5894
rect 4656 5807 4663 5833
rect 4716 5767 4723 5863
rect 4756 5856 4783 5863
rect 4676 5387 4683 5533
rect 4696 5487 4703 5713
rect 4756 5596 4763 5856
rect 4796 5667 4803 6093
rect 4816 5727 4823 6013
rect 4776 5560 4783 5563
rect 4773 5547 4787 5560
rect 4836 5527 4843 6513
rect 4876 6116 4883 6393
rect 4916 6380 4923 6383
rect 4913 6367 4927 6380
rect 4916 6287 4923 6353
rect 4913 6120 4927 6133
rect 4916 6116 4923 6120
rect 4956 6116 4963 6233
rect 4996 6187 5003 6533
rect 5016 6287 5023 6572
rect 4896 5967 4903 6083
rect 4936 5987 4943 6083
rect 4996 5967 5003 6114
rect 4936 5896 4943 5952
rect 5016 5927 5023 6273
rect 4956 5767 4963 5863
rect 5016 5767 5023 5892
rect 4967 5756 4983 5763
rect 4976 5596 4983 5756
rect 5036 5747 5043 6896
rect 5056 6767 5063 6873
rect 5056 6087 5063 6732
rect 5076 6727 5083 6956
rect 5096 6687 5103 7133
rect 5116 6707 5123 7633
rect 5196 7487 5203 7633
rect 5216 7567 5223 7853
rect 5236 7607 5243 8533
rect 5256 8407 5263 8913
rect 5276 8847 5283 8972
rect 5296 8967 5303 9153
rect 5316 8716 5323 9171
rect 5396 9167 5403 9473
rect 5416 9267 5423 9503
rect 5456 9467 5463 9503
rect 5436 9207 5443 9253
rect 5456 9206 5463 9393
rect 5476 9187 5483 9253
rect 5496 9248 5503 9373
rect 5536 9347 5543 10032
rect 5556 9967 5563 10356
rect 5656 10276 5663 10313
rect 5576 10107 5583 10274
rect 5556 9307 5563 9833
rect 5576 9407 5583 10054
rect 5596 9687 5603 10233
rect 5636 10227 5643 10243
rect 5627 10216 5643 10227
rect 5627 10213 5640 10216
rect 5696 10056 5703 10693
rect 5716 10287 5723 10752
rect 5736 10247 5743 11133
rect 5796 11063 5803 11243
rect 5796 11056 5823 11063
rect 5796 10796 5823 10803
rect 5796 10727 5803 10796
rect 5856 10687 5863 10763
rect 5767 10583 5780 10587
rect 5767 10576 5783 10583
rect 5816 10576 5823 10613
rect 5767 10573 5780 10576
rect 5896 10543 5903 11243
rect 5796 10427 5803 10532
rect 5616 9543 5623 10053
rect 5676 9967 5683 10023
rect 5716 10007 5723 10023
rect 5716 9867 5723 9993
rect 5776 9987 5783 10393
rect 5836 10367 5843 10543
rect 5876 10536 5903 10543
rect 5693 9767 5707 9773
rect 5656 9667 5663 9723
rect 5656 9548 5663 9573
rect 5716 9567 5723 9712
rect 5596 9536 5623 9543
rect 5556 9236 5563 9293
rect 5596 9287 5603 9536
rect 5593 9240 5607 9252
rect 5596 9236 5603 9240
rect 5356 9016 5363 9093
rect 5393 9028 5407 9033
rect 5336 8687 5343 8973
rect 5276 8567 5283 8683
rect 5356 8627 5363 8953
rect 5416 8787 5423 8983
rect 5256 8167 5263 8393
rect 5276 8387 5283 8553
rect 5296 8287 5303 8473
rect 5316 8447 5323 8613
rect 5356 8496 5363 8573
rect 5376 8527 5383 8733
rect 5396 8607 5403 8653
rect 5416 8567 5423 8633
rect 5436 8627 5443 8714
rect 5396 8496 5403 8533
rect 5456 8467 5463 9153
rect 5476 8747 5483 8972
rect 5496 8927 5503 9234
rect 5576 9200 5583 9203
rect 5573 9187 5587 9200
rect 5516 8947 5523 9093
rect 5636 9067 5643 9273
rect 5656 9187 5663 9433
rect 5696 9387 5703 9534
rect 5696 9207 5703 9333
rect 5716 9183 5723 9553
rect 5736 9207 5743 9793
rect 5756 9407 5763 9853
rect 5776 9347 5783 9853
rect 5796 9447 5803 10313
rect 5876 10276 5883 10536
rect 5836 9767 5843 10243
rect 5896 9783 5903 10473
rect 5916 10056 5923 10953
rect 5936 10327 5943 11094
rect 5956 10083 5963 10573
rect 5976 10527 5983 11243
rect 6036 11096 6043 11133
rect 6076 11057 6083 11243
rect 6236 11096 6263 11103
rect 6056 10808 6063 10833
rect 6096 10796 6103 10873
rect 6156 10767 6163 10794
rect 6076 10540 6083 10543
rect 5976 10246 5983 10333
rect 5956 10076 5983 10083
rect 5876 9776 5903 9783
rect 5876 9768 5883 9776
rect 5916 9756 5923 9793
rect 5816 9627 5823 9753
rect 5856 9720 5863 9723
rect 5836 9687 5843 9713
rect 5853 9707 5867 9720
rect 5896 9687 5903 9723
rect 5833 9540 5847 9553
rect 5836 9536 5843 9540
rect 5876 9536 5883 9673
rect 5900 9503 5913 9507
rect 5896 9496 5913 9503
rect 5900 9493 5913 9496
rect 5856 9327 5863 9492
rect 5876 9207 5883 9353
rect 5696 9176 5723 9183
rect 5596 9016 5603 9053
rect 5656 8976 5683 8983
rect 5513 8720 5527 8733
rect 5516 8716 5523 8720
rect 5487 8683 5500 8687
rect 5487 8676 5503 8683
rect 5487 8673 5500 8676
rect 5376 8443 5383 8463
rect 5536 8463 5543 8613
rect 5596 8496 5603 8753
rect 5636 8687 5643 8933
rect 5656 8627 5663 8953
rect 5536 8456 5563 8463
rect 5376 8436 5403 8443
rect 5316 8196 5323 8393
rect 5256 7467 5263 8132
rect 5296 8087 5303 8163
rect 5276 7847 5283 7974
rect 5296 7927 5303 7993
rect 5136 6906 5143 7373
rect 5156 7227 5163 7423
rect 5176 7347 5183 7393
rect 5196 7167 5203 7423
rect 5276 7367 5283 7673
rect 5296 7367 5303 7913
rect 5316 7687 5323 8093
rect 5336 7723 5343 8153
rect 5356 8107 5363 8433
rect 5376 8247 5383 8313
rect 5356 7987 5363 8053
rect 5376 7976 5383 8233
rect 5396 8067 5403 8436
rect 5416 8307 5423 8452
rect 5416 8127 5423 8293
rect 5456 8047 5463 8373
rect 5516 8196 5523 8293
rect 5476 8156 5503 8163
rect 5413 7980 5427 7993
rect 5416 7976 5423 7980
rect 5396 7940 5403 7943
rect 5356 7907 5363 7933
rect 5393 7927 5407 7940
rect 5336 7716 5353 7723
rect 5356 7676 5363 7713
rect 5416 7687 5423 7893
rect 5436 7843 5443 7943
rect 5476 7867 5483 8156
rect 5436 7836 5463 7843
rect 5336 7547 5343 7643
rect 5413 7627 5427 7633
rect 5356 7387 5363 7613
rect 5436 7607 5443 7674
rect 5416 7456 5423 7592
rect 5456 7467 5463 7836
rect 5336 7207 5343 7313
rect 5176 7027 5183 7154
rect 5253 7160 5267 7173
rect 5256 7156 5263 7160
rect 5193 7107 5207 7113
rect 5316 7123 5323 7173
rect 5336 7126 5343 7193
rect 5296 7116 5323 7123
rect 5207 6993 5213 7007
rect 5173 6940 5187 6953
rect 5176 6936 5183 6940
rect 5196 6807 5203 6903
rect 5176 6636 5183 6713
rect 5196 6648 5203 6673
rect 5076 6487 5083 6634
rect 5156 6600 5163 6603
rect 5153 6587 5167 6600
rect 5236 6547 5243 6973
rect 5256 6523 5263 7073
rect 5276 6967 5283 6993
rect 5296 6987 5303 7116
rect 5356 7087 5363 7352
rect 5376 7067 5383 7353
rect 5396 7127 5403 7412
rect 5436 7387 5443 7423
rect 5456 7367 5463 7413
rect 5316 6967 5323 6993
rect 5416 6983 5423 7353
rect 5476 7168 5483 7713
rect 5496 7427 5503 8013
rect 5516 7607 5523 8073
rect 5536 7627 5543 8093
rect 5556 8087 5563 8456
rect 5576 8407 5583 8463
rect 5616 8447 5623 8463
rect 5576 8227 5583 8372
rect 5576 8087 5583 8213
rect 5596 8147 5603 8413
rect 5616 8307 5623 8433
rect 5556 7847 5563 8033
rect 5616 8027 5623 8253
rect 5636 8027 5643 8273
rect 5613 7980 5627 7992
rect 5656 7987 5663 8453
rect 5616 7976 5623 7980
rect 5636 7647 5643 7773
rect 5536 7227 5543 7473
rect 5456 7047 5463 7123
rect 5496 7087 5503 7123
rect 5447 6993 5453 7007
rect 5476 7003 5483 7053
rect 5476 6996 5503 7003
rect 5416 6976 5443 6983
rect 5276 6667 5283 6813
rect 5296 6547 5303 6773
rect 5236 6516 5263 6523
rect 5116 6447 5123 6473
rect 5107 6423 5120 6427
rect 5107 6416 5123 6423
rect 5107 6413 5120 6416
rect 5136 6380 5143 6383
rect 5133 6367 5147 6380
rect 5216 6367 5223 6433
rect 5236 6367 5243 6516
rect 5316 6507 5323 6953
rect 5393 6940 5407 6953
rect 5396 6936 5403 6940
rect 5436 6936 5443 6976
rect 5376 6707 5383 6892
rect 5396 6687 5403 6833
rect 5416 6727 5423 6903
rect 5456 6607 5463 6713
rect 5476 6707 5483 6973
rect 5476 6607 5483 6634
rect 5356 6600 5363 6603
rect 5353 6587 5367 6600
rect 5496 6606 5503 6996
rect 5516 6947 5523 7053
rect 5536 6903 5543 7113
rect 5556 7087 5563 7333
rect 5576 7203 5583 7593
rect 5636 7456 5643 7612
rect 5656 7527 5663 7713
rect 5676 7627 5683 8976
rect 5696 8643 5703 9176
rect 5736 8907 5743 9172
rect 5756 8967 5763 9193
rect 5816 9187 5823 9203
rect 5816 9176 5833 9187
rect 5820 9173 5833 9176
rect 5816 9016 5823 9153
rect 5853 9020 5867 9033
rect 5896 9027 5903 9473
rect 5856 9016 5863 9020
rect 5836 8947 5843 8983
rect 5760 8743 5773 8747
rect 5756 8733 5773 8743
rect 5756 8716 5763 8733
rect 5776 8680 5783 8683
rect 5773 8667 5787 8680
rect 5696 8636 5713 8643
rect 5696 8387 5703 8612
rect 5716 8508 5723 8633
rect 5716 8447 5723 8494
rect 5716 8227 5723 8333
rect 5736 8267 5743 8651
rect 5816 8647 5823 8893
rect 5756 8467 5763 8494
rect 5776 8347 5783 8632
rect 5856 8623 5863 8953
rect 5876 8907 5883 8983
rect 5876 8827 5883 8893
rect 5836 8616 5863 8623
rect 5836 8587 5843 8616
rect 5876 8607 5883 8713
rect 5896 8687 5903 8973
rect 5856 8496 5863 8553
rect 5836 8460 5843 8463
rect 5833 8447 5847 8460
rect 5756 8196 5783 8203
rect 5716 8127 5723 8163
rect 5776 8147 5783 8196
rect 5696 7647 5703 7973
rect 5576 7196 5603 7203
rect 5576 7063 5583 7154
rect 5596 7127 5603 7196
rect 5616 7127 5623 7423
rect 5716 7407 5723 8013
rect 5736 7387 5743 8133
rect 5756 7747 5763 8113
rect 5816 7976 5823 8353
rect 5836 8067 5843 8194
rect 5856 7988 5863 8433
rect 5876 8427 5883 8463
rect 5876 8147 5883 8373
rect 5916 8367 5923 9433
rect 5936 9067 5943 9393
rect 5936 8847 5943 9013
rect 5956 8947 5963 9973
rect 5976 8887 5983 10076
rect 5996 10027 6003 10532
rect 6073 10527 6087 10540
rect 6116 10487 6123 10713
rect 6196 10687 6203 10752
rect 6176 10587 6183 10613
rect 6196 10427 6203 10673
rect 6076 10276 6083 10413
rect 6116 10276 6123 10373
rect 5996 9287 6003 10013
rect 6016 9487 6023 10273
rect 6196 10247 6203 10413
rect 6136 10207 6143 10243
rect 6216 10127 6223 10733
rect 6236 10463 6243 11096
rect 6296 11057 6303 11243
rect 6316 10796 6323 11033
rect 6296 10760 6303 10763
rect 6293 10747 6307 10760
rect 6396 10747 6403 11243
rect 6496 11096 6503 11173
rect 6416 10747 6423 11094
rect 6556 11063 6563 11093
rect 6476 11060 6483 11063
rect 6473 11047 6487 11060
rect 6516 11056 6563 11063
rect 6296 10576 6303 10693
rect 6256 10487 6263 10543
rect 6236 10456 6263 10463
rect 6156 10056 6163 10113
rect 6056 9707 6063 10012
rect 6176 9987 6183 10023
rect 6136 9756 6143 9873
rect 6116 9647 6123 9723
rect 6036 9236 6043 9493
rect 6076 9443 6083 9503
rect 6076 9436 6103 9443
rect 6016 9200 6023 9203
rect 5996 8927 6003 9193
rect 6013 9187 6027 9200
rect 5953 8720 5967 8733
rect 5956 8716 5963 8720
rect 5996 8716 6003 8813
rect 6016 8767 6023 9152
rect 6076 9043 6083 9413
rect 6096 9387 6103 9436
rect 6116 9167 6123 9493
rect 6136 9467 6143 9534
rect 6056 9036 6083 9043
rect 6056 9016 6063 9036
rect 6096 9016 6103 9153
rect 6116 8963 6123 8983
rect 6087 8956 6123 8963
rect 6016 8647 6023 8683
rect 5956 8287 5963 8533
rect 5996 8387 6003 8533
rect 5976 8227 5983 8293
rect 5896 8127 5903 8213
rect 6016 8163 6023 8573
rect 6056 8547 6063 8913
rect 6076 8547 6083 8733
rect 6096 8667 6103 8733
rect 6073 8523 6087 8533
rect 6056 8520 6087 8523
rect 6056 8516 6083 8520
rect 6056 8496 6063 8516
rect 6096 8507 6103 8593
rect 6116 8587 6123 8933
rect 6136 8687 6143 8973
rect 6136 8467 6143 8652
rect 6080 8464 6093 8467
rect 6076 8457 6093 8464
rect 6080 8453 6093 8457
rect 6156 8447 6163 9713
rect 6176 9307 6183 9653
rect 6196 9507 6203 9993
rect 6216 9767 6223 10023
rect 6256 9727 6263 10456
rect 6356 10276 6363 10733
rect 6456 10687 6463 10873
rect 6496 10766 6503 10853
rect 6556 10796 6563 10833
rect 6596 10796 6603 11133
rect 6696 10947 6703 11063
rect 6736 11060 6743 11063
rect 6733 11047 6747 11060
rect 6813 10800 6827 10813
rect 6816 10796 6823 10800
rect 6536 10687 6543 10763
rect 6576 10760 6583 10763
rect 6573 10747 6587 10760
rect 6636 10747 6643 10794
rect 6736 10687 6743 10794
rect 6276 9727 6283 10073
rect 6316 10007 6323 10243
rect 6376 10223 6383 10673
rect 6476 10587 6483 10633
rect 6656 10576 6703 10583
rect 6736 10576 6743 10613
rect 6536 10447 6543 10543
rect 6356 10216 6383 10223
rect 6356 10007 6363 10216
rect 6396 10087 6403 10232
rect 6393 10060 6407 10073
rect 6396 10056 6403 10060
rect 6353 9760 6367 9773
rect 6356 9756 6363 9760
rect 6296 9536 6303 9713
rect 6336 9536 6343 9573
rect 6376 9527 6383 9673
rect 6236 9236 6243 9492
rect 6176 8807 6183 9234
rect 6276 9203 6283 9433
rect 6316 9387 6323 9503
rect 6216 9167 6223 9203
rect 6256 9196 6283 9203
rect 6196 8847 6203 8873
rect 6216 8807 6223 9053
rect 6236 8867 6243 9173
rect 6256 8987 6263 9196
rect 6296 9067 6303 9353
rect 6336 9187 6343 9473
rect 6376 9403 6383 9513
rect 6396 9447 6403 9993
rect 6416 9727 6423 9754
rect 6356 9396 6383 9403
rect 6296 8827 6303 8983
rect 6207 8736 6243 8743
rect 6236 8716 6243 8736
rect 6236 8508 6243 8613
rect 6256 8607 6263 8683
rect 6296 8647 6303 8792
rect 6293 8547 6307 8553
rect 6273 8500 6287 8513
rect 6276 8496 6283 8500
rect 5936 8160 5943 8163
rect 5976 8160 5983 8163
rect 5933 8147 5947 8160
rect 5973 8147 5987 8160
rect 5996 8156 6023 8163
rect 5896 7943 5903 7993
rect 5836 7907 5843 7943
rect 5876 7940 5903 7943
rect 5873 7936 5903 7940
rect 5873 7927 5887 7936
rect 5796 7688 5803 7893
rect 5836 7676 5843 7713
rect 5896 7647 5903 7813
rect 5776 7427 5783 7632
rect 5916 7627 5923 7974
rect 5527 6896 5543 6903
rect 5556 7056 5583 7063
rect 5256 6428 5263 6493
rect 4596 5376 4623 5383
rect 4596 5287 4603 5376
rect 4736 5356 4743 5473
rect 4756 5407 4763 5513
rect 4896 5487 4903 5593
rect 4996 5543 5003 5552
rect 4947 5536 5003 5543
rect 4856 5360 4863 5363
rect 4853 5347 4867 5360
rect 4536 4887 4543 5013
rect 4556 4836 4563 4933
rect 4596 4847 4603 5113
rect 4616 4927 4623 5032
rect 4616 4836 4623 4913
rect 4536 4267 4543 4793
rect 4636 4787 4643 5293
rect 4696 5287 4703 5323
rect 4696 5247 4703 5273
rect 4756 5223 4763 5333
rect 4996 5307 5003 5513
rect 5036 5356 5043 5653
rect 5056 5627 5063 5913
rect 5056 5507 5063 5592
rect 5076 5483 5083 6313
rect 5136 6116 5143 6273
rect 5096 5527 5103 6072
rect 5156 5896 5163 5953
rect 5116 5807 5123 5893
rect 5216 5866 5223 6113
rect 5116 5627 5123 5793
rect 5176 5647 5183 5863
rect 5236 5847 5243 6353
rect 5173 5600 5187 5612
rect 5176 5596 5183 5600
rect 5256 5607 5263 6414
rect 5296 6387 5303 6453
rect 5356 6416 5363 6533
rect 5393 6420 5407 6433
rect 5436 6427 5443 6593
rect 5396 6416 5403 6420
rect 5276 5787 5283 6233
rect 5296 5847 5303 6173
rect 5316 6127 5323 6413
rect 5376 6380 5383 6383
rect 5416 6380 5423 6383
rect 5373 6367 5387 6380
rect 5413 6367 5427 6380
rect 5313 6067 5327 6073
rect 5416 5967 5423 6092
rect 5436 5927 5443 6013
rect 5456 6007 5463 6572
rect 5476 6227 5483 6572
rect 5476 6100 5483 6103
rect 5473 6087 5487 6100
rect 5456 5907 5463 5972
rect 5476 5967 5483 6073
rect 5516 5867 5523 6892
rect 5536 6567 5543 6693
rect 5556 6587 5563 7056
rect 5576 6967 5583 7033
rect 5596 7007 5603 7092
rect 5616 7047 5623 7073
rect 5636 6987 5643 7253
rect 5656 7067 5663 7373
rect 5696 7120 5703 7123
rect 5693 7107 5707 7120
rect 5633 6940 5647 6952
rect 5636 6936 5643 6940
rect 5656 6867 5663 6903
rect 5616 6727 5623 6813
rect 5616 6636 5623 6713
rect 5536 6267 5543 6493
rect 5596 6447 5603 6592
rect 5636 6423 5643 6603
rect 5696 6527 5703 7013
rect 5616 6416 5643 6423
rect 5596 6247 5603 6383
rect 5716 6267 5723 6634
rect 5736 6387 5743 7113
rect 5576 5896 5583 5993
rect 5296 5787 5303 5812
rect 5336 5687 5343 5863
rect 5376 5860 5383 5863
rect 5373 5847 5387 5860
rect 5556 5827 5563 5863
rect 5296 5627 5303 5673
rect 5056 5476 5083 5483
rect 4756 5216 4783 5223
rect 4676 5076 4683 5113
rect 4696 5040 4703 5043
rect 4693 5027 4707 5040
rect 4667 5023 4680 5027
rect 4667 5013 4683 5023
rect 4596 4336 4603 4773
rect 4656 4667 4663 4992
rect 4676 4963 4683 5013
rect 4736 4967 4743 5043
rect 4776 5027 4783 5216
rect 4796 5067 4803 5153
rect 4676 4956 4703 4963
rect 4676 4787 4683 4933
rect 4696 4556 4703 4956
rect 4716 4727 4723 4933
rect 4816 4907 4823 5193
rect 4836 4856 4843 5233
rect 4856 4947 4863 5273
rect 5056 5247 5063 5476
rect 5096 5356 5103 5453
rect 5116 5303 5123 5573
rect 5136 5467 5143 5594
rect 5196 5407 5203 5563
rect 5276 5563 5283 5583
rect 5316 5566 5323 5633
rect 5516 5576 5523 5733
rect 5536 5587 5543 5633
rect 5256 5556 5283 5563
rect 5256 5543 5263 5556
rect 5227 5536 5263 5543
rect 5216 5447 5223 5493
rect 5316 5403 5323 5513
rect 5336 5427 5343 5572
rect 5316 5396 5343 5403
rect 5116 5296 5143 5303
rect 4876 4987 4883 5153
rect 4936 5076 4943 5213
rect 4956 5040 4963 5043
rect 4916 4903 4923 5032
rect 4953 5027 4967 5040
rect 4996 5007 5003 5113
rect 4916 4896 4943 4903
rect 4867 4853 4873 4867
rect 4676 4343 4683 4523
rect 4676 4336 4703 4343
rect 4556 4287 4563 4334
rect 4573 4287 4587 4292
rect 4567 4193 4573 4207
rect 4676 4147 4683 4173
rect 4696 4147 4703 4336
rect 4716 4227 4723 4512
rect 4756 4287 4763 4833
rect 4776 4287 4783 4812
rect 4836 4368 4843 4593
rect 4856 4527 4863 4573
rect 4893 4560 4907 4573
rect 4936 4568 4943 4896
rect 4956 4868 4963 4973
rect 5016 4947 5023 5193
rect 5136 5147 5143 5296
rect 5036 5047 5043 5133
rect 5196 5108 5203 5393
rect 5336 5376 5343 5396
rect 5536 5376 5543 5453
rect 5236 5096 5243 5253
rect 5256 5167 5263 5374
rect 5356 5207 5363 5343
rect 5556 5287 5563 5343
rect 5376 5227 5383 5253
rect 5040 5026 5060 5027
rect 5047 5013 5053 5026
rect 5076 4987 5083 5093
rect 4996 4896 5063 4903
rect 4996 4867 5003 4896
rect 4956 4607 4963 4854
rect 5013 4860 5027 4873
rect 5016 4856 5023 4860
rect 5056 4856 5063 4896
rect 5096 4863 5103 5093
rect 5153 5080 5167 5093
rect 5156 5076 5163 5080
rect 5116 4887 5123 5033
rect 5176 5040 5183 5043
rect 5173 5027 5187 5040
rect 5256 5007 5263 5053
rect 5096 4856 5123 4863
rect 5036 4767 5043 4823
rect 4896 4556 4903 4560
rect 4876 4336 4883 4393
rect 4896 4347 4903 4473
rect 4556 4107 4563 4133
rect 4473 3907 4487 3913
rect 4473 3900 4493 3907
rect 4476 3896 4493 3900
rect 4480 3893 4493 3896
rect 4476 3707 4483 3873
rect 4236 3456 4263 3463
rect 4176 3347 4183 3443
rect 4136 3296 4143 3333
rect 4096 3163 4103 3233
rect 4116 3183 4123 3252
rect 4176 3247 4183 3333
rect 4116 3176 4143 3183
rect 4096 3156 4123 3163
rect 4036 3087 4043 3113
rect 4036 3027 4043 3052
rect 4076 3027 4083 3053
rect 4096 2996 4103 3133
rect 4116 3007 4123 3156
rect 4136 3087 4143 3176
rect 4016 2867 4023 2893
rect 4036 2767 4043 2793
rect 3956 2740 3963 2743
rect 3896 2027 3903 2293
rect 3916 1967 3923 2733
rect 3953 2727 3967 2740
rect 3996 2723 4003 2743
rect 3976 2716 4003 2723
rect 3936 2423 3943 2474
rect 3936 2416 3963 2423
rect 3736 1827 3743 1953
rect 3916 1926 3923 1953
rect 3656 1587 3663 1613
rect 3676 1547 3683 1593
rect 3716 1567 3723 1703
rect 3776 1587 3783 1753
rect 3796 1607 3803 1923
rect 3916 1887 3923 1912
rect 3896 1807 3903 1873
rect 3936 1767 3943 2193
rect 3956 2187 3963 2416
rect 3976 2407 3983 2716
rect 4056 2476 4063 2793
rect 4076 2747 4083 2963
rect 4073 2507 4087 2513
rect 4096 2487 4103 2933
rect 4116 2788 4123 2913
rect 3996 2367 4003 2432
rect 3976 2107 3983 2333
rect 4016 2303 4023 2393
rect 4036 2327 4043 2443
rect 4076 2367 4083 2432
rect 4016 2296 4043 2303
rect 4036 2256 4043 2296
rect 4096 2226 4103 2353
rect 4016 2220 4023 2223
rect 4013 2207 4027 2220
rect 4056 2147 4063 2223
rect 3996 1968 4003 2133
rect 4096 2127 4103 2212
rect 4036 1956 4043 2073
rect 3776 1547 3783 1573
rect 3773 1467 3787 1473
rect 3696 1367 3703 1403
rect 3496 1047 3503 1213
rect 3613 1167 3627 1172
rect 3547 963 3560 967
rect 3547 953 3563 963
rect 3493 920 3507 933
rect 3556 943 3563 953
rect 3556 940 3583 943
rect 3556 936 3587 940
rect 3533 920 3547 932
rect 3573 928 3587 936
rect 3496 916 3503 920
rect 3536 916 3543 920
rect 3236 696 3243 733
rect 3216 587 3223 663
rect 3136 396 3163 403
rect 3296 403 3303 883
rect 3456 886 3463 913
rect 3433 700 3447 713
rect 3436 696 3443 700
rect 3516 666 3523 872
rect 3556 447 3563 883
rect 3616 607 3623 1033
rect 3636 787 3643 1233
rect 3656 1187 3663 1214
rect 3676 947 3683 1293
rect 3696 1187 3703 1253
rect 3756 1227 3763 1393
rect 3796 1248 3803 1533
rect 3816 1467 3823 1734
rect 3996 1736 4003 1873
rect 3836 1307 3843 1553
rect 3876 1527 3883 1633
rect 3896 1443 3903 1733
rect 3916 1607 3923 1633
rect 3876 1436 3903 1443
rect 3916 1436 3923 1593
rect 3936 1487 3943 1613
rect 3976 1587 3983 1703
rect 3956 1436 3963 1493
rect 3996 1447 4003 1573
rect 4076 1547 4083 1953
rect 4136 1487 4143 3052
rect 4176 2947 4183 2993
rect 4156 2867 4163 2893
rect 4176 2807 4183 2833
rect 4196 2827 4203 3073
rect 4216 2907 4223 3294
rect 4236 2947 4243 3456
rect 4256 3227 4263 3333
rect 4276 3203 4283 3693
rect 4476 3567 4483 3613
rect 4476 3516 4483 3553
rect 4296 3347 4303 3514
rect 4333 3467 4347 3473
rect 4376 3447 4383 3514
rect 4407 3483 4420 3487
rect 4407 3480 4423 3483
rect 4407 3473 4427 3480
rect 4413 3467 4427 3473
rect 4336 3327 4343 3393
rect 4356 3296 4363 3373
rect 4396 3327 4403 3353
rect 4416 3263 4423 3333
rect 4436 3327 4443 3433
rect 4256 3196 4283 3203
rect 4256 2963 4263 3196
rect 4336 3023 4343 3263
rect 4376 3256 4423 3263
rect 4396 3147 4403 3256
rect 4416 3063 4423 3213
rect 4396 3056 4423 3063
rect 4336 3016 4363 3023
rect 4256 2956 4283 2963
rect 4256 2907 4263 2956
rect 4173 2780 4187 2793
rect 4176 2776 4183 2780
rect 4196 1967 4203 2743
rect 4216 2647 4223 2693
rect 4256 2607 4263 2793
rect 4276 2687 4283 2933
rect 4296 2746 4303 2813
rect 4316 2667 4323 2933
rect 4336 2787 4343 2973
rect 4356 2947 4363 3016
rect 4396 2966 4403 3056
rect 4436 3043 4443 3313
rect 4416 3036 4443 3043
rect 4416 2907 4423 3036
rect 4436 2927 4443 3013
rect 4396 2776 4403 2853
rect 4436 2788 4443 2813
rect 4456 2787 4463 3353
rect 4516 3303 4523 3613
rect 4536 3486 4543 3653
rect 4556 3527 4563 3783
rect 4576 3627 4583 3992
rect 4596 3947 4603 4093
rect 4536 3367 4543 3393
rect 4576 3347 4583 3513
rect 4596 3327 4603 3933
rect 4616 3527 4623 4133
rect 4796 4123 4803 4333
rect 4796 4116 4823 4123
rect 4656 3787 4663 4013
rect 4636 3363 4643 3472
rect 4676 3367 4683 3473
rect 4636 3356 4663 3363
rect 4496 3296 4523 3303
rect 4496 3027 4503 3296
rect 4616 3303 4623 3333
rect 4596 3296 4623 3303
rect 4516 3207 4523 3273
rect 4576 3243 4583 3263
rect 4556 3236 4583 3243
rect 4516 2996 4523 3113
rect 4556 3067 4563 3236
rect 4216 2547 4223 2573
rect 4276 2547 4283 2633
rect 4353 2627 4367 2633
rect 4316 2587 4323 2613
rect 4416 2527 4423 2743
rect 4247 2513 4253 2527
rect 4296 2476 4303 2513
rect 4216 2327 4223 2474
rect 4276 2367 4283 2443
rect 4316 2436 4343 2443
rect 4296 2347 4303 2413
rect 4336 2367 4343 2436
rect 4256 2307 4263 2333
rect 4296 2256 4303 2333
rect 4236 2187 4243 2223
rect 4336 2183 4343 2353
rect 4356 2226 4363 2473
rect 4336 2176 4353 2183
rect 4176 1927 4183 1954
rect 4236 1956 4243 2013
rect 4216 1887 4223 1923
rect 4176 1736 4183 1813
rect 4256 1748 4263 1923
rect 4196 1607 4203 1703
rect 4156 1547 4163 1573
rect 3856 1267 3863 1433
rect 3876 1406 3883 1436
rect 3833 1220 3847 1233
rect 3876 1227 3883 1333
rect 3836 1216 3843 1220
rect 3816 1127 3823 1183
rect 3696 886 3703 1053
rect 3776 916 3783 1033
rect 3816 1007 3823 1113
rect 3876 1067 3883 1133
rect 3696 607 3703 663
rect 3616 487 3623 593
rect 3836 547 3843 953
rect 3896 847 3903 1253
rect 3916 1167 3923 1193
rect 3936 1107 3943 1392
rect 4016 1367 4023 1453
rect 3956 1167 3963 1233
rect 4096 1223 4103 1433
rect 4136 1327 4143 1403
rect 4096 1216 4123 1223
rect 4116 1186 4123 1216
rect 4036 1127 4043 1183
rect 3967 883 3980 887
rect 4056 886 4063 1133
rect 3967 876 3983 883
rect 3967 873 3980 876
rect 4136 787 4143 1213
rect 4216 967 4223 1453
rect 4236 1183 4243 1313
rect 4256 1267 4263 1473
rect 4276 1216 4283 1293
rect 4336 1223 4343 1813
rect 4356 1436 4363 2173
rect 4376 2087 4383 2393
rect 4416 2107 4423 2313
rect 4456 2307 4463 2733
rect 4476 2487 4483 2893
rect 4496 2476 4503 2773
rect 4556 2747 4563 3013
rect 4536 2476 4543 2673
rect 4576 2507 4583 3213
rect 4636 3187 4643 3333
rect 4656 2907 4663 3356
rect 4696 3343 4703 3973
rect 4716 3947 4723 4003
rect 4796 3987 4803 4034
rect 4816 3947 4823 4116
rect 4716 3828 4723 3933
rect 4836 3927 4843 4273
rect 4736 3816 4743 3913
rect 4776 3816 4783 3853
rect 4756 3747 4763 3783
rect 4796 3607 4803 3783
rect 4856 3747 4863 4213
rect 4876 4048 4883 4173
rect 4916 4043 4923 4353
rect 4936 4147 4943 4453
rect 4976 4287 4983 4393
rect 5056 4336 5063 4653
rect 5116 4607 5123 4856
rect 5136 4647 5143 4973
rect 5276 4947 5283 5063
rect 5296 4927 5303 5113
rect 5396 5056 5403 5133
rect 5556 5103 5563 5273
rect 5536 5096 5563 5103
rect 5536 4967 5543 5096
rect 5576 5027 5583 5063
rect 5347 4893 5353 4907
rect 5136 4516 5163 4523
rect 5096 4336 5103 4453
rect 5156 4348 5163 4516
rect 5016 4306 5023 4333
rect 5076 4300 5083 4303
rect 5073 4287 5087 4300
rect 4896 4036 4923 4043
rect 4896 4006 4903 4036
rect 4976 4036 4983 4252
rect 5056 4167 5063 4253
rect 5156 4247 5163 4334
rect 4893 3987 4907 3992
rect 4916 3927 4923 3953
rect 4916 3707 4923 3813
rect 4676 3336 4703 3343
rect 4676 3087 4683 3336
rect 4696 3027 4703 3293
rect 4716 3266 4723 3573
rect 4736 3486 4743 3513
rect 4756 3487 4763 3553
rect 4836 3547 4843 3573
rect 4776 3467 4783 3533
rect 4856 3516 4863 3633
rect 4896 3567 4903 3693
rect 4736 3227 4743 3313
rect 4836 3296 4843 3353
rect 4856 3308 4863 3393
rect 4816 3227 4823 3263
rect 4716 2996 4723 3153
rect 4776 2963 4783 3013
rect 4696 2847 4703 2963
rect 4736 2956 4783 2963
rect 4733 2847 4747 2853
rect 4616 2723 4623 2743
rect 4616 2716 4643 2723
rect 4596 2446 4603 2473
rect 4516 2387 4523 2443
rect 4536 2256 4543 2353
rect 4436 2226 4443 2253
rect 4436 1956 4443 1993
rect 4476 1956 4483 2153
rect 4436 1736 4443 1853
rect 4456 1827 4463 1923
rect 4476 1847 4483 1893
rect 4496 1887 4503 1923
rect 4536 1887 4543 2073
rect 4476 1716 4483 1773
rect 4396 1400 4403 1403
rect 4393 1387 4407 1400
rect 4336 1216 4363 1223
rect 4333 1183 4347 1193
rect 4236 1176 4263 1183
rect 4316 1180 4347 1183
rect 4316 1176 4343 1180
rect 4356 1047 4363 1216
rect 4213 920 4227 932
rect 4216 916 4223 920
rect 4256 916 4263 953
rect 4156 847 4163 913
rect 3876 696 3883 733
rect 4116 696 4123 733
rect 3896 660 3903 663
rect 3893 647 3907 660
rect 4096 627 4103 663
rect 4136 627 4143 663
rect 3276 396 3303 403
rect 3356 396 3363 433
rect 3420 423 3433 427
rect 3416 413 3433 423
rect 3416 396 3423 413
rect 2916 147 2923 174
rect 2856 127 2863 143
rect 3196 146 3203 393
rect 3233 347 3247 353
rect 3256 307 3263 333
rect 3256 176 3263 272
rect 3276 227 3283 396
rect 3316 360 3323 363
rect 3313 347 3327 360
rect 3296 247 3303 313
rect 3376 287 3383 363
rect 3556 287 3563 412
rect 3576 366 3583 453
rect 3956 427 3963 473
rect 4196 447 4203 883
rect 4236 847 4243 883
rect 3687 413 3693 427
rect 3720 423 3733 427
rect 3716 413 3733 423
rect 3716 396 3723 413
rect 3913 400 3927 413
rect 3953 400 3967 413
rect 3916 396 3923 400
rect 3956 396 3963 400
rect 3676 327 3683 363
rect 3736 327 3743 373
rect 3756 247 3763 293
rect 3316 143 3323 174
rect 3956 176 3963 233
rect 4096 188 4103 433
rect 4176 360 4183 363
rect 4173 347 4187 360
rect 4216 347 4223 693
rect 4296 627 4303 913
rect 4316 847 4323 933
rect 4376 747 4383 913
rect 4396 886 4403 1213
rect 4416 927 4423 1703
rect 4436 1327 4443 1393
rect 4456 1227 4463 1693
rect 4476 1216 4483 1513
rect 4516 1248 4523 1813
rect 4576 1783 4583 2253
rect 4596 1847 4603 2432
rect 4616 1827 4623 2493
rect 4636 2047 4643 2716
rect 4656 2147 4663 2743
rect 4676 2367 4683 2473
rect 4676 2226 4683 2353
rect 4696 2267 4703 2773
rect 4756 2746 4763 2893
rect 4796 2847 4803 2893
rect 4816 2887 4823 3173
rect 4727 2713 4733 2727
rect 4716 2487 4723 2593
rect 4776 2507 4783 2833
rect 4816 2787 4823 2852
rect 4836 2827 4843 3233
rect 4896 3187 4903 3453
rect 4916 3207 4923 3373
rect 4936 3287 4943 3973
rect 4953 3967 4967 3971
rect 4996 3907 5003 4003
rect 5036 3816 5043 3933
rect 5056 3827 5063 4153
rect 4956 3667 4963 3773
rect 4956 3407 4963 3514
rect 4976 3467 4983 3783
rect 4996 3367 5003 3733
rect 5076 3627 5083 4133
rect 5096 3567 5103 4233
rect 5176 4227 5183 4873
rect 5196 4167 5203 4893
rect 5216 4826 5223 4893
rect 5276 4803 5283 4823
rect 5256 4796 5283 4803
rect 5236 4447 5243 4713
rect 5256 4267 5263 4796
rect 5293 4560 5307 4573
rect 5296 4556 5303 4560
rect 5336 4556 5343 4753
rect 5356 4667 5363 4872
rect 5376 4787 5383 4853
rect 5376 4556 5383 4613
rect 5296 4336 5303 4413
rect 5316 4367 5323 4512
rect 5356 4427 5363 4523
rect 5356 4307 5363 4353
rect 5256 4036 5263 4073
rect 5116 4007 5123 4034
rect 5156 4003 5163 4034
rect 5296 4007 5303 4133
rect 5156 3996 5183 4003
rect 5016 3487 5023 3514
rect 5036 3427 5043 3553
rect 5116 3516 5123 3813
rect 5156 3687 5163 3893
rect 5053 3308 5067 3313
rect 4936 3087 4943 3233
rect 4956 3187 4963 3293
rect 5096 3267 5103 3333
rect 5036 3247 5043 3263
rect 4896 3008 4903 3073
rect 4876 2996 4893 3003
rect 4876 2947 4883 2996
rect 4973 3000 4987 3013
rect 4976 2996 4983 3000
rect 5016 2966 5023 3173
rect 4836 2776 4843 2813
rect 4856 2807 4863 2893
rect 4896 2867 4903 2893
rect 4876 2776 4883 2853
rect 4796 2723 4803 2773
rect 4956 2746 4963 2963
rect 4796 2716 4823 2723
rect 4796 2647 4803 2693
rect 4816 2687 4823 2716
rect 4816 2446 4823 2673
rect 4836 2667 4843 2713
rect 4896 2687 4903 2743
rect 4916 2587 4923 2693
rect 4736 2347 4743 2443
rect 4776 2440 4783 2443
rect 4773 2427 4787 2440
rect 4756 2256 4763 2313
rect 4796 2227 4803 2254
rect 4676 1956 4683 1993
rect 4716 1956 4723 1993
rect 4736 1967 4743 2223
rect 4776 2047 4783 2193
rect 4816 2167 4823 2253
rect 4796 1927 4803 1954
rect 4556 1776 4583 1783
rect 4536 1716 4543 1753
rect 4556 1727 4563 1776
rect 4576 1467 4583 1753
rect 4816 1747 4823 1953
rect 4836 1927 4843 2573
rect 4976 2527 4983 2933
rect 4996 2547 5003 2653
rect 5016 2607 5023 2952
rect 4856 1727 4863 2493
rect 4896 2427 4903 2513
rect 5016 2446 5023 2493
rect 4947 2403 4960 2407
rect 4947 2393 4963 2403
rect 4876 2347 4883 2393
rect 4916 2347 4923 2373
rect 4936 2268 4943 2372
rect 4956 2327 4963 2393
rect 4976 2387 4983 2432
rect 5036 2407 5043 3233
rect 5116 3027 5123 3353
rect 5136 3147 5143 3333
rect 5156 3247 5163 3413
rect 5156 3023 5163 3113
rect 5176 3107 5183 3996
rect 5196 3947 5203 4003
rect 5196 3823 5203 3933
rect 5216 3887 5223 3913
rect 5196 3816 5223 3823
rect 5256 3816 5263 3873
rect 5316 3827 5323 4213
rect 5376 4083 5383 4313
rect 5416 4267 5423 4913
rect 5487 4903 5500 4907
rect 5487 4893 5503 4903
rect 5496 4856 5503 4893
rect 5536 4856 5543 4932
rect 5576 4927 5583 5013
rect 5576 4867 5583 4913
rect 5596 4887 5603 5313
rect 5616 5127 5623 5813
rect 5636 5263 5643 5453
rect 5656 5287 5663 5553
rect 5716 5467 5723 5973
rect 5736 5863 5743 5993
rect 5756 5987 5763 7113
rect 5776 6267 5783 7373
rect 5796 7127 5803 7553
rect 5836 7456 5843 7513
rect 5796 6947 5803 7092
rect 5816 7087 5823 7413
rect 5836 6968 5843 7393
rect 5856 7387 5863 7423
rect 5916 7407 5923 7513
rect 5936 7347 5943 8053
rect 5956 7907 5963 8113
rect 5976 7927 5983 8073
rect 5956 7187 5963 7893
rect 5976 7547 5983 7673
rect 5976 7507 5983 7533
rect 5976 7307 5983 7454
rect 5896 7087 5903 7123
rect 5976 7123 5983 7293
rect 5956 7116 5983 7123
rect 5936 7103 5943 7112
rect 5916 7096 5943 7103
rect 5876 6847 5883 7073
rect 5896 6767 5903 6953
rect 5916 6747 5923 7096
rect 5896 6683 5903 6713
rect 5936 6687 5943 6953
rect 5956 6767 5963 7116
rect 5996 7087 6003 8156
rect 6036 8107 6043 8393
rect 6056 8127 6063 8194
rect 6033 7980 6047 7993
rect 6036 7976 6043 7980
rect 6076 7976 6083 8073
rect 6096 8027 6103 8432
rect 6196 8407 6203 8494
rect 6116 7976 6123 8313
rect 6256 8247 6263 8463
rect 6176 8196 6183 8233
rect 6213 8200 6227 8213
rect 6216 8196 6223 8200
rect 6156 8147 6163 8163
rect 6147 8136 6163 8147
rect 6147 8133 6160 8136
rect 6056 7940 6063 7943
rect 6053 7927 6067 7940
rect 6096 7907 6103 7943
rect 6076 7707 6083 7833
rect 6076 7643 6083 7693
rect 6056 7636 6083 7643
rect 6016 7127 6023 7613
rect 6096 7607 6103 7773
rect 6073 7460 6087 7473
rect 6076 7456 6083 7460
rect 6056 7420 6063 7423
rect 6053 7407 6067 7420
rect 6116 7407 6123 7913
rect 6066 7400 6067 7407
rect 6056 7367 6063 7393
rect 6036 7007 6043 7213
rect 6056 7147 6063 7233
rect 6076 7168 6083 7393
rect 6136 7247 6143 7693
rect 6156 7267 6163 8113
rect 6176 8047 6183 8093
rect 6176 7827 6183 8012
rect 6196 7947 6203 8163
rect 6256 8147 6263 8212
rect 6276 8127 6283 8273
rect 6176 7527 6183 7733
rect 6216 7676 6223 7753
rect 6236 7707 6243 8053
rect 6316 8003 6323 8773
rect 6336 8686 6343 8733
rect 6336 8547 6343 8633
rect 6356 8567 6363 9396
rect 6376 9107 6383 9333
rect 6436 9236 6443 9613
rect 6456 9427 6463 10274
rect 6476 10068 6483 10353
rect 6536 10288 6543 10313
rect 6576 10276 6583 10493
rect 6636 10487 6643 10573
rect 6656 10443 6663 10576
rect 6796 10567 6803 10763
rect 6756 10540 6763 10543
rect 6753 10527 6767 10540
rect 6856 10527 6863 11133
rect 6936 11096 6943 11133
rect 6916 11047 6923 11063
rect 7076 11047 7083 11133
rect 7376 11096 7383 11133
rect 7816 11096 7823 11133
rect 6916 10827 6923 11033
rect 7116 11027 7123 11063
rect 7036 10796 7043 10973
rect 7116 10947 7123 11013
rect 7073 10800 7087 10813
rect 7076 10796 7083 10800
rect 6936 10747 6943 10793
rect 7056 10747 7063 10763
rect 6996 10576 7003 10693
rect 7056 10587 7063 10733
rect 6647 10436 6663 10443
rect 6636 10187 6643 10433
rect 6696 10247 6703 10274
rect 6736 10227 6743 10473
rect 6816 10276 6823 10393
rect 6856 10387 6863 10513
rect 6896 10487 6903 10574
rect 7116 10547 7123 10794
rect 6936 10467 6943 10543
rect 6976 10540 6983 10543
rect 6973 10527 6987 10540
rect 6856 10276 6863 10313
rect 6896 10243 6903 10274
rect 6796 10227 6803 10243
rect 6476 9807 6483 10054
rect 6476 9548 6483 9793
rect 6496 9767 6503 10113
rect 6636 10056 6643 10113
rect 6556 9987 6563 10054
rect 6616 9947 6623 10023
rect 6656 10020 6663 10023
rect 6653 10007 6667 10020
rect 6536 9756 6543 9873
rect 6576 9756 6583 9793
rect 6616 9768 6623 9853
rect 6556 9703 6563 9723
rect 6556 9696 6583 9703
rect 6476 9487 6483 9534
rect 6416 9167 6423 9203
rect 6376 8647 6383 8893
rect 6396 8887 6403 9053
rect 6416 8863 6423 9153
rect 6516 9087 6523 9293
rect 6556 9287 6563 9433
rect 6576 9307 6583 9696
rect 6596 9647 6603 9723
rect 6596 9607 6603 9633
rect 6596 9507 6603 9534
rect 6476 8986 6483 9073
rect 6556 9023 6563 9273
rect 6556 9016 6583 9023
rect 6516 8927 6523 8983
rect 6396 8856 6423 8863
rect 6336 8227 6343 8313
rect 6356 8287 6363 8513
rect 6376 8367 6383 8633
rect 6396 8587 6403 8856
rect 6496 8716 6503 8833
rect 6576 8747 6583 9016
rect 6440 8663 6453 8667
rect 6436 8653 6453 8663
rect 6416 8567 6423 8593
rect 6296 7996 6323 8003
rect 6296 7988 6303 7996
rect 6336 7976 6343 8192
rect 6356 8103 6363 8273
rect 6376 8207 6383 8353
rect 6396 8307 6403 8533
rect 6436 8507 6443 8653
rect 6476 8547 6483 8683
rect 6516 8647 6523 8672
rect 6516 8476 6523 8633
rect 6596 8523 6603 9413
rect 6616 9207 6623 9693
rect 6696 9587 6703 9793
rect 6716 9707 6723 10133
rect 6736 9787 6743 10053
rect 6736 9536 6743 9773
rect 6756 9727 6763 10193
rect 6796 9867 6803 10213
rect 6836 10207 6843 10243
rect 6876 10236 6903 10243
rect 6816 9967 6823 10173
rect 6876 10056 6883 10236
rect 6936 10207 6943 10333
rect 6976 10087 6983 10373
rect 7016 10347 7023 10532
rect 7116 10387 7123 10533
rect 7136 10427 7143 10673
rect 7056 10276 7063 10373
rect 7036 10240 7043 10243
rect 7033 10227 7047 10240
rect 6976 10027 6983 10052
rect 6896 10020 6903 10023
rect 6893 10007 6907 10020
rect 7056 10007 7063 10073
rect 7116 10056 7123 10313
rect 7096 10007 7103 10023
rect 7087 9996 7103 10007
rect 7087 9993 7100 9996
rect 6676 9236 6683 9373
rect 6716 9236 6723 9333
rect 6656 9167 6663 9203
rect 6756 9016 6763 9153
rect 6796 9016 6803 9633
rect 6836 9507 6843 9713
rect 6836 9127 6843 9234
rect 6856 9207 6863 9953
rect 6876 9747 6883 9933
rect 7056 9756 7063 9993
rect 6876 9527 6883 9712
rect 6916 9687 6923 9754
rect 6956 9727 6963 9754
rect 6956 9407 6963 9503
rect 6996 9367 7003 9673
rect 7056 9506 7063 9533
rect 6916 9236 6923 9313
rect 7076 9243 7083 9713
rect 7136 9536 7143 9653
rect 7156 9647 7163 11013
rect 7176 10767 7183 10933
rect 7196 10827 7203 11093
rect 7296 11027 7303 11094
rect 7396 11060 7403 11063
rect 7393 11047 7407 11060
rect 7347 10833 7353 10847
rect 7296 10796 7303 10833
rect 7340 10803 7353 10807
rect 7336 10796 7353 10803
rect 7340 10793 7353 10796
rect 7276 10647 7283 10763
rect 7316 10760 7323 10763
rect 7313 10747 7327 10760
rect 7196 10576 7203 10613
rect 7236 10576 7243 10613
rect 7356 10547 7363 10752
rect 7216 10540 7223 10543
rect 7213 10527 7227 10540
rect 7256 10276 7263 10393
rect 7316 10287 7323 10313
rect 7336 10243 7343 10493
rect 7376 10327 7383 10813
rect 7416 10743 7423 10793
rect 7436 10767 7443 10993
rect 7476 10947 7483 11094
rect 7916 11066 7923 11093
rect 7476 10887 7483 10933
rect 7487 10833 7493 10847
rect 7516 10827 7523 11033
rect 7636 11023 7643 11063
rect 7616 11016 7643 11023
rect 7567 10836 7603 10843
rect 7416 10736 7443 10743
rect 7436 10576 7443 10736
rect 7456 10667 7463 10813
rect 7533 10800 7547 10813
rect 7573 10800 7587 10813
rect 7596 10808 7603 10836
rect 7536 10796 7543 10800
rect 7576 10796 7583 10800
rect 7496 10547 7503 10653
rect 7407 10536 7423 10543
rect 7236 10240 7243 10243
rect 7276 10240 7283 10243
rect 7233 10227 7247 10240
rect 7273 10227 7287 10240
rect 7316 10236 7343 10243
rect 7316 10056 7323 10236
rect 7396 10147 7403 10533
rect 7176 9727 7183 10054
rect 7296 10003 7303 10012
rect 7296 9996 7323 10003
rect 7176 9536 7183 9573
rect 7196 9563 7203 9993
rect 7316 9887 7323 9996
rect 7416 9967 7423 10293
rect 7436 10227 7443 10413
rect 7536 10367 7543 10433
rect 7473 10280 7487 10293
rect 7476 10276 7483 10280
rect 7516 10276 7523 10313
rect 7516 10056 7523 10193
rect 7556 10068 7563 10333
rect 7496 10020 7503 10023
rect 7493 10007 7507 10020
rect 7236 9756 7243 9813
rect 7276 9768 7283 9873
rect 7596 9827 7603 10573
rect 7616 10507 7623 11016
rect 7836 10987 7843 11063
rect 7656 10576 7663 10633
rect 7696 10507 7703 10543
rect 7656 10287 7663 10453
rect 7676 10276 7683 10393
rect 7616 10026 7623 10173
rect 7656 10026 7663 10233
rect 7696 10167 7703 10243
rect 7736 10240 7743 10243
rect 7733 10227 7747 10240
rect 7796 10227 7803 10713
rect 7896 10576 7903 10794
rect 7916 10787 7923 10953
rect 7936 10907 7943 11073
rect 7936 10587 7943 10793
rect 7956 10547 7963 11052
rect 7996 10808 8003 11113
rect 8273 11100 8287 11113
rect 8276 11096 8283 11100
rect 8956 11096 8963 11133
rect 9073 11127 9087 11133
rect 8876 11066 8883 11093
rect 8096 11007 8103 11063
rect 8296 10927 8303 11063
rect 8336 11047 8343 11063
rect 8316 11036 8333 11043
rect 8036 10796 8043 10913
rect 8216 10808 8223 10833
rect 8253 10828 8267 10833
rect 8156 10767 8163 10794
rect 8080 10663 8093 10667
rect 8076 10653 8093 10663
rect 7876 10523 7883 10532
rect 7876 10516 7903 10523
rect 7856 10288 7863 10333
rect 7816 10247 7823 10274
rect 7336 9727 7343 9754
rect 7256 9647 7263 9723
rect 7296 9707 7303 9723
rect 7416 9707 7423 9754
rect 7196 9556 7223 9563
rect 7216 9506 7223 9556
rect 7156 9500 7163 9503
rect 7153 9487 7167 9500
rect 7236 9487 7243 9533
rect 7296 9463 7303 9693
rect 7276 9456 7303 9463
rect 7176 9248 7183 9433
rect 7076 9236 7093 9243
rect 7096 9207 7103 9234
rect 6896 9167 6903 9203
rect 6616 8647 6623 9014
rect 6896 8996 6923 9003
rect 6776 8827 6783 8983
rect 6856 8927 6863 8963
rect 6916 8863 6923 8996
rect 6916 8860 6943 8863
rect 6916 8856 6947 8860
rect 6933 8847 6947 8856
rect 7016 8827 7023 8913
rect 6873 8720 6887 8733
rect 6876 8716 6883 8720
rect 6916 8716 6923 8773
rect 6756 8686 6763 8713
rect 6596 8516 6623 8523
rect 6556 8496 6573 8503
rect 6407 8223 6420 8227
rect 6407 8213 6423 8223
rect 6416 8196 6423 8213
rect 6396 8160 6403 8163
rect 6393 8147 6407 8160
rect 6436 8127 6443 8163
rect 6356 8096 6383 8103
rect 6196 7327 6203 7573
rect 6236 7487 6243 7643
rect 6276 7456 6283 7633
rect 6316 7468 6323 7753
rect 6356 7727 6363 7793
rect 6376 7767 6383 8096
rect 6476 8067 6483 8373
rect 6496 8027 6503 8453
rect 6516 8087 6523 8393
rect 6396 7807 6403 7853
rect 6196 7207 6203 7313
rect 6133 7160 6147 7173
rect 6136 7156 6143 7160
rect 6216 7163 6223 7453
rect 6356 7447 6363 7674
rect 6376 7647 6383 7674
rect 6256 7387 6263 7423
rect 6396 7367 6403 7772
rect 6436 7747 6443 7973
rect 6456 7767 6463 7973
rect 6476 7847 6483 7993
rect 6556 7987 6563 8496
rect 6573 8480 6587 8493
rect 6576 8476 6583 8480
rect 6616 8407 6623 8516
rect 6896 8486 6903 8683
rect 6936 8487 6943 8653
rect 6856 8476 6883 8483
rect 6856 8327 6863 8476
rect 6847 8316 6863 8327
rect 6847 8313 6860 8316
rect 6633 8223 6647 8233
rect 6616 8220 6647 8223
rect 6616 8216 6643 8220
rect 6616 8196 6623 8216
rect 6593 8107 6607 8113
rect 6507 7983 6520 7987
rect 6507 7976 6523 7983
rect 6507 7973 6520 7976
rect 6576 7956 6583 8013
rect 6536 7940 6543 7943
rect 6533 7927 6547 7940
rect 6547 7916 6563 7923
rect 6476 7688 6483 7812
rect 6536 7646 6543 7733
rect 6256 7207 6263 7352
rect 6216 7156 6243 7163
rect 6076 7047 6083 7154
rect 6056 6983 6063 7013
rect 6096 6987 6103 7093
rect 6116 7063 6123 7123
rect 6156 7120 6163 7123
rect 6153 7107 6167 7120
rect 6196 7103 6203 7123
rect 6176 7096 6203 7103
rect 6116 7056 6143 7063
rect 6036 6976 6063 6983
rect 5976 6906 5983 6973
rect 6036 6936 6043 6976
rect 5896 6680 5923 6683
rect 5896 6676 5927 6680
rect 5796 6527 5803 6673
rect 5836 6636 5843 6673
rect 5913 6667 5927 6676
rect 5816 6347 5823 6383
rect 5816 6227 5823 6333
rect 5856 6107 5863 6353
rect 5896 6307 5903 6592
rect 5936 6487 5943 6673
rect 5956 6607 5963 6713
rect 5976 6467 5983 6673
rect 5936 6267 5943 6383
rect 5976 6347 5983 6453
rect 5776 6067 5783 6103
rect 5796 5896 5803 6093
rect 5836 5907 5843 6013
rect 5736 5856 5763 5863
rect 5736 5687 5743 5813
rect 5736 5567 5743 5673
rect 5756 5376 5763 5856
rect 5776 5667 5783 5713
rect 5816 5667 5823 5863
rect 5796 5447 5803 5614
rect 5816 5527 5823 5613
rect 5816 5487 5823 5513
rect 5676 5346 5683 5374
rect 5636 5256 5663 5263
rect 5656 5063 5663 5256
rect 5676 5083 5683 5332
rect 5696 5227 5703 5253
rect 5736 5247 5743 5343
rect 5776 5340 5783 5343
rect 5773 5327 5787 5340
rect 5816 5327 5823 5373
rect 5836 5303 5843 5853
rect 5856 5627 5863 6072
rect 5876 5867 5883 6253
rect 6016 6247 6023 6653
rect 6036 6327 6043 6833
rect 6056 6647 6063 6892
rect 6116 6727 6123 6934
rect 6136 6787 6143 7056
rect 6156 6827 6163 6993
rect 6136 6636 6143 6673
rect 6076 6307 6083 6553
rect 6176 6547 6183 7096
rect 6196 6687 6203 7073
rect 6236 6963 6243 7156
rect 6256 6987 6263 7154
rect 6276 7087 6283 7333
rect 6296 7067 6303 7233
rect 6276 6963 6283 7013
rect 6296 6967 6303 6993
rect 6216 6956 6243 6963
rect 6256 6956 6283 6963
rect 6133 6420 6147 6433
rect 6136 6416 6143 6420
rect 6216 6423 6223 6956
rect 6256 6936 6263 6956
rect 6316 6887 6323 7253
rect 6336 7107 6343 7353
rect 6416 7267 6423 7633
rect 6456 7367 6463 7643
rect 6496 7587 6503 7632
rect 6556 7467 6563 7916
rect 6576 7547 6583 7853
rect 6596 7527 6603 7713
rect 6616 7427 6623 8133
rect 6676 8107 6683 8152
rect 6716 8067 6723 8194
rect 6796 8187 6803 8253
rect 6816 8087 6823 8293
rect 6836 8107 6843 8153
rect 6876 8107 6883 8163
rect 6916 8067 6923 8173
rect 6936 8127 6943 8293
rect 6956 8147 6963 8733
rect 6976 8627 6983 8693
rect 6633 7960 6647 7973
rect 6636 7956 6643 7960
rect 6676 7767 6683 7993
rect 6976 7987 6983 8533
rect 6996 8127 7003 8672
rect 7036 8507 7043 8773
rect 7036 8347 7043 8472
rect 7056 8467 7063 8813
rect 7156 8787 7163 8994
rect 7216 8807 7223 9453
rect 7276 9187 7283 9456
rect 7296 9147 7303 9233
rect 7316 9203 7323 9613
rect 7436 9587 7443 9773
rect 7473 9760 7487 9773
rect 7476 9756 7483 9760
rect 7436 9506 7443 9533
rect 7456 9527 7463 9713
rect 7496 9687 7503 9723
rect 7536 9720 7543 9723
rect 7533 9707 7547 9720
rect 7576 9667 7583 9753
rect 7596 9707 7603 9813
rect 7616 9627 7623 9913
rect 7636 9548 7643 9873
rect 7676 9767 7683 10133
rect 7736 10056 7743 10192
rect 7813 10067 7827 10073
rect 7856 10026 7863 10053
rect 7707 9763 7720 9767
rect 7707 9756 7723 9763
rect 7756 9756 7763 9813
rect 7707 9753 7720 9756
rect 7736 9687 7743 9723
rect 7776 9720 7783 9723
rect 7773 9707 7787 9720
rect 7836 9707 7843 9773
rect 7696 9547 7703 9573
rect 7516 9467 7523 9513
rect 7556 9496 7583 9503
rect 7316 9196 7343 9203
rect 7276 8847 7283 9073
rect 7296 8947 7303 8994
rect 7136 8640 7143 8643
rect 7133 8627 7147 8640
rect 7076 8347 7083 8613
rect 7016 8227 7023 8253
rect 7036 8196 7043 8233
rect 6916 7956 6943 7963
rect 6816 7927 6823 7952
rect 6636 7643 6643 7753
rect 6756 7676 6783 7683
rect 6636 7636 6663 7643
rect 6776 7627 6783 7676
rect 6796 7607 6803 7713
rect 6696 7468 6703 7603
rect 6716 7456 6723 7533
rect 6496 7387 6503 7423
rect 6336 6987 6343 7013
rect 6336 6907 6343 6973
rect 6356 6867 6363 7053
rect 6316 6767 6323 6813
rect 6336 6787 6343 6853
rect 6376 6847 6383 7123
rect 6396 6907 6403 7053
rect 6476 6968 6483 7233
rect 6496 7127 6503 7253
rect 6536 7227 6543 7423
rect 6556 7127 6563 7413
rect 6656 7247 6663 7453
rect 6736 7307 6743 7423
rect 6816 7423 6823 7892
rect 6916 7807 6923 7956
rect 6976 7867 6983 7923
rect 6836 7467 6843 7674
rect 6876 7468 6883 7733
rect 6796 7416 6823 7423
rect 6236 6607 6243 6634
rect 6216 6416 6243 6423
rect 5896 5827 5903 6133
rect 5916 5967 5923 6113
rect 5936 6087 5943 6134
rect 5896 5707 5903 5813
rect 5956 5747 5963 6213
rect 5976 6067 5983 6213
rect 6096 6207 6103 6373
rect 5993 6127 6007 6133
rect 6013 6120 6027 6133
rect 6016 6116 6023 6120
rect 6056 6116 6063 6173
rect 6116 6167 6123 6373
rect 6156 6327 6163 6383
rect 6196 6380 6203 6383
rect 6193 6367 6207 6380
rect 6173 6120 6187 6133
rect 6176 6116 6183 6120
rect 6016 5896 6023 5953
rect 6036 5927 6043 6083
rect 6076 5947 6083 6083
rect 6216 5947 6223 6333
rect 6236 6047 6243 6416
rect 6256 6327 6263 6753
rect 6356 6667 6363 6733
rect 6353 6640 6367 6653
rect 6356 6636 6363 6640
rect 6316 6547 6323 6573
rect 6276 6367 6283 6413
rect 6316 6347 6323 6533
rect 6336 6367 6343 6603
rect 6376 6600 6383 6603
rect 6373 6587 6387 6600
rect 6416 6527 6423 6953
rect 6516 6936 6563 6943
rect 6447 6903 6460 6907
rect 6447 6896 6463 6903
rect 6447 6893 6460 6896
rect 6556 6883 6563 6936
rect 6576 6906 6583 7213
rect 6613 7160 6627 7173
rect 6616 7156 6623 7160
rect 6596 6887 6603 7113
rect 6636 7027 6643 7123
rect 6616 6906 6623 6933
rect 6556 6876 6583 6883
rect 6436 6587 6443 6872
rect 6436 6416 6443 6453
rect 6456 6447 6463 6853
rect 6476 6707 6483 6833
rect 6476 6607 6483 6693
rect 6576 6667 6583 6876
rect 6596 6747 6603 6873
rect 6616 6747 6623 6773
rect 6416 6380 6423 6383
rect 6413 6367 6427 6380
rect 6296 6007 6303 6083
rect 6033 5907 6047 5913
rect 5893 5600 5907 5613
rect 5896 5596 5903 5600
rect 5816 5296 5843 5303
rect 5676 5076 5703 5083
rect 5636 5060 5663 5063
rect 5636 5056 5667 5060
rect 5616 4863 5623 5053
rect 5653 5047 5667 5056
rect 5596 4856 5623 4863
rect 5596 4848 5603 4856
rect 5676 4843 5683 4913
rect 5656 4836 5683 4843
rect 5436 4207 5443 4573
rect 5456 4527 5463 4812
rect 5516 4803 5523 4823
rect 5496 4796 5523 4803
rect 5496 4527 5503 4796
rect 5516 4407 5523 4673
rect 5556 4556 5563 4613
rect 5576 4587 5583 4653
rect 5636 4427 5643 4554
rect 5696 4527 5703 5076
rect 5756 4947 5763 5213
rect 5796 5027 5803 5113
rect 5816 5087 5823 5296
rect 5856 5247 5863 5413
rect 5876 5307 5883 5563
rect 5976 5487 5983 5653
rect 5996 5608 6003 5863
rect 6056 5807 6063 5894
rect 6076 5647 6083 5933
rect 6096 5687 6103 5893
rect 6116 5667 6123 5933
rect 6136 5643 6143 5913
rect 6213 5900 6227 5912
rect 6256 5907 6263 5953
rect 6216 5896 6223 5900
rect 6276 5866 6283 5933
rect 6196 5827 6203 5863
rect 6136 5636 6163 5643
rect 6016 5567 6023 5613
rect 5916 5267 5923 5433
rect 6036 5346 6043 5633
rect 6113 5600 6127 5613
rect 6116 5596 6123 5600
rect 6156 5596 6163 5636
rect 6056 5327 6063 5473
rect 6096 5346 6103 5513
rect 6116 5387 6123 5433
rect 5856 5127 5863 5233
rect 5827 5043 5840 5047
rect 5827 5036 5843 5043
rect 5827 5033 5840 5036
rect 5916 4947 5923 5253
rect 5936 5046 5943 5073
rect 5936 4846 5943 4873
rect 5956 4836 5963 5193
rect 5976 4907 5983 5293
rect 6116 5287 6123 5373
rect 5996 5067 6003 5133
rect 6053 5080 6067 5093
rect 6056 5076 6063 5080
rect 6036 5023 6043 5032
rect 6036 5016 6063 5023
rect 5716 4527 5723 4573
rect 5816 4556 5823 4693
rect 5856 4567 5863 4713
rect 5456 4327 5463 4373
rect 5596 4306 5603 4393
rect 5736 4387 5743 4554
rect 5756 4336 5763 4513
rect 5836 4407 5843 4523
rect 5656 4306 5663 4333
rect 5816 4307 5823 4334
rect 5356 4076 5383 4083
rect 5336 3786 5343 4033
rect 5196 3308 5203 3773
rect 5276 3447 5283 3783
rect 5356 3543 5363 4076
rect 5456 4048 5463 4273
rect 5556 4107 5563 4173
rect 5496 4036 5503 4093
rect 5436 3967 5443 4003
rect 5476 4000 5483 4003
rect 5473 3987 5487 4000
rect 5516 3816 5523 3853
rect 5396 3647 5403 3814
rect 5456 3667 5463 3783
rect 5476 3707 5483 3753
rect 5496 3727 5503 3783
rect 5556 3747 5563 4093
rect 5356 3536 5383 3543
rect 5336 3516 5363 3523
rect 5236 3296 5243 3393
rect 5276 3296 5283 3333
rect 5156 3016 5183 3023
rect 5176 3008 5183 3016
rect 5056 2927 5063 2994
rect 5036 2307 5043 2393
rect 4936 1956 4943 2053
rect 4956 2007 4963 2223
rect 4996 2127 5003 2193
rect 5016 2127 5023 2254
rect 5016 2087 5023 2113
rect 4876 1747 4883 1913
rect 4916 1887 4923 1923
rect 4716 1687 4723 1723
rect 4816 1716 4843 1723
rect 4736 1663 4743 1713
rect 4716 1656 4743 1663
rect 4596 1436 4603 1493
rect 4616 1467 4623 1533
rect 4536 1223 4543 1293
rect 4527 1216 4543 1223
rect 4496 947 4503 1183
rect 4556 1167 4563 1213
rect 4556 1067 4563 1113
rect 4576 1027 4583 1403
rect 4596 1087 4603 1333
rect 4376 696 4383 733
rect 4356 660 4363 663
rect 4353 647 4367 660
rect 4427 633 4433 647
rect 4336 607 4343 633
rect 4176 247 4183 333
rect 3296 136 3323 143
rect 2847 116 2863 127
rect 2847 113 2860 116
rect 3556 67 3563 173
rect 3796 107 3803 174
rect 4236 146 4243 433
rect 4356 396 4363 473
rect 4316 307 4323 393
rect 4456 366 4463 413
rect 4496 403 4503 773
rect 4596 727 4603 933
rect 4616 927 4623 1273
rect 4656 1087 4663 1573
rect 4696 1527 4703 1613
rect 4716 1448 4723 1656
rect 4816 1567 4823 1716
rect 4836 1587 4843 1653
rect 4876 1627 4883 1683
rect 4816 1566 4840 1567
rect 4816 1556 4833 1566
rect 4820 1553 4833 1556
rect 4736 1267 4743 1453
rect 4776 1436 4783 1533
rect 4796 1467 4803 1553
rect 4827 1493 4833 1507
rect 4796 1287 4803 1403
rect 4856 1327 4863 1573
rect 4876 1487 4883 1613
rect 4716 1240 4763 1243
rect 4716 1236 4767 1240
rect 4716 1216 4723 1236
rect 4753 1227 4767 1236
rect 4776 1186 4783 1253
rect 4696 1027 4703 1172
rect 4796 1167 4803 1213
rect 4647 943 4660 947
rect 4647 933 4663 943
rect 4656 916 4663 933
rect 4716 827 4723 1073
rect 4616 696 4623 813
rect 4516 627 4523 694
rect 4656 666 4663 713
rect 4556 547 4563 663
rect 4496 396 4523 403
rect 4616 396 4623 613
rect 4736 427 4743 893
rect 4756 886 4763 1133
rect 4816 1127 4823 1313
rect 4896 1287 4903 1673
rect 4916 1487 4923 1833
rect 4936 1767 4943 1853
rect 4936 1587 4943 1732
rect 4933 1507 4947 1513
rect 4956 1463 4963 1923
rect 4996 1823 5003 1953
rect 4976 1816 5003 1823
rect 4976 1567 4983 1816
rect 4996 1587 5003 1793
rect 5016 1507 5023 1713
rect 5036 1468 5043 2272
rect 5056 1847 5063 2673
rect 5076 2227 5083 2913
rect 5156 2807 5163 2963
rect 5113 2780 5127 2793
rect 5116 2776 5123 2780
rect 5096 2427 5103 2473
rect 5116 2327 5123 2713
rect 5156 2607 5163 2743
rect 5176 2523 5183 2773
rect 5196 2567 5203 2873
rect 5216 2788 5223 2953
rect 5236 2647 5243 2993
rect 5256 2967 5263 3263
rect 5256 2727 5263 2932
rect 5276 2707 5283 3233
rect 5296 3087 5303 3173
rect 5296 2867 5303 2893
rect 5316 2887 5323 3433
rect 5176 2516 5203 2523
rect 5173 2480 5187 2493
rect 5196 2487 5203 2516
rect 5176 2476 5183 2480
rect 5216 2387 5223 2533
rect 5076 1736 5083 1773
rect 5096 1767 5103 2293
rect 5173 2260 5187 2273
rect 5176 2256 5183 2260
rect 5216 2256 5223 2373
rect 5236 2267 5243 2593
rect 5156 2187 5163 2223
rect 5156 1968 5163 2093
rect 5176 1967 5183 2153
rect 5216 2143 5223 2193
rect 5196 2136 5223 2143
rect 5196 2067 5203 2136
rect 5236 1923 5243 2113
rect 5256 2107 5263 2513
rect 5276 2287 5283 2633
rect 5276 2187 5283 2252
rect 5296 2127 5303 2793
rect 5316 2783 5323 2833
rect 5336 2807 5343 3313
rect 5356 3007 5363 3516
rect 5376 3387 5383 3536
rect 5376 3187 5383 3373
rect 5376 2996 5383 3152
rect 5396 3027 5403 3633
rect 5416 3347 5423 3633
rect 5436 3303 5443 3553
rect 5456 3327 5463 3653
rect 5513 3520 5527 3533
rect 5516 3516 5523 3520
rect 5556 3516 5563 3693
rect 5576 3527 5583 4193
rect 5596 3308 5603 4153
rect 5700 4063 5713 4067
rect 5696 4053 5713 4063
rect 5696 4036 5703 4053
rect 5756 4007 5763 4253
rect 5416 3296 5463 3303
rect 5416 3027 5423 3296
rect 5476 3260 5483 3263
rect 5473 3247 5487 3260
rect 5476 3087 5483 3233
rect 5556 3187 5563 3293
rect 5616 3127 5623 3893
rect 5676 3867 5683 4003
rect 5716 4000 5723 4003
rect 5713 3987 5727 4000
rect 5776 3887 5783 4303
rect 5796 3907 5803 4233
rect 5693 3820 5707 3833
rect 5696 3816 5703 3820
rect 5756 3747 5763 3783
rect 5636 3267 5643 3533
rect 5656 3367 5663 3513
rect 5436 3003 5443 3033
rect 5416 2996 5443 3003
rect 5396 2927 5403 2963
rect 5356 2807 5363 2893
rect 5316 2776 5343 2783
rect 5376 2776 5383 2893
rect 5456 2803 5463 3013
rect 5596 2996 5603 3073
rect 5636 2996 5643 3253
rect 5656 3227 5663 3353
rect 5556 2960 5573 2963
rect 5553 2956 5573 2960
rect 5553 2947 5567 2956
rect 5436 2796 5463 2803
rect 5396 2707 5403 2743
rect 5316 2207 5323 2473
rect 5436 2387 5443 2796
rect 5456 2746 5463 2773
rect 5336 2307 5343 2373
rect 5336 2087 5343 2272
rect 5376 2263 5383 2373
rect 5516 2307 5523 2893
rect 5616 2887 5623 2963
rect 5356 2256 5383 2263
rect 5356 2167 5363 2256
rect 5416 2187 5423 2223
rect 5456 2220 5463 2223
rect 5453 2207 5467 2220
rect 5496 2127 5503 2253
rect 5516 2207 5523 2293
rect 5536 2187 5543 2873
rect 5613 2780 5627 2793
rect 5616 2776 5623 2780
rect 5596 2687 5603 2743
rect 5576 2547 5583 2653
rect 5676 2547 5683 3573
rect 5696 3447 5703 3693
rect 5776 3516 5783 3653
rect 5796 3547 5803 3814
rect 5816 3587 5823 4293
rect 5836 3787 5843 4173
rect 5856 4107 5863 4313
rect 5916 4207 5923 4693
rect 5936 4507 5943 4793
rect 5996 4767 6003 4803
rect 6036 4767 6043 4933
rect 6056 4707 6063 5016
rect 6113 4987 6127 4993
rect 6136 4927 6143 5563
rect 6176 5527 6183 5563
rect 6216 5387 6223 5653
rect 6236 5343 6243 5831
rect 6256 5427 6263 5733
rect 6316 5547 6323 6033
rect 6336 5847 6343 6313
rect 6336 5687 6343 5733
rect 6356 5667 6363 6193
rect 6376 6087 6383 6333
rect 6396 6007 6403 6153
rect 6416 5967 6423 6233
rect 6476 6207 6483 6572
rect 6496 6347 6503 6634
rect 6516 6127 6523 6653
rect 6576 6636 6583 6653
rect 6536 6167 6543 6372
rect 6556 6167 6563 6513
rect 6376 5687 6383 5893
rect 6416 5827 6423 5863
rect 6416 5627 6423 5813
rect 6496 5787 6503 6072
rect 6467 5753 6473 5767
rect 6373 5600 6387 5613
rect 6436 5603 6443 5673
rect 6376 5596 6383 5600
rect 6416 5596 6443 5603
rect 6193 5327 6207 5332
rect 6216 5336 6243 5343
rect 6156 4987 6163 5313
rect 6156 4903 6163 4952
rect 6136 4896 6163 4903
rect 5956 4567 5963 4593
rect 6016 4556 6023 4613
rect 6076 4588 6083 4853
rect 6116 4687 6123 4893
rect 6116 4627 6123 4673
rect 5993 4547 6007 4553
rect 5976 4336 5983 4393
rect 6036 4367 6043 4523
rect 5956 4127 5963 4303
rect 5996 4227 6003 4303
rect 6076 4267 6083 4493
rect 6136 4287 6143 4896
rect 6176 4867 6183 5253
rect 6196 4903 6203 5273
rect 6216 4967 6223 5336
rect 6256 5076 6263 5392
rect 6293 5080 6307 5093
rect 6316 5087 6323 5373
rect 6336 5267 6343 5513
rect 6356 5387 6363 5433
rect 6396 5408 6403 5563
rect 6456 5447 6463 5593
rect 6476 5566 6483 5653
rect 6476 5346 6483 5373
rect 6296 5076 6303 5080
rect 6233 4967 6247 4973
rect 6196 4900 6223 4903
rect 6196 4896 6227 4900
rect 6213 4887 6227 4896
rect 6193 4860 6207 4873
rect 6196 4856 6203 4860
rect 6236 4856 6243 4913
rect 6156 4307 6163 4833
rect 6216 4820 6223 4823
rect 6213 4807 6227 4820
rect 6316 4807 6323 4873
rect 6176 4427 6183 4673
rect 6196 4336 6203 4573
rect 6276 4556 6283 4793
rect 6316 4667 6323 4793
rect 6336 4607 6343 5193
rect 6256 4520 6263 4523
rect 6253 4507 6267 4520
rect 6216 4287 6223 4303
rect 6207 4276 6223 4287
rect 6207 4273 6220 4276
rect 6136 4247 6143 4273
rect 5856 3907 5863 4033
rect 5856 3543 5863 3872
rect 5876 3567 5883 4073
rect 5896 4068 5903 4093
rect 5956 4036 5983 4043
rect 5896 3707 5903 3893
rect 5976 3867 5983 4036
rect 5916 3647 5923 3693
rect 5976 3647 5983 3783
rect 6016 3667 6023 4113
rect 6036 3828 6043 4073
rect 6076 3807 6083 3893
rect 6096 3828 6103 4193
rect 6176 4047 6183 4253
rect 6216 4087 6223 4253
rect 6216 4036 6243 4043
rect 6116 3927 6123 4033
rect 6136 3967 6143 4003
rect 6236 3827 6243 4036
rect 6156 3780 6163 3783
rect 6153 3767 6167 3780
rect 6276 3747 6283 3913
rect 5856 3536 5883 3543
rect 5756 3407 5763 3483
rect 5747 3296 5763 3303
rect 5696 2746 5703 2813
rect 5576 2227 5583 2443
rect 5696 2327 5703 2474
rect 5656 2256 5663 2293
rect 5696 2256 5703 2313
rect 5716 2287 5723 3113
rect 5756 3063 5763 3296
rect 5796 3267 5803 3483
rect 5836 3447 5843 3503
rect 5756 3056 5783 3063
rect 5776 2947 5783 3056
rect 5856 3023 5863 3373
rect 5876 3147 5883 3536
rect 5936 3503 5943 3613
rect 6236 3587 6243 3633
rect 6236 3536 6243 3573
rect 5896 3496 5943 3503
rect 5896 3407 5903 3473
rect 6176 3403 6183 3433
rect 6156 3396 6183 3403
rect 5916 3296 5923 3373
rect 6156 3296 6163 3396
rect 5936 3227 5943 3263
rect 5856 3016 5883 3023
rect 5876 2996 5883 3016
rect 5916 2967 5923 3033
rect 5756 2607 5763 2774
rect 5816 2740 5823 2743
rect 5813 2727 5827 2740
rect 5807 2696 5833 2703
rect 5776 2307 5783 2443
rect 5756 2227 5763 2293
rect 5636 2220 5643 2223
rect 5633 2207 5647 2220
rect 5676 2203 5683 2223
rect 5716 2220 5723 2223
rect 5713 2207 5727 2220
rect 5676 2196 5703 2203
rect 5496 2087 5503 2113
rect 5276 1987 5283 2073
rect 5136 1887 5143 1923
rect 5216 1916 5243 1923
rect 5216 1887 5223 1916
rect 5056 1627 5063 1653
rect 4956 1456 5003 1463
rect 4996 1436 5003 1456
rect 4836 947 4843 1033
rect 4856 1007 4863 1273
rect 4913 1220 4927 1233
rect 4916 1216 4923 1220
rect 4876 1186 4883 1213
rect 4936 1067 4943 1183
rect 4896 967 4903 993
rect 4896 916 4903 953
rect 4816 847 4823 914
rect 4816 787 4823 833
rect 4813 700 4827 713
rect 4816 696 4823 700
rect 4796 660 4803 663
rect 4856 660 4863 663
rect 4793 647 4807 660
rect 4853 647 4867 660
rect 4836 396 4843 433
rect 4876 403 4883 883
rect 4976 743 4983 1403
rect 4996 1247 5003 1293
rect 5016 1267 5023 1403
rect 4956 736 4983 743
rect 4876 396 4903 403
rect 4156 140 4163 143
rect 4153 127 4167 140
rect 4256 87 4263 173
rect 4296 127 4303 173
rect 4316 146 4323 293
rect 4416 267 4423 363
rect 4476 67 4483 174
rect 4496 147 4503 373
rect 4516 366 4523 396
rect 4896 366 4903 396
rect 4936 366 4943 693
rect 4956 647 4963 736
rect 5056 727 5063 1373
rect 5076 1367 5083 1433
rect 5096 1387 5103 1453
rect 5116 1367 5123 1393
rect 5136 1387 5143 1593
rect 5076 1327 5083 1353
rect 5156 1243 5163 1753
rect 5176 1527 5183 1734
rect 5196 1707 5203 1833
rect 5216 1727 5223 1873
rect 5256 1867 5263 1943
rect 5276 1767 5283 1933
rect 5296 1907 5303 2033
rect 5436 1936 5443 2033
rect 5236 1507 5243 1753
rect 5296 1736 5303 1773
rect 5333 1740 5347 1753
rect 5336 1736 5343 1740
rect 5376 1706 5383 1833
rect 5536 1767 5543 2133
rect 5596 1976 5603 2013
rect 5636 1967 5643 2073
rect 5276 1647 5283 1703
rect 5396 1567 5403 1673
rect 5496 1627 5503 1713
rect 5576 1703 5583 1753
rect 5556 1696 5583 1703
rect 5233 1440 5247 1453
rect 5236 1436 5243 1440
rect 5216 1383 5223 1403
rect 5216 1376 5243 1383
rect 5136 1236 5163 1243
rect 5136 1216 5143 1236
rect 5176 1216 5183 1273
rect 5076 1127 5083 1193
rect 5236 1183 5243 1376
rect 5256 1247 5263 1403
rect 5116 1027 5123 1183
rect 5116 947 5123 1013
rect 5156 947 5163 1183
rect 5196 1127 5203 1183
rect 5216 1176 5243 1183
rect 5156 923 5163 933
rect 5136 916 5163 923
rect 4976 666 4983 713
rect 4993 707 5007 713
rect 5016 660 5023 663
rect 5013 647 5027 660
rect 4636 327 4643 352
rect 4816 287 4823 313
rect 4856 287 4863 363
rect 5036 327 5043 363
rect 4653 180 4667 193
rect 4896 188 4903 253
rect 4953 188 4967 193
rect 5096 188 5103 333
rect 4656 176 4663 180
rect 5136 146 5143 413
rect 5156 188 5163 793
rect 5176 267 5183 993
rect 5216 696 5223 1176
rect 5296 923 5303 1493
rect 5376 1406 5383 1473
rect 5336 1207 5343 1293
rect 5396 1216 5403 1473
rect 5476 1307 5483 1403
rect 5476 1186 5483 1233
rect 5536 1228 5543 1433
rect 5556 1347 5563 1493
rect 5276 916 5303 923
rect 5336 916 5343 1033
rect 5373 920 5387 933
rect 5376 916 5383 920
rect 5276 727 5283 916
rect 5316 807 5323 883
rect 5236 607 5243 663
rect 5256 396 5263 433
rect 5196 366 5203 393
rect 5236 287 5243 363
rect 5276 176 5323 183
rect 5316 147 5323 176
rect 4636 107 4643 143
rect 5176 67 5183 143
rect 5236 140 5243 143
rect 5233 127 5247 140
rect 5336 -24 5343 713
rect 5356 607 5363 872
rect 5496 767 5503 1213
rect 5516 1167 5523 1193
rect 5516 886 5523 973
rect 5556 916 5563 1333
rect 5596 1223 5603 1773
rect 5616 1407 5623 1933
rect 5636 1847 5643 1873
rect 5656 1667 5663 2013
rect 5676 1547 5683 2173
rect 5696 1687 5703 2196
rect 5716 1867 5723 2053
rect 5736 1947 5743 2033
rect 5756 1887 5763 2033
rect 5776 2007 5783 2272
rect 5796 2207 5803 2293
rect 5796 1968 5803 2193
rect 5816 2147 5823 2254
rect 5836 1956 5843 2353
rect 5856 2307 5863 2913
rect 5856 2207 5863 2293
rect 5896 2268 5903 2474
rect 5936 2387 5943 3013
rect 5976 2927 5983 3263
rect 6076 2996 6083 3293
rect 6276 3287 6283 3573
rect 6296 3276 6303 3493
rect 6316 3447 6323 4393
rect 6336 4306 6343 4433
rect 6356 4407 6363 5293
rect 6376 5167 6383 5343
rect 6416 5340 6423 5343
rect 6413 5327 6427 5340
rect 6496 5307 6503 5752
rect 6376 4647 6383 5153
rect 6396 4767 6403 5133
rect 6416 4947 6423 5093
rect 6456 5083 6463 5233
rect 6476 5147 6483 5253
rect 6436 5076 6463 5083
rect 6476 5076 6483 5112
rect 6516 5107 6523 6073
rect 6536 6067 6543 6153
rect 6556 6087 6563 6113
rect 6536 5527 6543 5953
rect 6556 5866 6563 5973
rect 6576 5767 6583 6553
rect 6636 6507 6643 6953
rect 6656 6787 6663 7093
rect 6656 6607 6663 6752
rect 6616 6428 6623 6453
rect 6656 6416 6663 6572
rect 6676 6567 6683 7113
rect 6716 7103 6723 7253
rect 6756 7107 6763 7313
rect 6776 7126 6783 7193
rect 6796 7127 6803 7416
rect 6836 7407 6843 7453
rect 6816 7347 6823 7373
rect 6896 7267 6903 7693
rect 6936 7676 6943 7733
rect 7016 7587 7023 8073
rect 7036 7947 7043 8033
rect 7036 7647 7043 7674
rect 6916 7426 6923 7533
rect 6976 7420 6983 7423
rect 6973 7407 6987 7420
rect 7056 7423 7063 8131
rect 7076 7707 7083 8153
rect 7096 7787 7103 8593
rect 7176 8536 7183 8573
rect 7236 8466 7243 8613
rect 7136 8327 7143 8373
rect 7126 8233 7127 8240
rect 7113 8227 7127 8233
rect 7116 8027 7123 8152
rect 7136 8107 7143 8233
rect 7176 8007 7183 8213
rect 7196 8167 7203 8393
rect 7256 8227 7263 8813
rect 7296 8727 7303 8933
rect 7276 8508 7283 8553
rect 7296 8307 7303 8513
rect 7316 8407 7323 9173
rect 7233 8200 7247 8213
rect 7236 8196 7243 8200
rect 7256 8087 7263 8163
rect 7173 7980 7187 7993
rect 7176 7976 7183 7980
rect 7116 7727 7123 7773
rect 7196 7707 7203 7943
rect 7256 7867 7263 8033
rect 7200 7643 7213 7647
rect 7156 7583 7163 7643
rect 7196 7636 7213 7643
rect 7200 7633 7213 7636
rect 7236 7627 7243 7674
rect 7256 7647 7263 7693
rect 7276 7647 7283 8093
rect 7296 7803 7303 8163
rect 7316 7827 7323 8153
rect 7336 7907 7343 9196
rect 7356 8767 7363 9093
rect 7376 9067 7383 9203
rect 7416 9147 7423 9203
rect 7376 8747 7383 9014
rect 7396 8728 7403 9073
rect 7456 9028 7463 9333
rect 7496 9027 7503 9293
rect 7516 8963 7523 9453
rect 7536 9087 7543 9492
rect 7556 9206 7563 9496
rect 7556 8987 7563 9192
rect 7507 8956 7523 8963
rect 7376 8607 7383 8683
rect 7436 8667 7443 8873
rect 7456 8687 7463 8853
rect 7496 8607 7503 8953
rect 7516 8767 7523 8913
rect 7576 8723 7583 9173
rect 7596 8947 7603 9203
rect 7676 9187 7683 9534
rect 7776 9243 7783 9593
rect 7876 9536 7883 10373
rect 7896 10327 7903 10516
rect 7896 9863 7903 10313
rect 7916 10287 7923 10543
rect 8036 10546 8043 10633
rect 8076 10627 8083 10653
rect 8093 10580 8107 10593
rect 8096 10576 8103 10580
rect 8136 10576 8143 10713
rect 8176 10587 8183 10653
rect 8196 10647 8203 10763
rect 8296 10763 8303 10913
rect 8316 10767 8323 11036
rect 8536 11027 8543 11063
rect 8716 11060 8723 11063
rect 8713 11047 8727 11060
rect 8756 10967 8763 11063
rect 8976 11027 8983 11063
rect 9036 10967 9043 11094
rect 8276 10756 8303 10763
rect 8156 10387 8163 10543
rect 7980 10283 7993 10287
rect 7976 10276 7993 10283
rect 7980 10273 7993 10276
rect 8116 10147 8123 10313
rect 8147 10283 8160 10287
rect 8147 10276 8163 10283
rect 8216 10276 8223 10493
rect 8276 10327 8283 10756
rect 8336 10727 8343 10793
rect 8313 10580 8327 10593
rect 8316 10576 8323 10580
rect 8356 10576 8363 10813
rect 8396 10766 8403 10873
rect 8456 10827 8463 10853
rect 8453 10800 8467 10813
rect 8493 10800 8507 10813
rect 8516 10808 8523 10853
rect 8456 10796 8463 10800
rect 8496 10796 8503 10800
rect 8436 10546 8443 10752
rect 8476 10647 8483 10763
rect 8553 10588 8567 10593
rect 8596 10576 8603 10833
rect 8736 10796 8743 10833
rect 8976 10796 9023 10803
rect 8656 10687 8663 10752
rect 8676 10707 8683 10763
rect 8376 10387 8383 10543
rect 8576 10540 8583 10543
rect 8616 10540 8623 10543
rect 8573 10527 8587 10540
rect 8613 10527 8627 10540
rect 8616 10387 8623 10513
rect 8656 10487 8663 10673
rect 8676 10527 8683 10693
rect 8716 10667 8723 10763
rect 9016 10727 9023 10796
rect 8836 10576 8843 10713
rect 9036 10607 9043 10793
rect 9076 10767 9083 10993
rect 8736 10507 8743 10553
rect 8756 10467 8763 10574
rect 8896 10546 8903 10573
rect 8773 10527 8787 10533
rect 8816 10487 8823 10543
rect 8413 10280 8427 10293
rect 8416 10276 8423 10280
rect 8456 10276 8463 10313
rect 8147 10273 8160 10276
rect 8136 10187 8143 10273
rect 8176 10207 8183 10243
rect 8396 10240 8403 10243
rect 8393 10227 8407 10240
rect 8376 10216 8393 10223
rect 8176 10167 8183 10193
rect 8196 10056 8203 10213
rect 7936 9987 7943 10053
rect 8296 10026 8303 10133
rect 8316 10127 8323 10153
rect 7896 9856 7913 9863
rect 7816 9427 7823 9503
rect 7916 9407 7923 9853
rect 7936 9763 7943 9973
rect 7976 9867 7983 10023
rect 7936 9756 7963 9763
rect 7996 9756 8003 9933
rect 8016 9927 8023 10023
rect 8256 9987 8263 10023
rect 8016 9887 8023 9913
rect 7916 9287 7923 9393
rect 7776 9236 7803 9243
rect 7836 9236 7843 9273
rect 7896 9203 7903 9253
rect 8016 9243 8023 9723
rect 8056 9607 8063 9754
rect 8156 9667 8163 9754
rect 8296 9726 8303 10012
rect 8316 10007 8323 10053
rect 8356 9987 8363 10054
rect 8376 10026 8383 10216
rect 8436 10207 8443 10243
rect 8496 10207 8503 10274
rect 8536 10207 8543 10293
rect 8596 10246 8603 10313
rect 8693 10280 8707 10293
rect 8696 10276 8703 10280
rect 8576 10236 8593 10243
rect 8476 10056 8483 10113
rect 8376 9947 8383 10012
rect 8436 9967 8443 9993
rect 8496 9967 8503 10023
rect 8456 9756 8463 9793
rect 8056 9536 8063 9593
rect 8116 9567 8123 9633
rect 8216 9527 8223 9723
rect 8476 9667 8483 9723
rect 8516 9723 8523 9754
rect 8507 9716 8523 9723
rect 8496 9647 8503 9712
rect 8076 9327 8083 9503
rect 8256 9467 8263 9573
rect 8313 9540 8327 9553
rect 8316 9536 8323 9540
rect 8296 9427 8303 9503
rect 8436 9467 8443 9513
rect 8456 9506 8463 9553
rect 8496 9536 8503 9633
rect 8536 9536 8543 9573
rect 8576 9543 8583 10236
rect 8676 10207 8683 10243
rect 8716 10127 8723 10232
rect 8736 10207 8743 10453
rect 8716 10056 8723 10113
rect 8576 9536 8603 9543
rect 8596 9506 8603 9536
rect 7996 9236 8023 9243
rect 7956 9207 7963 9234
rect 7876 9196 7903 9203
rect 7653 9020 7667 9033
rect 7656 9016 7663 9020
rect 7716 8983 7723 9013
rect 7816 8986 7823 9033
rect 7876 9016 7883 9196
rect 7636 8980 7643 8983
rect 7633 8967 7647 8980
rect 7676 8976 7723 8983
rect 7856 8927 7863 8983
rect 7556 8716 7583 8723
rect 7636 8716 7643 8913
rect 7536 8686 7543 8713
rect 7356 8147 7363 8573
rect 7453 8540 7467 8553
rect 7456 8536 7463 8540
rect 7496 8496 7523 8503
rect 7516 8467 7523 8496
rect 7376 8456 7403 8463
rect 7376 8367 7383 8456
rect 7356 8087 7363 8112
rect 7376 8087 7383 8353
rect 7396 8107 7403 8393
rect 7416 8127 7423 8253
rect 7436 8187 7443 8313
rect 7496 8196 7503 8293
rect 7516 8247 7523 8432
rect 7536 8327 7543 8533
rect 7556 8407 7563 8716
rect 7676 8683 7683 8893
rect 7656 8676 7683 8683
rect 7656 8663 7663 8676
rect 7636 8656 7663 8663
rect 7576 8367 7583 8653
rect 7596 8267 7603 8573
rect 7616 8447 7623 8613
rect 7636 8387 7643 8656
rect 7696 8496 7703 8714
rect 7716 8687 7723 8773
rect 7736 8507 7743 8593
rect 7776 8507 7783 8833
rect 7876 8716 7883 8773
rect 7976 8707 7983 9053
rect 7996 8787 8003 9236
rect 8073 9240 8087 9253
rect 8076 9236 8083 9240
rect 8056 9200 8063 9203
rect 8053 9187 8067 9200
rect 8116 9187 8123 9313
rect 8196 9248 8203 9353
rect 8276 9236 8283 9333
rect 8416 9248 8423 9273
rect 8456 9236 8463 9333
rect 8016 8986 8023 9133
rect 8096 9016 8103 9093
rect 8156 8986 8163 9033
rect 8196 8907 8203 9234
rect 8256 9027 8263 9203
rect 8316 9016 8323 9053
rect 8416 8947 8423 9234
rect 8476 9187 8483 9203
rect 8476 9176 8493 9187
rect 8480 9173 8493 9176
rect 7996 8700 8003 8703
rect 7816 8483 7823 8673
rect 7856 8486 7863 8683
rect 7896 8607 7903 8683
rect 7936 8587 7943 8692
rect 7993 8687 8007 8700
rect 8036 8627 8043 8833
rect 8176 8696 8183 8733
rect 7796 8476 7823 8483
rect 7676 8427 7683 8452
rect 7796 8327 7803 8476
rect 8096 8476 8123 8483
rect 7596 8163 7603 8214
rect 7476 8127 7483 8163
rect 7576 8156 7603 8163
rect 7376 8086 7400 8087
rect 7376 8076 7393 8086
rect 7380 8073 7393 8076
rect 7376 7976 7383 8053
rect 7456 7947 7463 7973
rect 7296 7796 7323 7803
rect 7136 7576 7163 7583
rect 7036 7416 7063 7423
rect 6893 7160 6907 7173
rect 6896 7156 6903 7160
rect 6696 7096 6723 7103
rect 6696 6967 6703 7096
rect 6876 7007 6883 7123
rect 6753 6980 6767 6993
rect 6756 6976 6763 6980
rect 6836 6906 6843 6993
rect 6896 6948 6903 7013
rect 6916 6847 6923 7112
rect 6936 7087 6943 7173
rect 7016 7167 7023 7213
rect 6956 7087 6963 7154
rect 7036 7067 7043 7416
rect 7096 7387 7103 7573
rect 7116 7247 7123 7513
rect 7136 7327 7143 7576
rect 7156 7287 7163 7553
rect 7196 7456 7203 7613
rect 7236 7456 7243 7533
rect 7276 7507 7283 7612
rect 7216 7307 7223 7423
rect 7167 7276 7183 7283
rect 6936 6847 6943 6933
rect 6696 6587 6703 6613
rect 6716 6567 6723 6773
rect 7016 6747 7023 6892
rect 7056 6727 7063 6753
rect 7036 6667 7043 6693
rect 6756 6567 6763 6603
rect 6796 6527 6803 6603
rect 6676 6380 6683 6383
rect 6633 6367 6647 6372
rect 6673 6367 6687 6380
rect 6736 6307 6743 6433
rect 6716 6247 6723 6293
rect 6756 6267 6763 6473
rect 6776 6428 6783 6453
rect 6816 6367 6823 6553
rect 6836 6507 6843 6593
rect 6856 6567 6863 6603
rect 6916 6527 6923 6613
rect 6836 6423 6843 6493
rect 6936 6487 6943 6653
rect 7033 6640 7047 6653
rect 7036 6636 7043 6640
rect 7027 6443 7040 6447
rect 7027 6440 7043 6443
rect 7027 6433 7047 6440
rect 6836 6416 6863 6423
rect 7033 6427 7047 6433
rect 6616 6043 6623 6114
rect 6636 6047 6643 6213
rect 6716 6163 6723 6193
rect 6736 6187 6743 6213
rect 6716 6156 6743 6163
rect 6676 6080 6683 6083
rect 6673 6067 6687 6080
rect 6596 6036 6623 6043
rect 6596 6027 6603 6036
rect 6576 5647 6583 5732
rect 6556 5636 6573 5643
rect 6536 5207 6543 5473
rect 6533 5127 6547 5133
rect 6520 5083 6533 5087
rect 6516 5076 6533 5083
rect 6436 4927 6443 5076
rect 6520 5073 6533 5076
rect 6456 4883 6463 5033
rect 6476 4888 6483 5013
rect 6436 4876 6463 4883
rect 6436 4856 6443 4876
rect 6376 4526 6383 4593
rect 6396 4336 6403 4613
rect 6416 4607 6423 4812
rect 6516 4727 6523 4953
rect 6476 4568 6483 4693
rect 6516 4556 6523 4593
rect 6536 4583 6543 4793
rect 6556 4747 6563 5636
rect 6596 5623 6603 6013
rect 6656 5896 6663 5933
rect 6736 5867 6743 6156
rect 6756 6086 6763 6113
rect 6776 6027 6783 6353
rect 6876 6347 6883 6383
rect 6916 6347 6923 6383
rect 6876 6167 6883 6333
rect 6916 6187 6923 6233
rect 6936 6227 6943 6372
rect 6956 6267 6963 6383
rect 6636 5827 6643 5863
rect 6756 5866 6763 5953
rect 6776 5843 6783 5894
rect 6756 5836 6783 5843
rect 6616 5667 6623 5753
rect 6576 5616 6603 5623
rect 6576 5343 6583 5616
rect 6596 5560 6603 5563
rect 6593 5547 6607 5560
rect 6656 5527 6663 5563
rect 6696 5383 6703 5733
rect 6676 5376 6703 5383
rect 6576 5336 6603 5343
rect 6576 5167 6583 5193
rect 6576 5047 6583 5093
rect 6576 4827 6583 4854
rect 6556 4627 6563 4673
rect 6536 4576 6553 4583
rect 6556 4556 6563 4573
rect 6496 4367 6503 4523
rect 6536 4483 6543 4523
rect 6536 4476 6563 4483
rect 6416 4227 6423 4303
rect 6356 4006 6363 4213
rect 6496 4167 6503 4353
rect 6416 4036 6423 4153
rect 6436 3947 6443 4003
rect 6356 3816 6363 3853
rect 6476 3787 6483 3814
rect 6456 3776 6473 3783
rect 6456 3667 6463 3776
rect 6356 3507 6363 3633
rect 6316 3367 6323 3412
rect 6376 3407 6383 3613
rect 6433 3520 6447 3533
rect 6456 3527 6463 3653
rect 6436 3516 6443 3520
rect 6416 3387 6423 3483
rect 6516 3467 6523 4393
rect 6536 4348 6543 4413
rect 6556 4387 6563 4476
rect 6596 4407 6603 5336
rect 6656 5207 6663 5343
rect 6716 5327 6723 5813
rect 6736 5307 6743 5594
rect 6756 5327 6763 5836
rect 6776 5487 6783 5793
rect 6796 5747 6803 6153
rect 6907 6134 6913 6147
rect 6900 6133 6920 6134
rect 6853 6120 6867 6133
rect 6856 6116 6863 6120
rect 6816 6007 6823 6113
rect 6956 6027 6963 6133
rect 6976 6107 6983 6293
rect 6996 6227 7003 6293
rect 7056 6287 7063 6573
rect 6876 5896 6883 6013
rect 6796 5566 6803 5613
rect 6816 5527 6823 5853
rect 6856 5627 6863 5863
rect 6936 5647 6943 5993
rect 6876 5596 6883 5633
rect 6956 5627 6963 6013
rect 6976 5847 6983 5893
rect 6996 5866 7003 6113
rect 7016 6087 7023 6114
rect 7036 5967 7043 6253
rect 7056 5947 7063 6233
rect 7076 6127 7083 6953
rect 7096 6867 7103 6934
rect 7096 6587 7103 6853
rect 7116 6527 7123 6953
rect 7136 6507 7143 6934
rect 7136 6416 7143 6472
rect 7156 6467 7163 7053
rect 7176 6967 7183 7276
rect 7256 7247 7263 7423
rect 7196 6943 7203 7233
rect 7216 7027 7223 7073
rect 7176 6936 7203 6943
rect 7236 6936 7243 7053
rect 7276 7047 7283 7373
rect 7296 6967 7303 7693
rect 7316 7567 7323 7796
rect 7396 7747 7403 7943
rect 7480 7923 7493 7927
rect 7476 7913 7493 7923
rect 7436 7703 7443 7833
rect 7476 7827 7483 7913
rect 7436 7696 7463 7703
rect 7376 7640 7383 7643
rect 7136 6116 7143 6173
rect 7176 6127 7183 6936
rect 7216 6847 7223 6903
rect 7216 6647 7223 6753
rect 7256 6636 7263 6833
rect 7316 6783 7323 7493
rect 7356 7387 7363 7633
rect 7373 7627 7387 7640
rect 7376 7587 7383 7613
rect 7376 7287 7383 7453
rect 7396 7207 7403 7473
rect 7416 7467 7423 7513
rect 7436 7487 7443 7673
rect 7456 7627 7463 7696
rect 7476 7527 7483 7673
rect 7496 7587 7503 7833
rect 7456 7347 7463 7393
rect 7456 7223 7463 7333
rect 7476 7247 7483 7423
rect 7456 7216 7483 7223
rect 7456 7126 7463 7193
rect 7476 7168 7483 7216
rect 7436 7047 7443 7073
rect 7456 7027 7463 7112
rect 7496 7107 7503 7373
rect 7516 7347 7523 8113
rect 7576 8047 7583 8156
rect 7556 8036 7573 8043
rect 7556 7887 7563 8036
rect 7596 7976 7603 8053
rect 7636 7976 7643 8013
rect 7656 7940 7663 7943
rect 7653 7927 7667 7940
rect 7536 7876 7553 7883
rect 7536 7507 7543 7876
rect 7516 7307 7523 7333
rect 7336 6867 7343 6934
rect 7356 6907 7363 6993
rect 7376 6887 7383 7013
rect 7476 6987 7483 7033
rect 7516 7027 7523 7272
rect 7536 7127 7543 7472
rect 7556 7147 7563 7573
rect 7576 7547 7583 7643
rect 7616 7640 7623 7643
rect 7613 7627 7627 7640
rect 7576 7387 7583 7493
rect 7576 7163 7583 7313
rect 7596 7267 7603 7613
rect 7636 7487 7643 7633
rect 7676 7607 7683 7674
rect 7696 7627 7703 7713
rect 7716 7587 7723 8013
rect 7736 7647 7743 8053
rect 7696 7456 7703 7533
rect 7736 7467 7743 7612
rect 7756 7487 7763 8073
rect 7776 7907 7783 7974
rect 7796 7747 7803 8073
rect 7836 8067 7843 8373
rect 7876 8087 7883 8183
rect 7896 8027 7903 8313
rect 7936 8303 7943 8333
rect 8096 8327 8103 8476
rect 7936 8296 7963 8303
rect 7936 7956 7943 8133
rect 7956 8047 7963 8296
rect 7976 8147 7983 8313
rect 8136 8287 8143 8393
rect 8196 8196 8203 8293
rect 8096 8087 8103 8172
rect 8236 8167 8243 8493
rect 8256 8447 8263 8493
rect 8276 8447 8283 8933
rect 8316 8747 8323 8873
rect 8333 8748 8347 8753
rect 8176 8107 8183 8163
rect 7876 7647 7883 7893
rect 7896 7887 7903 7923
rect 8056 7767 8063 7963
rect 8076 7676 8083 7813
rect 7896 7547 7903 7613
rect 7916 7567 7923 7674
rect 8056 7640 8063 7643
rect 8053 7627 8067 7640
rect 7616 7223 7623 7453
rect 7716 7247 7723 7423
rect 7756 7400 7763 7403
rect 7736 7287 7743 7393
rect 7753 7387 7767 7400
rect 7727 7236 7743 7243
rect 7596 7216 7623 7223
rect 7596 7187 7603 7216
rect 7576 7156 7623 7163
rect 7520 6903 7533 6907
rect 7416 6787 7423 6893
rect 7436 6867 7443 6893
rect 7296 6776 7323 6783
rect 7296 6656 7303 6776
rect 7196 6086 7203 6513
rect 7216 6247 7223 6513
rect 7236 6367 7243 6603
rect 7276 6483 7283 6573
rect 7356 6527 7363 6713
rect 7456 6683 7463 6873
rect 7476 6747 7483 6903
rect 7516 6896 7533 6903
rect 7520 6893 7533 6896
rect 7556 6906 7563 6933
rect 7576 6807 7583 7113
rect 7596 6707 7603 7133
rect 7616 6907 7623 6933
rect 7436 6676 7463 6683
rect 7436 6627 7443 6676
rect 7453 6620 7467 6633
rect 7456 6616 7463 6620
rect 7596 6607 7603 6693
rect 7636 6687 7643 7073
rect 7656 6626 7663 6953
rect 7676 6947 7683 7083
rect 7716 6936 7723 6993
rect 7736 6967 7743 7236
rect 7756 6936 7763 7073
rect 7776 6967 7783 7253
rect 7816 7127 7823 7473
rect 7996 7156 8023 7163
rect 8016 7127 8023 7156
rect 7887 7123 7900 7127
rect 7887 7116 7903 7123
rect 7887 7113 7900 7116
rect 7796 7087 7803 7112
rect 7736 6867 7743 6903
rect 7636 6620 7643 6623
rect 7633 6607 7647 6620
rect 7256 6476 7283 6483
rect 6913 5600 6927 5613
rect 6916 5596 6923 5600
rect 6816 5487 6823 5513
rect 6856 5507 6863 5563
rect 6956 5527 6963 5613
rect 6776 5346 6783 5373
rect 6753 5267 6767 5273
rect 6796 5263 6803 5433
rect 6936 5347 6943 5374
rect 6787 5256 6803 5263
rect 6813 5267 6827 5273
rect 6696 5127 6703 5233
rect 6756 5187 6763 5232
rect 6636 4967 6643 5113
rect 6776 5103 6783 5253
rect 6796 5207 6803 5233
rect 6836 5127 6843 5311
rect 6776 5096 6803 5103
rect 6693 5080 6707 5092
rect 6696 5076 6703 5080
rect 6656 5047 6663 5073
rect 6616 4823 6623 4873
rect 6696 4856 6703 4993
rect 6716 4967 6723 5043
rect 6616 4816 6643 4823
rect 6616 4467 6623 4573
rect 6636 4547 6643 4816
rect 6676 4687 6683 4823
rect 6596 4336 6603 4372
rect 6556 3783 6563 4334
rect 6613 4287 6627 4292
rect 6616 4187 6623 4233
rect 6636 4227 6643 4253
rect 6616 4036 6623 4133
rect 6656 4047 6663 4173
rect 6696 4143 6703 4733
rect 6716 4647 6723 4823
rect 6756 4627 6763 5032
rect 6796 4927 6803 5013
rect 6816 4907 6823 5053
rect 6836 4667 6843 5063
rect 6736 4556 6743 4613
rect 6716 4167 6723 4453
rect 6736 4307 6743 4493
rect 6756 4347 6763 4523
rect 6696 4136 6723 4143
rect 6653 3947 6667 3953
rect 6696 3947 6703 4093
rect 6616 3816 6623 3853
rect 6556 3776 6583 3783
rect 6576 3503 6583 3776
rect 6636 3747 6643 3783
rect 6716 3547 6723 4136
rect 6736 3627 6743 4293
rect 6756 3967 6763 4193
rect 6756 3647 6763 3953
rect 6776 3907 6783 4093
rect 6796 4043 6803 4633
rect 6836 4483 6843 4613
rect 6856 4507 6863 5273
rect 6876 5267 6883 5343
rect 6916 5207 6923 5233
rect 6956 5227 6963 5353
rect 6976 5247 6983 5413
rect 6996 5187 7003 5393
rect 7016 5267 7023 5933
rect 7096 5896 7103 5973
rect 7116 5927 7123 6083
rect 7156 6027 7163 6083
rect 7013 5247 7027 5253
rect 7036 5207 7043 5613
rect 7136 5596 7143 5733
rect 7156 5627 7163 5913
rect 7176 5866 7183 5953
rect 7196 5847 7203 5894
rect 7056 5507 7063 5594
rect 7196 5567 7203 5713
rect 7076 5376 7083 5473
rect 7116 5383 7123 5563
rect 7156 5527 7163 5563
rect 7116 5376 7143 5383
rect 6936 5067 6943 5113
rect 6956 5056 6963 5133
rect 6896 4856 6903 4933
rect 6836 4476 6863 4483
rect 6856 4336 6863 4476
rect 6876 4387 6883 4812
rect 6956 4607 6963 4823
rect 6996 4767 7003 4854
rect 7016 4827 7023 4893
rect 6956 4556 6963 4593
rect 6896 4367 6903 4533
rect 6936 4487 6943 4523
rect 6916 4476 6933 4483
rect 6916 4343 6923 4476
rect 6896 4336 6923 4343
rect 6836 4300 6843 4303
rect 6876 4300 6883 4303
rect 6833 4287 6847 4300
rect 6873 4287 6887 4300
rect 6976 4287 6983 4512
rect 7016 4283 7023 4673
rect 7036 4307 7043 4553
rect 7096 4527 7103 5293
rect 7136 5127 7143 5376
rect 7116 5003 7123 5053
rect 7136 5027 7143 5063
rect 7156 5007 7163 5513
rect 7176 5107 7183 5253
rect 7116 4996 7143 5003
rect 7116 4847 7123 4973
rect 7136 4947 7143 4996
rect 7216 4887 7223 6113
rect 7236 5287 7243 6193
rect 7256 5947 7263 6476
rect 7276 5923 7283 6453
rect 7296 6347 7303 6453
rect 7356 6447 7363 6513
rect 7376 6416 7383 6453
rect 7356 6307 7363 6372
rect 7396 6347 7403 6383
rect 7436 6347 7443 6473
rect 7476 6387 7483 6513
rect 7496 6267 7503 6493
rect 7516 6447 7523 6513
rect 7516 6307 7523 6393
rect 7536 6267 7543 6414
rect 7356 6116 7363 6153
rect 7396 6116 7403 6233
rect 7556 6207 7563 6453
rect 7596 6416 7603 6513
rect 7716 6443 7723 6673
rect 7696 6436 7723 6443
rect 7696 6407 7703 6436
rect 7296 6047 7303 6093
rect 7336 6007 7343 6072
rect 7376 6063 7383 6083
rect 7376 6060 7403 6063
rect 7376 6056 7407 6060
rect 7393 6047 7407 6056
rect 7256 5916 7283 5923
rect 7256 5867 7263 5916
rect 7356 5896 7363 5953
rect 7376 5908 7383 6033
rect 7256 5383 7263 5653
rect 7276 5587 7283 5773
rect 7336 5727 7343 5863
rect 7296 5407 7303 5613
rect 7356 5596 7363 5733
rect 7396 5596 7403 5653
rect 7416 5623 7423 6073
rect 7516 6047 7523 6073
rect 7556 5983 7563 6153
rect 7636 6123 7643 6383
rect 7676 6356 7703 6363
rect 7696 6343 7703 6356
rect 7696 6336 7723 6343
rect 7656 6187 7663 6233
rect 7636 6116 7663 6123
rect 7556 5976 7583 5983
rect 7496 5683 7503 5933
rect 7576 5747 7583 5976
rect 7636 5947 7643 6013
rect 7616 5787 7623 5893
rect 7636 5867 7643 5912
rect 7636 5767 7643 5853
rect 7496 5676 7523 5683
rect 7416 5616 7433 5623
rect 7433 5600 7447 5613
rect 7493 5600 7507 5613
rect 7516 5607 7523 5676
rect 7436 5596 7443 5600
rect 7496 5596 7503 5600
rect 7256 5376 7283 5383
rect 7316 5376 7323 5553
rect 7376 5507 7383 5563
rect 7296 5267 7303 5343
rect 7336 5336 7363 5343
rect 7356 5247 7363 5336
rect 7236 4927 7243 5193
rect 7316 5147 7323 5233
rect 7416 5207 7423 5553
rect 7536 5483 7543 5653
rect 7616 5627 7623 5713
rect 7636 5687 7643 5713
rect 7656 5667 7663 6116
rect 7556 5507 7563 5613
rect 7536 5476 7563 5483
rect 7256 5007 7263 5063
rect 7153 4860 7167 4873
rect 7236 4863 7243 4892
rect 7276 4868 7283 4933
rect 7156 4856 7163 4860
rect 7216 4856 7243 4863
rect 7136 4647 7143 4823
rect 7236 4727 7243 4833
rect 7256 4563 7263 4834
rect 7276 4667 7283 4854
rect 7296 4687 7303 5113
rect 7316 5027 7323 5063
rect 7316 4947 7323 5013
rect 7316 4727 7323 4912
rect 7336 4887 7343 4973
rect 7356 4863 7363 5193
rect 7456 5187 7463 5453
rect 7476 5367 7483 5393
rect 7556 5376 7563 5476
rect 7656 5467 7663 5613
rect 7676 5407 7683 6333
rect 7696 6086 7703 6153
rect 7696 5866 7703 6013
rect 7716 5927 7723 6336
rect 7736 6207 7743 6793
rect 7796 6567 7803 6993
rect 7816 6507 7823 7113
rect 7836 6527 7843 7093
rect 7896 6636 7903 7013
rect 7956 6936 7963 6973
rect 7993 6940 8007 6953
rect 7996 6936 8003 6940
rect 7936 6787 7943 6903
rect 7976 6867 7983 6903
rect 8036 6887 8043 6953
rect 7976 6648 7983 6853
rect 7960 6603 7973 6607
rect 7916 6507 7923 6603
rect 7956 6596 7973 6603
rect 7960 6593 7973 6596
rect 7996 6567 8003 6873
rect 7836 6400 7843 6403
rect 7833 6387 7847 6400
rect 8016 6396 8023 6593
rect 7736 6067 7743 6172
rect 7756 6087 7763 6253
rect 7856 6128 7863 6153
rect 7776 6083 7783 6114
rect 7776 6076 7803 6083
rect 7756 5896 7763 5973
rect 7796 5908 7803 6076
rect 7836 6027 7843 6083
rect 7816 5907 7823 5953
rect 7776 5860 7783 5863
rect 7773 5847 7787 5860
rect 7816 5827 7823 5853
rect 7836 5847 7843 5992
rect 7856 5827 7863 5894
rect 7696 5447 7703 5753
rect 7696 5387 7703 5433
rect 7716 5346 7723 5433
rect 7536 5207 7543 5343
rect 7576 5287 7583 5343
rect 7736 5287 7743 5552
rect 7756 5547 7763 5633
rect 7816 5596 7823 5733
rect 7856 5687 7863 5713
rect 7876 5647 7883 5893
rect 7796 5560 7803 5563
rect 7793 5547 7807 5560
rect 7836 5447 7843 5563
rect 7896 5527 7903 6193
rect 7916 5507 7923 6253
rect 7976 6247 7983 6393
rect 7956 5907 7963 6153
rect 7996 5967 8003 6353
rect 8036 6267 8043 6513
rect 8056 6467 8063 7533
rect 8076 7447 8083 7553
rect 8096 7547 8103 7674
rect 8116 7527 8123 7733
rect 8136 7607 8143 7753
rect 8116 7483 8123 7513
rect 8096 7476 8123 7483
rect 8096 7436 8103 7476
rect 8116 7407 8123 7453
rect 8156 7436 8163 7553
rect 8076 7127 8083 7393
rect 8096 7103 8103 7373
rect 8116 7107 8123 7333
rect 8176 7287 8183 7613
rect 8196 7327 8203 8033
rect 8236 7956 8243 8013
rect 8216 7387 8223 7913
rect 8256 7727 8263 8033
rect 8276 7987 8283 8353
rect 8296 8147 8303 8633
rect 8316 8467 8323 8573
rect 8336 8547 8343 8593
rect 8376 8496 8383 8753
rect 8396 8683 8403 8734
rect 8416 8707 8423 8813
rect 8436 8687 8443 9153
rect 8516 9016 8523 9173
rect 8536 9047 8543 9273
rect 8616 9248 8623 10053
rect 8756 10026 8763 10273
rect 8656 9967 8663 10023
rect 8836 9847 8843 10054
rect 8856 10026 8863 10532
rect 8996 10288 9003 10593
rect 9096 10588 9103 11113
rect 9173 11100 9187 11113
rect 9176 11096 9183 11100
rect 9633 11100 9647 11113
rect 9636 11096 9643 11100
rect 10256 11096 10263 11173
rect 9116 10766 9123 11033
rect 9156 10796 9163 10953
rect 9196 10887 9203 11063
rect 9236 10796 9243 10833
rect 9276 10766 9283 10873
rect 9356 10623 9363 11033
rect 9396 10796 9403 10873
rect 9416 10827 9423 11063
rect 9436 10796 9443 10833
rect 9476 10627 9483 11093
rect 9496 11066 9503 11093
rect 9616 10947 9623 11063
rect 9656 10796 9663 10893
rect 9576 10647 9583 10794
rect 9696 10787 9703 11052
rect 9356 10616 9373 10623
rect 9236 10576 9243 10613
rect 9036 10327 9043 10543
rect 9056 10246 9063 10453
rect 9096 10303 9103 10574
rect 9376 10546 9383 10613
rect 9256 10487 9263 10543
rect 9180 10303 9193 10307
rect 9087 10296 9103 10303
rect 9176 10293 9193 10303
rect 8936 10107 8943 10203
rect 8933 10060 8947 10072
rect 8936 10056 8943 10060
rect 8656 9720 8663 9723
rect 8653 9707 8667 9720
rect 8716 9707 8723 9773
rect 8896 9756 8903 9793
rect 8916 9787 8923 10023
rect 8796 9707 8803 9753
rect 8816 9723 8823 9754
rect 8816 9716 8843 9723
rect 8656 9506 8663 9693
rect 8776 9536 8783 9593
rect 8676 9303 8683 9533
rect 8796 9467 8803 9503
rect 8836 9467 8843 9716
rect 8916 9720 8923 9723
rect 8913 9707 8927 9720
rect 8976 9687 8983 10093
rect 9036 9727 9043 9754
rect 9056 9707 9063 10232
rect 9076 10087 9083 10293
rect 9176 10276 9183 10293
rect 9196 10207 9203 10243
rect 9236 10107 9243 10153
rect 9256 10147 9263 10473
rect 9316 10247 9323 10313
rect 9336 10227 9343 10433
rect 9376 10327 9383 10532
rect 9416 10327 9423 10613
rect 9576 10547 9583 10633
rect 9756 10547 9763 10813
rect 9520 10543 9533 10547
rect 9516 10536 9533 10543
rect 9520 10533 9533 10536
rect 9376 10276 9383 10313
rect 9420 10306 9433 10307
rect 9427 10293 9433 10306
rect 9396 10240 9403 10243
rect 9316 10216 9333 10223
rect 9076 9947 9083 10073
rect 9093 10067 9107 10073
rect 9173 10060 9187 10073
rect 9176 10056 9183 10060
rect 9296 10027 9303 10133
rect 9076 9723 9083 9933
rect 9116 9887 9123 10023
rect 9316 10007 9323 10216
rect 9356 10068 9363 10233
rect 9393 10227 9407 10240
rect 9396 10056 9403 10192
rect 9436 10187 9443 10243
rect 9376 10020 9383 10023
rect 9373 10007 9387 10020
rect 9416 9947 9423 10023
rect 9136 9756 9163 9763
rect 9076 9716 9103 9723
rect 9156 9707 9163 9756
rect 8916 9506 8923 9633
rect 8656 9296 8683 9303
rect 8613 9187 8627 9192
rect 8636 9163 8643 9293
rect 8616 9156 8643 9163
rect 8556 9016 8563 9093
rect 8616 9008 8623 9156
rect 8656 9087 8663 9296
rect 8936 9287 8943 9673
rect 8976 9536 8983 9652
rect 9016 9587 9023 9693
rect 9036 9467 9043 9503
rect 9016 9236 9023 9273
rect 8916 9187 8923 9234
rect 9056 9227 9063 9253
rect 8716 9156 8743 9163
rect 8456 8827 8463 8994
rect 8536 8887 8543 8983
rect 8576 8947 8583 8983
rect 8396 8676 8423 8683
rect 8416 8507 8423 8676
rect 8436 8488 8443 8513
rect 8456 8507 8463 8713
rect 8296 7956 8303 8013
rect 8316 7927 8323 8432
rect 8476 8347 8483 8793
rect 8496 8476 8503 8673
rect 8596 8667 8603 8714
rect 8516 8487 8523 8613
rect 8596 8587 8603 8653
rect 8616 8627 8623 8913
rect 8656 8847 8663 9033
rect 8676 8996 8683 9133
rect 8696 9007 8703 9073
rect 8716 8927 8723 9133
rect 8736 9107 8743 9156
rect 8860 9003 8873 9007
rect 8856 8996 8873 9003
rect 8860 8993 8873 8996
rect 8673 8827 8687 8833
rect 8696 8807 8703 8853
rect 8713 8827 8727 8833
rect 8736 8716 8743 8753
rect 8773 8720 8787 8733
rect 8776 8716 8783 8720
rect 8756 8587 8763 8683
rect 8796 8647 8803 8683
rect 8856 8647 8863 8973
rect 8956 8947 8963 9203
rect 8976 8996 8983 9033
rect 8996 9007 9003 9153
rect 9076 9067 9083 9553
rect 9096 9147 9103 9693
rect 9233 9540 9247 9553
rect 9236 9536 9243 9540
rect 9276 9536 9283 9573
rect 9476 9567 9483 10313
rect 9216 9487 9223 9503
rect 9213 9467 9227 9473
rect 9056 8967 9063 9013
rect 9116 9008 9123 9433
rect 9136 9127 9143 9453
rect 9196 9236 9203 9293
rect 9316 9267 9323 9533
rect 9416 9506 9423 9553
rect 9496 9548 9503 10413
rect 9776 10327 9783 11094
rect 9856 11060 9863 11063
rect 9853 11047 9867 11060
rect 9896 11007 9903 11063
rect 9796 10727 9803 10893
rect 9853 10800 9867 10813
rect 9856 10796 9863 10800
rect 9936 10767 9943 10833
rect 10096 10796 10103 10853
rect 10296 10796 10303 10933
rect 10356 10927 10363 11073
rect 10376 11066 10383 11093
rect 10456 11047 10463 11173
rect 10496 10987 10503 11063
rect 10536 11060 10543 11063
rect 10533 11047 10547 11060
rect 10636 11047 10643 11093
rect 10536 10887 10543 11033
rect 10516 10796 10523 10853
rect 10556 10808 10563 10833
rect 10376 10767 10383 10794
rect 9836 10727 9843 10763
rect 9856 10487 9863 10574
rect 10036 10547 10043 10574
rect 10056 10507 10063 10613
rect 10076 10543 10083 10653
rect 10316 10583 10323 10763
rect 10656 10766 10663 10973
rect 10676 10927 10683 11094
rect 10736 10987 10743 11063
rect 10776 11060 10783 11063
rect 10773 11047 10787 11060
rect 10676 10627 10683 10913
rect 10296 10576 10323 10583
rect 10076 10536 10093 10543
rect 10156 10507 10163 10543
rect 9593 10283 9607 10293
rect 9593 10280 9623 10283
rect 9596 10276 9623 10280
rect 9716 10236 9743 10243
rect 9736 10147 9743 10236
rect 9776 10147 9783 10313
rect 9516 9987 9523 10053
rect 9576 10023 9583 10093
rect 9613 10060 9627 10073
rect 9616 10056 9623 10060
rect 9576 10016 9603 10023
rect 9536 9756 9543 9813
rect 9576 9756 9583 9793
rect 9656 9768 9663 10023
rect 9776 9947 9783 10133
rect 9796 10087 9803 10273
rect 9836 10207 9843 10353
rect 9856 10246 9863 10473
rect 10296 10427 10303 10576
rect 10376 10540 10383 10543
rect 10373 10527 10387 10540
rect 10416 10527 10423 10613
rect 10536 10576 10543 10613
rect 10496 10546 10503 10573
rect 10556 10507 10563 10543
rect 10596 10447 10603 10532
rect 10156 10276 10203 10283
rect 9916 10187 9923 10243
rect 10056 10187 10063 10274
rect 9796 10026 9803 10073
rect 9896 10056 9903 10133
rect 9876 9987 9883 10023
rect 9696 9727 9703 9754
rect 9936 9727 9943 9813
rect 9956 9807 9963 10053
rect 10016 10026 10023 10173
rect 10136 10147 10143 10243
rect 10036 10007 10043 10133
rect 10196 10107 10203 10276
rect 10336 10187 10343 10243
rect 10136 10056 10143 10093
rect 10356 10056 10363 10213
rect 10376 10107 10383 10243
rect 10516 10107 10523 10353
rect 10556 10276 10563 10313
rect 10596 10276 10603 10353
rect 10636 10207 10643 10553
rect 10696 10546 10703 10973
rect 10816 10947 10823 11093
rect 10736 10796 10743 10873
rect 10767 10863 10780 10867
rect 10767 10853 10783 10863
rect 10776 10796 10783 10853
rect 11136 10847 11143 11094
rect 10796 10760 10803 10763
rect 10793 10747 10807 10760
rect 10896 10747 10903 10794
rect 10836 10627 10843 10693
rect 10836 10576 10843 10613
rect 10776 10540 10783 10543
rect 10596 10056 10603 10093
rect 10436 10026 10443 10053
rect 10076 10020 10083 10023
rect 10073 10007 10087 10020
rect 10036 9756 10043 9993
rect 10073 9987 10087 9993
rect 10296 9987 10303 10023
rect 9776 9687 9783 9723
rect 9447 9543 9460 9547
rect 9447 9536 9463 9543
rect 9447 9533 9460 9536
rect 9476 9500 9483 9503
rect 9416 9307 9423 9492
rect 9473 9487 9487 9500
rect 9533 9487 9547 9493
rect 9507 9363 9520 9367
rect 9507 9353 9523 9363
rect 9456 9236 9463 9293
rect 9216 9200 9223 9203
rect 9213 9187 9227 9200
rect 9376 9187 9383 9234
rect 9436 9200 9443 9203
rect 9433 9187 9447 9200
rect 9133 9000 9147 9013
rect 9136 8996 9143 9000
rect 9016 8927 9023 8963
rect 9056 8867 9063 8953
rect 8916 8687 8923 8714
rect 8536 8487 8543 8553
rect 8776 8476 8803 8483
rect 8336 7947 8343 8293
rect 8356 7887 8363 8153
rect 8376 8087 8383 8152
rect 8416 8107 8423 8163
rect 8276 7676 8283 7733
rect 8296 7727 8303 7773
rect 8236 7343 8243 7633
rect 8256 7367 8263 7643
rect 8236 7336 8263 7343
rect 8076 7096 8103 7103
rect 8076 6487 8083 7096
rect 8136 7007 8143 7273
rect 8176 7156 8183 7233
rect 8176 6987 8183 7093
rect 8176 6936 8183 6973
rect 8216 6936 8223 6993
rect 8236 6947 8243 7113
rect 8256 7107 8263 7336
rect 8276 7083 8283 7593
rect 8296 7367 8303 7513
rect 8256 7076 8283 7083
rect 8096 6587 8103 6733
rect 8256 6683 8263 7076
rect 8236 6676 8263 6683
rect 8096 6427 8103 6552
rect 8116 6547 8123 6593
rect 8136 6567 8143 6603
rect 8196 6587 8203 6623
rect 8076 6396 8103 6403
rect 8096 6327 8103 6396
rect 8116 6387 8123 6413
rect 8076 6128 8083 6293
rect 8116 6167 8123 6352
rect 8056 6080 8063 6083
rect 8053 6067 8067 6080
rect 8036 5908 8043 5953
rect 7936 5727 7943 5893
rect 8076 5866 8083 5953
rect 8096 5908 8103 6072
rect 7976 5787 7983 5863
rect 7936 5567 7943 5594
rect 7820 5426 7840 5427
rect 7820 5423 7833 5426
rect 7816 5413 7833 5423
rect 7816 5403 7823 5413
rect 7796 5396 7823 5403
rect 7796 5376 7803 5396
rect 7836 5343 7843 5392
rect 7816 5336 7843 5343
rect 7616 5207 7623 5233
rect 7596 5127 7603 5193
rect 7656 5096 7663 5233
rect 7493 5060 7507 5073
rect 7496 5056 7503 5060
rect 7696 4947 7703 5273
rect 7716 5007 7723 5073
rect 7756 5067 7763 5193
rect 7796 4947 7803 5233
rect 7336 4856 7363 4863
rect 7336 4826 7343 4856
rect 7416 4856 7423 4893
rect 7436 4667 7443 4823
rect 7247 4556 7263 4563
rect 7116 4467 7123 4554
rect 7093 4340 7107 4353
rect 7096 4336 7103 4340
rect 7076 4300 7083 4303
rect 7073 4287 7087 4300
rect 7016 4276 7043 4283
rect 6796 4036 6823 4043
rect 6856 4036 6863 4153
rect 6916 4007 6923 4053
rect 6936 4007 6943 4093
rect 6876 3967 6883 4003
rect 6956 4006 6963 4153
rect 6996 4107 7003 4233
rect 7036 4087 7043 4276
rect 7053 4267 7067 4273
rect 7116 4127 7123 4303
rect 7156 4207 7163 4273
rect 7176 4147 7183 4353
rect 7196 4227 7203 4373
rect 7093 4040 7107 4053
rect 7096 4036 7103 4040
rect 6807 3943 6820 3947
rect 6807 3933 6823 3943
rect 6816 3907 6823 3933
rect 6776 3687 6783 3853
rect 6796 3747 6803 3873
rect 6836 3816 6843 3853
rect 6536 3407 6543 3503
rect 6556 3496 6583 3503
rect 6556 3347 6563 3496
rect 6576 3303 6583 3453
rect 6556 3296 6583 3303
rect 6096 3027 6103 3173
rect 5996 2967 6003 2994
rect 6047 2963 6060 2967
rect 6047 2956 6063 2963
rect 6047 2953 6060 2956
rect 6096 2887 6103 2963
rect 6116 2827 6123 2853
rect 5976 2476 5983 2773
rect 6076 2747 6083 2774
rect 5996 2707 6003 2743
rect 6056 2740 6063 2743
rect 6053 2727 6067 2740
rect 6016 2476 6023 2713
rect 5996 2347 6003 2443
rect 5736 1736 5743 1773
rect 5756 1767 5763 1852
rect 5816 1743 5823 1923
rect 5816 1736 5843 1743
rect 5756 1687 5763 1703
rect 5673 1440 5687 1453
rect 5713 1440 5727 1453
rect 5676 1436 5683 1440
rect 5716 1436 5723 1440
rect 5576 1216 5603 1223
rect 5576 1007 5583 1216
rect 5676 1216 5683 1273
rect 5756 1187 5763 1673
rect 5776 1406 5783 1433
rect 5616 1007 5623 1183
rect 5696 1103 5703 1183
rect 5727 1113 5733 1127
rect 5676 1096 5703 1103
rect 5596 928 5603 993
rect 5396 347 5403 753
rect 5576 727 5583 883
rect 5476 716 5533 723
rect 5416 666 5423 713
rect 5476 708 5483 716
rect 5627 713 5633 727
rect 5496 627 5503 663
rect 5496 396 5503 433
rect 5556 427 5563 693
rect 5576 647 5583 673
rect 5476 360 5483 363
rect 5516 360 5523 363
rect 5473 347 5487 360
rect 5513 347 5527 360
rect 5536 327 5543 353
rect 5556 347 5563 413
rect 5656 366 5663 733
rect 5676 587 5683 1096
rect 5816 916 5823 1093
rect 5836 923 5843 1736
rect 5856 1706 5863 1813
rect 5876 1748 5883 2093
rect 5896 1926 5903 1953
rect 5916 1907 5923 2223
rect 5956 2220 5963 2223
rect 5953 2207 5967 2220
rect 5936 1867 5943 1993
rect 5956 1887 5963 2013
rect 5996 1963 6003 2253
rect 6016 2027 6023 2393
rect 6036 2107 6043 2443
rect 6076 2067 6083 2453
rect 6136 2307 6143 2773
rect 6156 2407 6163 3233
rect 6176 3067 6183 3263
rect 6216 3207 6223 3263
rect 6316 3246 6323 3273
rect 6416 3267 6423 3283
rect 6556 3267 6563 3296
rect 6596 3276 6603 3393
rect 6236 2966 6243 3013
rect 6316 2996 6323 3033
rect 6236 2776 6243 2893
rect 6176 2307 6183 2533
rect 6236 2476 6243 2513
rect 6276 2476 6283 2533
rect 6216 2367 6223 2443
rect 6316 2443 6323 2633
rect 6296 2436 6323 2443
rect 6136 2256 6143 2293
rect 6216 2227 6223 2254
rect 5976 1956 6003 1963
rect 6036 1956 6043 2033
rect 6076 2007 6083 2053
rect 5896 1507 5903 1853
rect 5916 1467 5923 1753
rect 5936 1467 5943 1793
rect 5976 1767 5983 1956
rect 5996 1736 6003 1793
rect 6016 1787 6023 1813
rect 6056 1716 6063 1813
rect 5976 1700 5983 1703
rect 5973 1687 5987 1700
rect 6096 1686 6103 1873
rect 6116 1716 6123 1993
rect 6136 1787 6143 1953
rect 5906 1453 5907 1460
rect 5893 1440 5907 1453
rect 5896 1436 5903 1440
rect 5896 1216 5903 1293
rect 5956 1186 5963 1453
rect 5853 1107 5867 1113
rect 5876 927 5883 1183
rect 5916 967 5923 1183
rect 5976 1087 5983 1633
rect 5996 1507 6003 1613
rect 5996 1406 6003 1453
rect 5836 916 5863 923
rect 5796 747 5803 883
rect 5696 547 5703 663
rect 5756 660 5763 663
rect 5753 647 5767 660
rect 5776 627 5783 694
rect 5476 176 5483 233
rect 5516 176 5523 253
rect 5656 127 5663 352
rect 5756 188 5763 533
rect 5856 447 5863 916
rect 5936 827 5943 1053
rect 5976 1007 5983 1073
rect 5976 916 5983 993
rect 6036 967 6043 1573
rect 6076 1307 6083 1403
rect 6093 1220 6107 1233
rect 6096 1216 6103 1220
rect 6136 1216 6143 1313
rect 6156 1247 6163 2053
rect 6176 1927 6183 1993
rect 6236 1967 6243 2253
rect 6276 1956 6283 2173
rect 6296 2067 6303 2436
rect 6316 2223 6323 2373
rect 6336 2267 6343 2963
rect 6416 2927 6423 3253
rect 6516 2883 6523 2963
rect 6516 2876 6543 2883
rect 6536 2827 6543 2876
rect 6396 2647 6403 2793
rect 6453 2780 6467 2793
rect 6456 2776 6463 2780
rect 6416 2627 6423 2774
rect 6536 2747 6543 2813
rect 6356 2256 6363 2293
rect 6316 2216 6343 2223
rect 6216 1926 6223 1953
rect 6216 1827 6223 1912
rect 6336 1827 6343 2216
rect 6376 1926 6383 2223
rect 6416 2067 6423 2613
rect 6476 2476 6483 2653
rect 6436 1867 6443 2413
rect 6456 2047 6463 2443
rect 6476 2147 6483 2273
rect 6496 2267 6503 2443
rect 6536 2288 6543 2493
rect 6596 2447 6603 3073
rect 6616 2307 6623 3333
rect 6676 3283 6683 3313
rect 6656 3276 6683 3283
rect 6696 3187 6703 3373
rect 6716 3267 6723 3293
rect 6736 2996 6743 3033
rect 6636 2966 6643 2993
rect 6756 2927 6763 2963
rect 6716 2776 6723 2913
rect 6636 2547 6643 2774
rect 6736 2607 6743 2743
rect 6716 2476 6723 2533
rect 6796 2523 6803 3393
rect 6816 3327 6823 3633
rect 6876 3536 6883 3573
rect 6876 3367 6883 3413
rect 6916 3387 6923 3953
rect 6833 3300 6847 3313
rect 6836 3296 6843 3300
rect 6836 2747 6843 2813
rect 6856 2746 6863 3263
rect 6876 2667 6883 3253
rect 6936 3167 6943 3533
rect 6976 3267 6983 4034
rect 7036 3967 7043 3993
rect 6996 3767 7003 3814
rect 7116 3787 7123 3814
rect 7136 3807 7143 3873
rect 7056 3767 7063 3783
rect 7156 3767 7163 4113
rect 7056 3756 7073 3767
rect 7060 3753 7073 3756
rect 7133 3727 7147 3733
rect 7176 3723 7183 4073
rect 7196 3747 7203 4192
rect 7216 4007 7223 4453
rect 7236 4287 7243 4554
rect 7256 3867 7263 4532
rect 7276 4527 7283 4593
rect 7296 4303 7303 4633
rect 7316 4547 7323 4653
rect 7416 4556 7423 4593
rect 7336 4407 7343 4493
rect 7356 4467 7363 4523
rect 7396 4467 7403 4523
rect 7336 4336 7343 4393
rect 7436 4307 7443 4513
rect 7456 4307 7463 4713
rect 7296 4296 7323 4303
rect 7293 4207 7307 4213
rect 7276 4036 7283 4153
rect 7356 4147 7363 4293
rect 7336 4036 7363 4043
rect 7356 3927 7363 4036
rect 7376 4007 7383 4253
rect 7276 3816 7283 3913
rect 7336 3807 7343 3873
rect 7396 3827 7403 4273
rect 7256 3780 7263 3783
rect 7253 3767 7267 3780
rect 7176 3716 7203 3723
rect 6996 3047 7003 3673
rect 7016 3323 7023 3573
rect 7036 3507 7043 3633
rect 7076 3516 7083 3653
rect 7096 3480 7103 3483
rect 7093 3467 7107 3480
rect 7156 3467 7163 3514
rect 7036 3407 7043 3453
rect 7016 3316 7033 3323
rect 7033 3300 7047 3313
rect 7036 3296 7043 3300
rect 7136 3266 7143 3293
rect 7056 3227 7063 3263
rect 6916 3003 6923 3033
rect 6916 2996 6943 3003
rect 7036 2956 7063 2963
rect 6936 2776 6943 2833
rect 6907 2743 6920 2747
rect 6996 2746 7003 2913
rect 6907 2736 6923 2743
rect 6907 2733 6920 2736
rect 7016 2627 7023 2753
rect 7056 2687 7063 2956
rect 7076 2627 7083 3153
rect 7156 2776 7163 3133
rect 7176 3087 7183 3613
rect 7196 2943 7203 3716
rect 7216 2996 7223 3333
rect 7236 3147 7243 3753
rect 7296 3727 7303 3783
rect 7256 3303 7263 3553
rect 7336 3516 7343 3693
rect 7396 3667 7403 3813
rect 7316 3407 7323 3483
rect 7356 3347 7363 3472
rect 7256 3296 7283 3303
rect 7296 3260 7303 3263
rect 7293 3247 7307 3260
rect 7376 3247 7383 3313
rect 7256 2960 7263 2963
rect 7253 2947 7267 2960
rect 7196 2936 7223 2943
rect 7216 2747 7223 2936
rect 6796 2516 6823 2523
rect 6773 2503 6787 2513
rect 6767 2500 6787 2503
rect 6767 2496 6783 2500
rect 6816 2466 6823 2516
rect 6676 2440 6683 2443
rect 6673 2427 6687 2440
rect 6796 2347 6803 2463
rect 6916 2456 6923 2493
rect 6496 2087 6503 2253
rect 6636 2236 6643 2313
rect 6656 2227 6663 2273
rect 6596 2147 6603 2203
rect 6553 2047 6567 2053
rect 6476 1956 6483 1993
rect 6576 1923 6583 1954
rect 6496 1843 6503 1923
rect 6476 1836 6503 1843
rect 6476 1726 6483 1836
rect 6396 1716 6423 1723
rect 6396 1567 6403 1716
rect 6296 1448 6303 1473
rect 6336 1436 6343 1493
rect 6456 1487 6463 1672
rect 6056 916 6063 1033
rect 6096 907 6103 1133
rect 6136 1127 6143 1153
rect 6156 1107 6163 1183
rect 5953 700 5967 713
rect 5956 696 5963 700
rect 6036 687 6043 872
rect 6116 787 6123 973
rect 6136 747 6143 1073
rect 6196 886 6203 1273
rect 6216 1147 6223 1253
rect 6247 1153 6253 1167
rect 6276 947 6283 1233
rect 6296 916 6303 1293
rect 6353 1220 6367 1233
rect 6356 1216 6363 1220
rect 6336 1107 6343 1183
rect 6336 1067 6343 1093
rect 6196 723 6203 872
rect 6176 716 6203 723
rect 6176 696 6183 716
rect 6216 696 6223 813
rect 6236 807 6243 883
rect 6316 880 6323 883
rect 6313 867 6327 880
rect 5976 660 5983 663
rect 5973 647 5987 660
rect 6276 666 6283 733
rect 5996 623 6003 653
rect 5947 616 6003 623
rect 5956 396 5963 433
rect 5996 367 6003 394
rect 5896 267 5903 363
rect 5936 327 5943 363
rect 5893 188 5907 193
rect 5956 183 5963 293
rect 5936 176 5963 183
rect 5856 147 5863 174
rect 6016 147 6023 633
rect 6156 396 6163 663
rect 6213 627 6227 633
rect 6226 620 6227 627
rect 6236 367 6243 613
rect 6180 363 6193 367
rect 6136 207 6143 363
rect 6176 356 6193 363
rect 6180 353 6193 356
rect 6140 183 6153 187
rect 6136 176 6153 183
rect 6140 173 6153 176
rect 6276 147 6283 313
rect 6316 267 6323 793
rect 6356 747 6363 914
rect 6376 666 6383 933
rect 6436 886 6443 1393
rect 6476 1287 6483 1493
rect 6476 1107 6483 1214
rect 6496 916 6503 1813
rect 6516 1436 6523 1633
rect 6536 1527 6543 1923
rect 6556 1916 6583 1923
rect 6556 1887 6563 1916
rect 6556 1707 6563 1873
rect 6576 1607 6583 1733
rect 6576 1403 6583 1593
rect 6556 1396 6583 1403
rect 6596 1307 6603 1913
rect 6616 1228 6623 2073
rect 6676 1926 6683 2033
rect 6736 1956 6743 2033
rect 6756 1987 6763 2243
rect 6776 1956 6783 2133
rect 6896 2087 6903 2333
rect 6933 2240 6947 2253
rect 6956 2248 6963 2293
rect 6936 2236 6943 2240
rect 6956 2147 6963 2234
rect 6656 1736 6663 1773
rect 6816 1767 6823 2033
rect 6836 1847 6843 1973
rect 6876 1927 6883 1954
rect 6693 1740 6707 1753
rect 6696 1736 6703 1740
rect 6896 1736 6903 2013
rect 6916 1887 6923 2053
rect 7016 2027 7023 2333
rect 6993 1960 7007 1973
rect 6996 1956 7003 1960
rect 6976 1847 6983 1923
rect 7016 1767 7023 1923
rect 6636 1307 6643 1693
rect 6676 1647 6683 1703
rect 6876 1683 6883 1703
rect 6876 1676 6903 1683
rect 6756 1436 6763 1533
rect 6896 1467 6903 1676
rect 6916 1647 6923 1703
rect 6793 1440 6807 1453
rect 6796 1436 6803 1440
rect 6776 1367 6783 1403
rect 6816 1400 6823 1403
rect 6813 1387 6827 1400
rect 6856 1367 6863 1453
rect 6916 1443 6923 1612
rect 6896 1436 6923 1443
rect 6556 1180 6563 1183
rect 6553 1167 6567 1180
rect 6616 1087 6623 1214
rect 6776 1216 6783 1293
rect 6656 1187 6663 1213
rect 6756 1147 6763 1183
rect 6476 727 6483 872
rect 6516 708 6523 883
rect 6556 880 6563 883
rect 6553 867 6567 880
rect 6556 807 6563 853
rect 6596 767 6603 914
rect 6616 807 6623 973
rect 6756 916 6763 953
rect 6696 767 6703 853
rect 6416 647 6423 663
rect 6407 636 6423 647
rect 6407 633 6420 636
rect 6336 396 6363 403
rect 6336 207 6343 396
rect 6476 367 6483 394
rect 6356 247 6363 273
rect 6356 176 6363 233
rect 6416 146 6423 173
rect 6436 87 6443 352
rect 6536 176 6543 393
rect 6556 367 6563 753
rect 6613 700 6627 713
rect 6616 696 6623 700
rect 6696 696 6703 753
rect 6736 723 6743 883
rect 6736 716 6763 723
rect 6596 408 6603 533
rect 6636 396 6643 493
rect 6736 467 6743 693
rect 6756 607 6763 716
rect 6776 666 6783 813
rect 6816 687 6823 713
rect 6836 607 6843 1172
rect 6856 886 6863 1013
rect 6896 696 6903 1436
rect 6936 1147 6943 1553
rect 6956 1427 6963 1733
rect 6996 1507 7003 1693
rect 7016 1687 7023 1753
rect 7056 1627 7063 2593
rect 7136 2547 7143 2743
rect 7156 2567 7163 2593
rect 7107 2456 7123 2463
rect 7076 2267 7083 2393
rect 7076 1747 7083 1953
rect 7096 1736 7103 2273
rect 7116 1847 7123 2456
rect 7176 2443 7183 2732
rect 7156 2436 7183 2443
rect 7136 1927 7143 2212
rect 7156 2187 7163 2436
rect 7196 2343 7203 2493
rect 7216 2466 7223 2673
rect 7216 2367 7223 2452
rect 7236 2407 7243 2853
rect 7256 2446 7263 2933
rect 7276 2927 7283 3133
rect 7196 2336 7223 2343
rect 7216 2256 7223 2336
rect 7256 2256 7263 2293
rect 7276 2283 7283 2873
rect 7296 2307 7303 2593
rect 7316 2587 7323 2952
rect 7416 2887 7423 4293
rect 7436 3627 7443 4233
rect 7456 3827 7463 4272
rect 7476 3867 7483 4673
rect 7516 4423 7523 4893
rect 7536 4836 7543 4933
rect 7576 4827 7583 4933
rect 7716 4836 7743 4843
rect 7556 4467 7563 4793
rect 7596 4556 7603 4653
rect 7496 4416 7523 4423
rect 7496 4387 7503 4416
rect 7616 4407 7623 4523
rect 7716 4487 7723 4813
rect 7736 4807 7743 4836
rect 7816 4747 7823 5336
rect 7856 5327 7863 5493
rect 7956 5467 7963 5773
rect 7967 5456 7983 5463
rect 7876 5247 7883 5373
rect 7896 5346 7903 5413
rect 7976 5383 7983 5456
rect 7996 5427 8003 5633
rect 8036 5608 8043 5813
rect 8076 5747 8083 5852
rect 8096 5663 8103 5894
rect 8116 5787 8123 6013
rect 8096 5656 8123 5663
rect 8076 5596 8083 5633
rect 7956 5376 7983 5383
rect 8016 5376 8023 5553
rect 8056 5388 8063 5473
rect 7836 5107 7843 5153
rect 7896 5076 7903 5332
rect 7956 5323 7963 5376
rect 8036 5327 8043 5343
rect 7956 5316 7983 5323
rect 7876 5040 7883 5043
rect 7836 4836 7843 5033
rect 7873 5027 7887 5040
rect 7916 4987 7923 5033
rect 7936 5027 7943 5074
rect 7916 4806 7923 4933
rect 7816 4556 7823 4613
rect 7876 4568 7883 4713
rect 7796 4520 7803 4523
rect 7793 4507 7807 4520
rect 7856 4487 7863 4523
rect 7516 4048 7523 4393
rect 7536 4306 7543 4373
rect 7556 4036 7563 4073
rect 7596 3987 7603 4034
rect 7616 4027 7623 4113
rect 7676 4067 7683 4473
rect 7836 4336 7843 4373
rect 7696 4307 7703 4334
rect 7816 4127 7823 4292
rect 7856 4227 7863 4292
rect 7896 4247 7903 4693
rect 7936 4307 7943 4933
rect 7956 4407 7963 5293
rect 7976 4907 7983 5316
rect 8016 5316 8033 5323
rect 7976 4167 7983 4593
rect 7996 4487 8003 5311
rect 8016 5127 8023 5316
rect 8016 4707 8023 5113
rect 8036 5047 8043 5292
rect 8096 5227 8103 5513
rect 8116 5487 8123 5656
rect 8116 5076 8123 5413
rect 8136 5347 8143 6473
rect 8156 5623 8163 5973
rect 8176 5687 8183 6533
rect 8216 6386 8223 6613
rect 8236 6167 8243 6676
rect 8276 6667 8283 6973
rect 8256 6620 8263 6623
rect 8253 6607 8267 6620
rect 8296 6447 8303 6993
rect 8316 6907 8323 7753
rect 8336 7607 8343 7833
rect 8356 7468 8363 7773
rect 8376 7647 8383 7973
rect 8416 7567 8423 8093
rect 8436 7847 8443 8153
rect 8456 7827 8463 8253
rect 8496 8167 8503 8373
rect 8536 8343 8543 8452
rect 8536 8336 8563 8343
rect 8496 7976 8503 8013
rect 8536 7988 8543 8273
rect 8556 8147 8563 8336
rect 8593 8200 8607 8213
rect 8596 8196 8603 8200
rect 8676 8196 8683 8293
rect 8476 7807 8483 7833
rect 8516 7707 8523 7943
rect 8473 7680 8487 7693
rect 8536 7683 8543 7773
rect 8476 7676 8483 7680
rect 8516 7676 8543 7683
rect 8456 7640 8463 7643
rect 8453 7627 8467 7640
rect 8376 7487 8383 7553
rect 8420 7423 8433 7427
rect 8376 7347 8383 7423
rect 8416 7416 8433 7423
rect 8420 7413 8433 7416
rect 8376 7167 8383 7273
rect 8416 7267 8423 7393
rect 8416 7156 8423 7253
rect 8436 7227 8443 7333
rect 8456 7176 8463 7493
rect 8476 7387 8483 7453
rect 8336 6787 8343 7093
rect 8396 7067 8403 7123
rect 8496 7027 8503 7093
rect 8393 6940 8407 6953
rect 8516 6947 8523 7553
rect 8556 7487 8563 7673
rect 8576 7646 8583 7973
rect 8576 7587 8583 7632
rect 8596 7567 8603 8133
rect 8716 7976 8723 8333
rect 8776 8327 8783 8476
rect 8856 8287 8863 8413
rect 8876 8387 8883 8593
rect 8893 8480 8907 8493
rect 8936 8483 8943 8853
rect 9116 8847 9123 8994
rect 9016 8716 9023 8773
rect 9176 8747 9183 9053
rect 9196 8716 9223 8723
rect 9196 8686 9203 8716
rect 8996 8486 9003 8683
rect 9033 8667 9047 8672
rect 9276 8663 9283 8833
rect 9256 8656 9283 8663
rect 8896 8476 8903 8480
rect 8936 8476 8963 8483
rect 8756 8107 8763 8213
rect 8796 8067 8803 8233
rect 8916 8196 8923 8233
rect 8936 8207 8943 8476
rect 9256 8476 9263 8656
rect 9336 8407 9343 8873
rect 9356 8446 9363 8493
rect 8996 8186 9003 8293
rect 9196 8176 9203 8313
rect 9356 8216 9363 8393
rect 9396 8267 9403 8853
rect 9416 8716 9423 9113
rect 9516 9107 9523 9353
rect 9436 8996 9443 9093
rect 9536 9003 9543 9273
rect 9556 9206 9563 9233
rect 9576 9123 9583 9573
rect 9713 9540 9727 9553
rect 9716 9536 9723 9540
rect 9696 9447 9703 9503
rect 9556 9116 9583 9123
rect 9556 9006 9563 9116
rect 9516 8996 9543 9003
rect 9476 8927 9483 8952
rect 9436 8307 9443 8494
rect 9013 8167 9027 8172
rect 8856 8160 8863 8163
rect 8896 8160 8903 8163
rect 8836 8127 8843 8152
rect 8853 8147 8867 8160
rect 8893 8147 8907 8160
rect 8816 7947 8823 8013
rect 8836 7988 8843 8013
rect 8736 7940 8743 7943
rect 8636 7527 8643 7933
rect 8733 7927 8747 7940
rect 8776 7936 8803 7943
rect 8733 7680 8747 7693
rect 8736 7676 8743 7680
rect 8536 7427 8543 7453
rect 8556 7426 8563 7473
rect 8636 7420 8643 7423
rect 8633 7407 8647 7420
rect 8696 7307 8703 7454
rect 8716 7407 8723 7493
rect 8396 6936 8403 6940
rect 8576 6936 8583 7013
rect 8596 7007 8603 7033
rect 8636 6847 8643 6903
rect 8536 6567 8543 6813
rect 8596 6656 8603 6713
rect 8636 6623 8643 6653
rect 8556 6448 8563 6623
rect 8616 6616 8643 6623
rect 8296 6380 8303 6383
rect 8293 6367 8307 6380
rect 8336 6247 8343 6372
rect 8293 6120 8307 6133
rect 8296 6116 8303 6120
rect 8216 5908 8223 5993
rect 8256 5896 8263 6013
rect 8276 5967 8283 6083
rect 8336 6067 8343 6114
rect 8196 5787 8203 5853
rect 8236 5767 8243 5863
rect 8276 5843 8283 5852
rect 8256 5836 8283 5843
rect 8256 5647 8263 5836
rect 8156 5616 8183 5623
rect 8156 5527 8163 5594
rect 8096 4927 8103 5043
rect 8136 5023 8143 5032
rect 8116 5016 8143 5023
rect 8116 4887 8123 5016
rect 8073 4860 8087 4873
rect 8076 4856 8083 4860
rect 8116 4856 8123 4873
rect 8136 4867 8143 4913
rect 8076 4556 8083 4733
rect 8096 4607 8103 4823
rect 8156 4767 8163 4893
rect 8176 4643 8183 5616
rect 8196 5567 8203 5613
rect 8233 5600 8247 5613
rect 8236 5596 8243 5600
rect 8276 5596 8283 5773
rect 8196 5307 8203 5513
rect 8256 5427 8263 5563
rect 8296 5527 8303 5563
rect 8296 5387 8303 5413
rect 8280 5343 8293 5347
rect 8156 4636 8183 4643
rect 8113 4560 8127 4573
rect 8116 4556 8123 4560
rect 8016 4526 8023 4553
rect 8056 4336 8063 4473
rect 8096 4343 8103 4523
rect 8096 4336 8123 4343
rect 8036 4187 8043 4303
rect 7556 3787 7563 3973
rect 7436 3187 7443 3393
rect 7456 3167 7463 3773
rect 7476 3087 7483 3693
rect 7496 3647 7503 3713
rect 7576 3587 7583 3814
rect 7596 3747 7603 3893
rect 7616 3827 7623 3913
rect 7516 3516 7523 3573
rect 7536 3308 7543 3433
rect 7596 3387 7603 3514
rect 7560 3266 7573 3267
rect 7516 3227 7523 3263
rect 7567 3253 7573 3266
rect 7596 3247 7603 3293
rect 7473 3000 7487 3013
rect 7476 2996 7483 3000
rect 7393 2780 7407 2793
rect 7396 2776 7403 2780
rect 7456 2768 7463 2913
rect 7276 2276 7303 2283
rect 7176 1956 7183 1993
rect 7216 1968 7223 2173
rect 7296 2087 7303 2276
rect 7136 1736 7143 1873
rect 7196 1787 7203 1912
rect 7256 1867 7263 1993
rect 7256 1767 7263 1793
rect 6996 1436 7003 1493
rect 7033 1440 7047 1453
rect 7036 1436 7043 1440
rect 7016 1400 7023 1403
rect 7013 1387 7027 1400
rect 7053 1347 7067 1353
rect 6993 1220 7007 1233
rect 6996 1216 7003 1220
rect 6936 883 6943 1133
rect 6976 1127 6983 1183
rect 7016 1087 7023 1183
rect 7056 947 7063 1233
rect 7076 1167 7083 1434
rect 7096 1267 7103 1673
rect 7156 1607 7163 1703
rect 7276 1567 7283 1973
rect 7296 1527 7303 1973
rect 7316 1747 7323 2433
rect 7336 2323 7343 2613
rect 7356 2476 7363 2713
rect 7376 2707 7383 2743
rect 7416 2423 7423 2693
rect 7436 2527 7443 2713
rect 7396 2416 7423 2423
rect 7336 2316 7363 2323
rect 7336 2187 7343 2293
rect 7336 1923 7343 2133
rect 7356 2087 7363 2316
rect 7376 2067 7383 2173
rect 7396 2047 7403 2416
rect 7436 2283 7443 2353
rect 7456 2307 7463 2573
rect 7496 2503 7503 3153
rect 7516 2947 7523 3213
rect 7616 3147 7623 3813
rect 7516 2756 7523 2833
rect 7496 2496 7523 2503
rect 7436 2276 7463 2283
rect 7456 2256 7463 2276
rect 7373 1960 7387 1973
rect 7376 1956 7383 1960
rect 7416 1956 7423 2013
rect 7496 1947 7503 2473
rect 7336 1916 7363 1923
rect 7356 1736 7363 1916
rect 7436 1706 7443 1853
rect 7476 1707 7483 1734
rect 7336 1647 7343 1703
rect 7376 1567 7383 1703
rect 7256 1467 7263 1513
rect 7136 1327 7143 1433
rect 7156 1347 7163 1453
rect 7216 1383 7223 1403
rect 7216 1376 7243 1383
rect 7176 1327 7183 1353
rect 7236 1347 7243 1376
rect 7256 1267 7263 1403
rect 7236 1216 7243 1253
rect 7276 1187 7283 1214
rect 7216 1087 7223 1183
rect 6993 920 7007 933
rect 6996 916 7003 920
rect 7036 916 7083 923
rect 7076 887 7083 916
rect 6936 876 6963 883
rect 6776 327 6783 473
rect 6796 366 6803 493
rect 6816 396 6823 553
rect 6876 423 6883 663
rect 6956 663 6963 876
rect 6976 708 6983 883
rect 6936 656 6963 663
rect 6876 416 6903 423
rect 6796 188 6803 293
rect 6556 107 6563 143
rect 6596 136 6633 143
rect 6856 146 6863 233
rect 6816 67 6823 143
rect 6896 -24 6903 416
rect 6916 367 6923 394
rect 6936 107 6943 656
rect 6996 527 7003 753
rect 7016 747 7023 883
rect 7156 667 7163 813
rect 7116 660 7123 663
rect 7113 647 7127 660
rect 6956 287 6963 393
rect 7016 176 7023 433
rect 7056 396 7063 573
rect 7136 396 7143 433
rect 7076 327 7083 363
rect 6956 146 6963 173
rect 7036 27 7043 143
rect 7096 67 7103 253
rect 7176 146 7183 1073
rect 7296 1027 7303 1433
rect 7436 1400 7443 1403
rect 7433 1387 7447 1400
rect 7216 928 7223 953
rect 7253 920 7267 933
rect 7256 916 7263 920
rect 7296 847 7303 953
rect 7316 947 7323 1333
rect 7476 1223 7483 1693
rect 7496 1467 7503 1813
rect 7516 1748 7523 2496
rect 7556 2487 7563 3073
rect 7636 3027 7643 4053
rect 7727 4043 7740 4047
rect 7727 4036 7743 4043
rect 7727 4033 7740 4036
rect 7816 4047 7823 4113
rect 7656 3207 7663 3853
rect 7676 3827 7683 4032
rect 7696 3848 7703 4013
rect 7756 3927 7763 4003
rect 7816 3796 7823 3853
rect 7836 3807 7843 4153
rect 7956 4087 7963 4133
rect 7676 3527 7683 3773
rect 7716 3767 7723 3783
rect 7707 3753 7723 3767
rect 7696 3487 7703 3533
rect 7716 3528 7723 3753
rect 7796 3667 7803 3794
rect 7753 3520 7767 3533
rect 7756 3516 7763 3520
rect 7716 3447 7723 3473
rect 7736 3447 7743 3483
rect 7736 3407 7743 3433
rect 7796 3403 7803 3453
rect 7776 3396 7803 3403
rect 7776 3367 7783 3396
rect 7676 3267 7683 3353
rect 7713 3300 7727 3313
rect 7716 3296 7723 3300
rect 7796 3307 7803 3373
rect 7836 3283 7843 3573
rect 7856 3307 7863 4073
rect 7996 4036 8003 4173
rect 8076 4067 8083 4303
rect 8116 4287 8123 4336
rect 8116 4067 8123 4213
rect 8136 4147 8143 4334
rect 8033 4040 8047 4053
rect 8036 4036 8043 4040
rect 8076 4007 8083 4053
rect 8016 3967 8023 4003
rect 8156 3967 8163 4636
rect 8156 3827 8163 3953
rect 7996 3767 8003 3803
rect 8176 3803 8183 4613
rect 8196 4367 8203 5073
rect 8216 4627 8223 5333
rect 8236 4587 8243 5343
rect 8276 5336 8293 5343
rect 8280 5333 8293 5336
rect 8256 4827 8263 5253
rect 8276 4947 8283 5313
rect 8316 5088 8323 5373
rect 8336 5327 8343 5753
rect 8356 5547 8363 5673
rect 8356 5107 8363 5533
rect 8376 5427 8383 5594
rect 8396 5527 8403 6433
rect 8476 6387 8483 6414
rect 8576 6423 8583 6473
rect 8567 6416 8583 6423
rect 8476 6327 8483 6373
rect 8536 6367 8543 6383
rect 8527 6356 8543 6367
rect 8527 6353 8540 6356
rect 8596 6227 8603 6433
rect 8467 6143 8480 6147
rect 8467 6133 8483 6143
rect 8476 6116 8483 6133
rect 8456 6080 8463 6083
rect 8453 6067 8467 6080
rect 8496 6007 8503 6083
rect 8416 5856 8443 5863
rect 8416 5727 8423 5856
rect 8396 5327 8403 5433
rect 8376 5083 8383 5153
rect 8356 5076 8383 5083
rect 8316 4856 8323 4993
rect 8196 4247 8203 4353
rect 8236 4067 8243 4573
rect 8256 4487 8263 4753
rect 8276 4563 8283 4813
rect 8296 4707 8303 4823
rect 8336 4803 8343 4812
rect 8336 4796 8363 4803
rect 8356 4707 8363 4796
rect 8396 4763 8403 5193
rect 8416 4987 8423 5653
rect 8476 5596 8483 5733
rect 8496 5727 8503 5863
rect 8536 5787 8543 6053
rect 8556 5667 8563 6153
rect 8616 5607 8623 6616
rect 8636 5967 8643 6593
rect 8736 6416 8743 6773
rect 8756 6607 8763 7553
rect 8776 7347 8783 7873
rect 8796 7647 8803 7936
rect 8836 7627 8843 7873
rect 8876 7867 8883 8073
rect 8836 7456 8843 7493
rect 8856 7467 8863 7693
rect 8816 7403 8823 7412
rect 8816 7396 8843 7403
rect 8796 7087 8803 7143
rect 8816 7083 8823 7353
rect 8836 7267 8843 7396
rect 8807 7076 8823 7083
rect 8816 6948 8823 6973
rect 8856 6967 8863 7143
rect 8876 7087 8883 7853
rect 8896 7687 8903 8053
rect 8916 7988 8923 8113
rect 8916 7887 8923 7974
rect 9196 7976 9203 8013
rect 8996 7907 9003 7943
rect 9036 7927 9043 7943
rect 9036 7913 9053 7927
rect 9036 7867 9043 7913
rect 9027 7793 9033 7807
rect 8913 7680 8927 7693
rect 8916 7676 8923 7680
rect 8896 7387 8903 7454
rect 8853 6940 8867 6953
rect 8856 6936 8863 6940
rect 8896 6863 8903 7333
rect 8916 7107 8923 7613
rect 8996 7607 9003 7713
rect 8916 6887 8923 7072
rect 8896 6856 8923 6863
rect 8856 6636 8863 6833
rect 8836 6600 8843 6603
rect 8833 6587 8847 6600
rect 8836 6487 8843 6573
rect 8893 6567 8907 6573
rect 8813 6428 8827 6433
rect 8836 6386 8843 6433
rect 8867 6413 8873 6427
rect 8676 6116 8683 6373
rect 8716 6116 8723 6372
rect 8916 6347 8923 6856
rect 8936 6587 8943 7573
rect 9036 7547 9043 7673
rect 9056 7647 9063 7873
rect 8976 7407 8983 7493
rect 9076 7487 9083 7673
rect 9096 7587 9103 7973
rect 9216 7883 9223 7943
rect 9296 7927 9303 8213
rect 9216 7876 9243 7883
rect 9236 7707 9243 7876
rect 9316 7807 9323 8183
rect 9396 8127 9403 8193
rect 9416 8107 9423 8183
rect 9376 7988 9383 8093
rect 9456 8047 9463 8651
rect 9476 8507 9483 8913
rect 9516 8667 9523 8996
rect 9576 8686 9583 9093
rect 9636 8867 9643 9393
rect 9696 9107 9703 9203
rect 9716 9147 9723 9353
rect 9736 9327 9743 9503
rect 9776 9503 9783 9553
rect 9956 9536 9963 9573
rect 9856 9506 9863 9533
rect 9776 9496 9803 9503
rect 9753 9487 9767 9493
rect 9796 9467 9803 9496
rect 9976 9496 10003 9503
rect 9947 9475 9973 9482
rect 9996 9467 10003 9496
rect 10036 9327 10043 9534
rect 10076 9487 10083 9933
rect 10096 9747 10103 9913
rect 10336 9847 10343 10023
rect 10216 9756 10223 9813
rect 10436 9768 10443 10012
rect 10496 9927 10503 10054
rect 10656 10047 10663 10393
rect 10576 9987 10583 10023
rect 10696 9923 10703 10532
rect 10773 10527 10787 10540
rect 10716 9947 10723 10513
rect 10696 9916 10723 9923
rect 10473 9760 10487 9773
rect 10476 9756 10483 9760
rect 10196 9543 10203 9723
rect 10236 9687 10243 9723
rect 10236 9548 10243 9673
rect 10196 9536 10223 9543
rect 10093 9487 10107 9493
rect 10116 9407 10123 9534
rect 10216 9487 10223 9536
rect 9876 9236 9883 9273
rect 9916 9236 9923 9313
rect 9996 9207 10003 9234
rect 10036 9206 10043 9313
rect 10256 9248 10263 9633
rect 10380 9563 10393 9567
rect 10376 9553 10393 9563
rect 10376 9536 10383 9553
rect 10356 9500 10363 9503
rect 10353 9487 10367 9500
rect 10396 9407 10403 9503
rect 10316 9236 10323 9313
rect 9776 8927 9783 9003
rect 9896 8996 9903 9133
rect 9976 8996 10003 9003
rect 9936 8847 9943 8952
rect 9976 8887 9983 8996
rect 9533 8500 9547 8513
rect 9536 8496 9543 8500
rect 9576 8427 9583 8513
rect 9496 8327 9503 8393
rect 9476 8167 9483 8183
rect 9476 8067 9483 8153
rect 9413 7980 9427 7993
rect 9416 7976 9423 7980
rect 9336 7927 9343 7974
rect 9376 7947 9383 7974
rect 9436 7907 9443 7943
rect 9516 7887 9523 8373
rect 9596 8327 9603 8733
rect 9616 8707 9623 8833
rect 10036 8807 10043 9113
rect 10056 9008 10063 9153
rect 10096 8927 10103 9203
rect 10356 9147 10363 9203
rect 10356 9107 10363 9133
rect 10376 9083 10383 9353
rect 10356 9076 10383 9083
rect 10336 9006 10343 9053
rect 10356 8996 10363 9076
rect 10376 8956 10403 8963
rect 9633 8720 9647 8734
rect 9636 8716 9643 8720
rect 9676 8587 9683 8683
rect 9756 8607 9763 8653
rect 9776 8607 9783 8713
rect 9873 8700 9887 8713
rect 9876 8696 9883 8700
rect 10056 8647 10063 8703
rect 9753 8500 9767 8513
rect 9756 8496 9763 8500
rect 9956 8496 9963 8593
rect 9996 8508 10003 8533
rect 10116 8508 10123 8703
rect 9616 8307 9623 8493
rect 9816 8216 9823 8313
rect 9776 8180 9783 8183
rect 9756 8087 9763 8174
rect 9773 8167 9787 8180
rect 9576 7787 9583 7974
rect 9176 7587 9183 7643
rect 9107 7576 9123 7583
rect 9036 7420 9043 7423
rect 9033 7407 9047 7420
rect 8956 7307 8963 7373
rect 8956 6807 8963 7293
rect 9036 7267 9043 7393
rect 8976 6547 8983 7253
rect 9056 7156 9063 7233
rect 9116 7187 9123 7576
rect 9136 7168 9143 7473
rect 9176 7407 9183 7453
rect 9076 7067 9083 7123
rect 9116 7120 9123 7123
rect 9113 7107 9127 7120
rect 9076 6987 9083 7053
rect 9053 6940 9067 6953
rect 9096 6948 9103 7093
rect 9196 7063 9203 7632
rect 9216 7547 9223 7663
rect 9216 7426 9223 7533
rect 9256 7487 9263 7733
rect 9596 7703 9603 8013
rect 9696 7976 9703 8073
rect 9636 7923 9643 7943
rect 9636 7916 9663 7923
rect 9596 7696 9613 7703
rect 9656 7707 9663 7916
rect 9676 7907 9683 7943
rect 9276 7547 9283 7663
rect 9296 7523 9303 7654
rect 9316 7627 9323 7693
rect 9276 7516 9303 7523
rect 9276 7456 9283 7516
rect 9316 7456 9323 7513
rect 9256 7420 9263 7423
rect 9253 7407 9267 7420
rect 9396 7187 9403 7533
rect 9493 7460 9507 7473
rect 9496 7456 9503 7460
rect 9536 7456 9543 7553
rect 9516 7403 9523 7412
rect 9496 7396 9523 7403
rect 9496 7227 9503 7396
rect 9216 7087 9223 7132
rect 9256 7107 9263 7134
rect 9187 7056 9203 7063
rect 9056 6936 9063 6940
rect 9036 6887 9043 6903
rect 8996 6606 9003 6733
rect 9036 6707 9043 6873
rect 9116 6747 9123 6903
rect 9076 6567 9083 6603
rect 8973 6420 8987 6433
rect 8976 6416 8983 6420
rect 8756 6116 8763 6193
rect 8696 6007 8703 6083
rect 8736 6027 8743 6083
rect 8733 5908 8747 5913
rect 8676 5847 8683 5894
rect 8736 5603 8743 5713
rect 8753 5603 8767 5613
rect 8736 5600 8767 5603
rect 8736 5596 8763 5600
rect 8456 5560 8463 5563
rect 8453 5547 8467 5560
rect 8496 5507 8503 5563
rect 8560 5563 8573 5567
rect 8556 5556 8573 5563
rect 8560 5553 8573 5556
rect 8456 5376 8463 5473
rect 8536 5447 8543 5553
rect 8496 5376 8503 5413
rect 8476 5340 8483 5343
rect 8473 5327 8487 5340
rect 8516 5287 8523 5343
rect 8416 4787 8423 4893
rect 8436 4767 8443 5213
rect 8556 5207 8563 5513
rect 8553 5080 8567 5093
rect 8556 5076 8563 5080
rect 8596 5076 8603 5373
rect 8616 5287 8623 5553
rect 8636 5507 8643 5594
rect 8536 5027 8543 5043
rect 8396 4756 8423 4763
rect 8276 4556 8303 4563
rect 8333 4560 8347 4573
rect 8356 4567 8363 4693
rect 8336 4556 8343 4560
rect 8316 4503 8323 4523
rect 8316 4496 8343 4503
rect 8256 4336 8263 4373
rect 8276 4367 8283 4413
rect 8296 4227 8303 4303
rect 8213 4040 8227 4053
rect 8216 4036 8223 4040
rect 8256 4036 8263 4173
rect 8316 4007 8323 4473
rect 8336 4227 8343 4496
rect 8096 3796 8123 3803
rect 8176 3796 8203 3803
rect 8016 3743 8023 3793
rect 7996 3736 8023 3743
rect 7816 3276 7863 3283
rect 7876 3276 7883 3533
rect 7896 3367 7903 3633
rect 7736 3260 7743 3263
rect 7696 3203 7703 3253
rect 7733 3247 7747 3260
rect 7696 3196 7723 3203
rect 7696 2996 7703 3173
rect 7716 2867 7723 3196
rect 7776 3027 7783 3053
rect 7696 2647 7703 2763
rect 7796 2623 7803 3233
rect 7856 3207 7863 3276
rect 7816 2756 7823 3113
rect 7836 2767 7843 3193
rect 7876 2996 7883 3073
rect 7916 3007 7923 3553
rect 7976 3516 7983 3593
rect 7996 3567 8003 3736
rect 8096 3723 8103 3796
rect 8156 3756 8183 3763
rect 8096 3716 8123 3723
rect 7936 3487 7943 3514
rect 7996 3480 8003 3483
rect 7993 3467 8007 3480
rect 8096 3467 8103 3693
rect 8116 3647 8123 3716
rect 8056 3276 8083 3283
rect 8056 3127 8063 3253
rect 8076 3247 8083 3276
rect 8156 3223 8163 3733
rect 8176 3727 8183 3756
rect 8196 3523 8203 3796
rect 8176 3516 8203 3523
rect 8216 3516 8223 3813
rect 8256 3787 8263 3813
rect 8276 3667 8283 4003
rect 8336 3927 8343 4113
rect 8356 3947 8363 4513
rect 8327 3916 8343 3927
rect 8327 3913 8340 3916
rect 8376 3887 8383 4093
rect 8396 4048 8403 4353
rect 8416 4267 8423 4756
rect 8456 4587 8463 4973
rect 8436 4467 8443 4543
rect 8436 4167 8443 4373
rect 8456 4343 8463 4533
rect 8476 4367 8483 4913
rect 8536 4887 8543 5013
rect 8576 4927 8583 5043
rect 8627 5033 8633 5047
rect 8656 4947 8663 5133
rect 8696 5123 8703 5343
rect 8736 5287 8743 5343
rect 8776 5267 8783 5953
rect 8796 5866 8803 6133
rect 8816 5908 8823 6233
rect 8816 5667 8823 5894
rect 8836 5586 8843 6013
rect 8856 6007 8863 6173
rect 8896 6083 8903 6313
rect 8956 6287 8963 6383
rect 8953 6147 8967 6153
rect 8956 6116 8963 6133
rect 8996 6128 9003 6383
rect 9036 6167 9043 6473
rect 9056 6287 9063 6533
rect 9096 6187 9103 6593
rect 9116 6207 9123 6693
rect 9156 6607 9163 6934
rect 9176 6607 9183 7053
rect 9296 6936 9303 6993
rect 9336 6936 9343 6973
rect 9356 6900 9363 6903
rect 9353 6887 9367 6900
rect 9256 6507 9263 6603
rect 9356 6587 9363 6793
rect 9376 6687 9383 6892
rect 9396 6887 9403 6933
rect 9456 6907 9463 7013
rect 9476 6767 9483 6933
rect 9496 6807 9503 7213
rect 9556 7176 9563 7213
rect 9516 6947 9523 7143
rect 9596 7027 9603 7613
rect 9616 7307 9623 7493
rect 9656 7107 9663 7693
rect 9676 7667 9683 7793
rect 9676 7527 9683 7613
rect 9696 7503 9703 7873
rect 9736 7607 9743 7693
rect 9756 7547 9763 8052
rect 9796 7883 9803 8073
rect 9856 8027 9863 8313
rect 9876 8087 9883 8452
rect 9896 8387 9903 8494
rect 9896 8087 9903 8213
rect 9956 8167 9963 8313
rect 9916 8067 9923 8133
rect 9893 7980 9907 7993
rect 9896 7976 9903 7980
rect 9776 7876 9803 7883
rect 9776 7627 9783 7876
rect 9816 7727 9823 7974
rect 9813 7707 9827 7713
rect 9876 7703 9883 7943
rect 9936 7847 9943 7993
rect 9956 7927 9963 7993
rect 9976 7767 9983 8293
rect 9996 8207 10003 8433
rect 10016 8307 10023 8463
rect 10116 8447 10123 8494
rect 10016 8196 10023 8233
rect 10136 8147 10143 8833
rect 10236 8547 10243 8593
rect 10236 8496 10243 8533
rect 10276 8467 10283 8714
rect 10296 8687 10303 8833
rect 10376 8827 10383 8956
rect 10376 8748 10383 8813
rect 10436 8787 10443 9153
rect 10456 8847 10463 9593
rect 10476 8986 10483 9533
rect 10516 9503 10523 9753
rect 10616 9723 10623 9813
rect 10656 9756 10663 9913
rect 10616 9716 10643 9723
rect 10607 9553 10613 9567
rect 10636 9543 10643 9716
rect 10676 9703 10683 9712
rect 10616 9536 10643 9543
rect 10656 9696 10683 9703
rect 10496 9496 10523 9503
rect 10556 9500 10563 9503
rect 10496 9248 10503 9496
rect 10553 9487 10567 9500
rect 10516 9167 10523 9473
rect 10656 9203 10663 9696
rect 10716 9647 10723 9916
rect 10736 9607 10743 10493
rect 10776 10276 10783 10353
rect 10816 10276 10823 10393
rect 10796 10083 10803 10243
rect 10776 10080 10803 10083
rect 10773 10076 10803 10080
rect 10756 9787 10763 10073
rect 10773 10067 10787 10076
rect 10813 10060 10827 10073
rect 10816 10056 10823 10060
rect 10856 10056 10863 10393
rect 10896 9967 10903 10733
rect 10916 10546 10923 10573
rect 10916 10026 10923 10273
rect 10756 9726 10763 9773
rect 10816 9536 10823 9953
rect 10916 9756 10923 9813
rect 10936 9763 10943 10613
rect 10956 10588 10963 10793
rect 11076 10766 11083 10793
rect 11036 10760 11043 10763
rect 10993 10747 11007 10752
rect 11033 10747 11047 10760
rect 11236 10707 11243 10763
rect 11036 10576 11043 10613
rect 10956 10026 10963 10433
rect 10976 9768 10983 10053
rect 10936 9756 10963 9763
rect 10856 9647 10863 9723
rect 10853 9540 10867 9553
rect 10856 9536 10863 9540
rect 10796 9467 10803 9503
rect 10636 9196 10663 9203
rect 10676 9127 10683 9223
rect 10716 9127 10723 9413
rect 10956 9367 10963 9756
rect 10976 9607 10983 9754
rect 10996 9726 11003 10133
rect 11036 10107 11043 10193
rect 11036 10056 11043 10093
rect 11056 9987 11063 10023
rect 11136 9967 11143 10532
rect 11056 9536 11063 9952
rect 11156 9827 11163 10573
rect 11256 10507 11263 10543
rect 11176 10276 11203 10283
rect 11176 9983 11183 10276
rect 11296 10236 11323 10243
rect 11256 10147 11263 10203
rect 11316 10103 11323 10236
rect 11307 10096 11323 10103
rect 11296 10056 11303 10093
rect 11176 9976 11193 9983
rect 11196 9763 11203 9973
rect 11176 9756 11203 9763
rect 11116 9506 11123 9683
rect 11036 9427 11043 9503
rect 10736 9187 10743 9223
rect 10636 9016 10643 9053
rect 10696 8986 10703 9033
rect 10376 8683 10383 8734
rect 10356 8676 10383 8683
rect 10396 8667 10403 8703
rect 10456 8647 10463 8703
rect 10636 8696 10643 8833
rect 10776 8743 10783 9254
rect 10916 9216 10923 9353
rect 11076 9347 11083 9503
rect 10853 9020 10867 9033
rect 11016 9028 11023 9333
rect 11036 9220 11043 9223
rect 11033 9207 11047 9220
rect 10856 9016 10863 9020
rect 10836 8907 10843 8983
rect 11016 8986 11023 9014
rect 10776 8736 10793 8743
rect 10456 8587 10463 8633
rect 10453 8500 10467 8513
rect 10456 8496 10463 8500
rect 10176 8207 10183 8393
rect 10176 8147 10183 8193
rect 10016 7887 10023 8093
rect 10056 8087 10063 8133
rect 10076 8107 10083 8131
rect 10196 8107 10203 8153
rect 10076 7976 10083 8053
rect 9813 7680 9827 7693
rect 9856 7696 9883 7703
rect 9816 7676 9823 7680
rect 9856 7676 9863 7696
rect 9836 7640 9843 7643
rect 9833 7627 9847 7640
rect 9876 7607 9883 7643
rect 9996 7607 10003 7833
rect 10096 7807 10103 7943
rect 10136 7940 10143 7943
rect 10133 7927 10147 7940
rect 10016 7667 10023 7793
rect 10076 7676 10083 7713
rect 10113 7680 10127 7693
rect 10116 7676 10123 7680
rect 9676 7496 9703 7503
rect 9636 6903 9643 7093
rect 9676 7083 9683 7496
rect 9713 7487 9727 7493
rect 9796 7456 9803 7493
rect 9696 7426 9703 7453
rect 9856 7447 9863 7593
rect 10056 7587 10063 7643
rect 10096 7587 10103 7643
rect 10156 7643 10163 7933
rect 10196 7807 10203 7873
rect 10216 7727 10223 8173
rect 10236 7956 10243 8233
rect 10296 8196 10303 8433
rect 10336 8343 10343 8494
rect 10536 8483 10543 8573
rect 10576 8487 10583 8513
rect 10536 8476 10563 8483
rect 10336 8336 10363 8343
rect 10276 8160 10283 8163
rect 10273 8147 10287 8160
rect 10316 8067 10323 8163
rect 10356 8067 10363 8336
rect 10376 8087 10383 8453
rect 10396 8307 10403 8463
rect 10436 8460 10443 8463
rect 10433 8447 10447 8460
rect 10476 8407 10483 8453
rect 10516 8196 10523 8233
rect 10536 8227 10543 8476
rect 10596 8327 10603 8493
rect 10736 8480 10743 8483
rect 10733 8467 10747 8480
rect 10836 8367 10843 8872
rect 10856 8587 10863 8703
rect 10916 8647 10923 8703
rect 10853 8480 10867 8493
rect 10856 8476 10863 8480
rect 10876 8436 10903 8443
rect 10576 8166 10583 8213
rect 10496 8067 10503 8163
rect 10276 7807 10283 7953
rect 10416 7847 10423 7963
rect 10147 7636 10163 7643
rect 9896 7467 9903 7553
rect 9876 7436 9903 7443
rect 9596 6896 9643 6903
rect 9656 7076 9683 7083
rect 9656 6887 9663 7076
rect 9576 6807 9583 6833
rect 9527 6753 9533 6767
rect 9213 6420 9227 6433
rect 9216 6416 9223 6420
rect 9236 6247 9243 6383
rect 9356 6327 9363 6573
rect 9376 6387 9383 6673
rect 9476 6636 9483 6693
rect 9456 6600 9463 6603
rect 9453 6587 9467 6600
rect 9456 6527 9463 6573
rect 9496 6567 9503 6603
rect 9416 6416 9423 6453
rect 9453 6420 9467 6433
rect 9456 6416 9463 6420
rect 8896 6076 8943 6083
rect 8856 5787 8863 5993
rect 8876 5827 8883 5953
rect 8896 5627 8903 6033
rect 8916 5927 8923 6076
rect 8976 5967 8983 6083
rect 8996 5943 9003 6053
rect 9096 6047 9103 6103
rect 9116 6067 9123 6094
rect 9136 5987 9143 6233
rect 9256 6207 9263 6293
rect 9416 6287 9423 6313
rect 9436 6267 9443 6372
rect 9476 6148 9483 6233
rect 9376 6047 9383 6093
rect 8976 5936 9003 5943
rect 8976 5896 8983 5936
rect 9056 5887 9063 5913
rect 9076 5876 9103 5883
rect 8996 5827 9003 5863
rect 9096 5727 9103 5876
rect 9376 5876 9383 6033
rect 9196 5628 9203 5832
rect 9227 5713 9233 5727
rect 8676 5116 8703 5123
rect 8676 5027 8683 5116
rect 8533 4860 8547 4873
rect 8696 4867 8703 5074
rect 8716 5027 8723 5253
rect 8816 5107 8823 5533
rect 8836 5388 8843 5572
rect 8856 5547 8863 5583
rect 8896 5547 8903 5613
rect 9236 5587 9243 5713
rect 8856 5347 8863 5533
rect 8876 5247 8883 5453
rect 8956 5376 8963 5433
rect 9136 5376 9143 5553
rect 9176 5376 9183 5433
rect 8936 5340 8943 5343
rect 8933 5327 8947 5340
rect 9156 5340 9163 5343
rect 9196 5340 9203 5343
rect 8816 5076 8863 5083
rect 8856 5047 8863 5076
rect 8747 5043 8760 5047
rect 8747 5036 8763 5043
rect 8747 5033 8760 5036
rect 8796 5007 8803 5043
rect 8536 4856 8543 4860
rect 8496 4827 8503 4854
rect 8716 4856 8723 4973
rect 8496 4727 8503 4813
rect 8693 4803 8707 4813
rect 8693 4800 8723 4803
rect 8696 4796 8723 4800
rect 8716 4507 8723 4796
rect 8736 4787 8743 4823
rect 8776 4576 8783 4773
rect 8516 4407 8523 4433
rect 8536 4367 8543 4413
rect 8556 4387 8563 4433
rect 8456 4336 8483 4343
rect 8496 4127 8503 4292
rect 8513 4040 8527 4053
rect 8516 4036 8523 4040
rect 8256 3516 8263 3573
rect 8296 3547 8303 3853
rect 8336 3816 8343 3873
rect 8396 3867 8403 4034
rect 8456 4000 8463 4003
rect 8453 3987 8467 4000
rect 8413 3820 8427 3833
rect 8416 3816 8423 3820
rect 8456 3787 8463 3933
rect 8176 3327 8183 3516
rect 8236 3447 8243 3483
rect 8216 3407 8223 3433
rect 8220 3243 8233 3247
rect 8216 3233 8233 3243
rect 8156 3216 8183 3223
rect 7896 2746 7903 2793
rect 7867 2720 7883 2723
rect 7867 2716 7887 2720
rect 7873 2707 7887 2716
rect 7776 2616 7803 2623
rect 7536 2347 7543 2474
rect 7633 2480 7647 2493
rect 7696 2487 7703 2533
rect 7636 2476 7643 2480
rect 7696 2446 7703 2473
rect 7536 2247 7543 2333
rect 7576 2187 7583 2443
rect 7616 2407 7623 2443
rect 7636 2256 7643 2293
rect 7576 1956 7603 1963
rect 7576 1867 7583 1956
rect 7656 1923 7663 2153
rect 7676 2047 7683 2223
rect 7636 1916 7663 1923
rect 7576 1736 7583 1773
rect 7656 1747 7663 1893
rect 7716 1767 7723 2093
rect 7736 1827 7743 2593
rect 7756 2247 7763 2613
rect 7776 2227 7783 2616
rect 7856 2487 7863 2673
rect 7916 2527 7923 2753
rect 7936 2547 7943 2833
rect 7956 2647 7963 2773
rect 7876 2460 7883 2463
rect 7873 2447 7887 2460
rect 7876 2256 7883 2293
rect 7896 2263 7903 2453
rect 7916 2327 7923 2513
rect 7936 2327 7943 2463
rect 7956 2407 7963 2454
rect 7896 2256 7913 2263
rect 7836 1956 7843 2053
rect 7916 1927 7923 2254
rect 7816 1827 7823 1923
rect 7856 1827 7863 1923
rect 7936 1907 7943 2073
rect 7956 2007 7963 2313
rect 7976 1807 7983 2993
rect 8016 2687 8023 2994
rect 8036 2967 8043 3033
rect 8076 2907 8083 2963
rect 8116 2960 8123 2963
rect 8113 2947 8127 2960
rect 8116 2788 8123 2893
rect 8156 2607 8163 2774
rect 8176 2687 8183 3216
rect 8196 2947 8203 3233
rect 8196 2827 8203 2853
rect 8216 2847 8223 3233
rect 8256 2863 8263 3313
rect 8276 3087 8283 3353
rect 8236 2856 8263 2863
rect 8196 2647 8203 2792
rect 8216 2427 8223 2673
rect 8236 2567 8243 2856
rect 8256 2707 8263 2833
rect 8276 2788 8283 3073
rect 8296 3007 8303 3333
rect 8316 3247 8323 3713
rect 8356 3227 8363 3772
rect 8396 3747 8403 3783
rect 8316 2996 8323 3193
rect 8376 3087 8383 3653
rect 8476 3587 8483 3813
rect 8496 3607 8503 4003
rect 8516 3747 8523 3893
rect 8536 3786 8543 3853
rect 8436 3516 8443 3553
rect 8476 3516 8483 3573
rect 8536 3567 8543 3772
rect 8556 3547 8563 4373
rect 8716 4336 8723 4453
rect 8636 4307 8643 4334
rect 8776 4307 8783 4493
rect 8816 4307 8823 5013
rect 8836 4427 8843 4633
rect 8856 4387 8863 4813
rect 8696 4227 8703 4303
rect 8596 4087 8603 4193
rect 8576 3783 8583 3833
rect 8616 3828 8623 4053
rect 8636 3907 8643 4213
rect 8656 3887 8663 4153
rect 8716 4036 8723 4093
rect 8736 4067 8743 4292
rect 8796 4006 8803 4213
rect 8816 3867 8823 4034
rect 8856 3927 8863 4034
rect 8876 4007 8883 4853
rect 8896 4807 8903 5173
rect 8916 4867 8923 5093
rect 9036 5088 9043 5193
rect 8956 5027 8963 5074
rect 9116 5063 9123 5333
rect 9153 5327 9167 5340
rect 9193 5327 9207 5340
rect 9236 5327 9243 5513
rect 9256 5287 9263 5614
rect 9316 5307 9323 5713
rect 9336 5567 9343 5872
rect 9396 5727 9403 6103
rect 9436 5876 9443 5973
rect 9476 5847 9483 6134
rect 9387 5716 9403 5727
rect 9387 5713 9400 5716
rect 9356 5527 9363 5653
rect 9496 5627 9503 6353
rect 9516 5747 9523 6593
rect 9536 6447 9543 6613
rect 9556 6247 9563 6733
rect 9536 5887 9543 6173
rect 9576 6087 9583 6453
rect 9453 5600 9467 5613
rect 9456 5596 9463 5600
rect 9496 5566 9503 5613
rect 9416 5487 9423 5533
rect 9436 5527 9443 5563
rect 9416 5376 9423 5473
rect 9516 5447 9523 5733
rect 9576 5527 9583 5973
rect 9596 5727 9603 6873
rect 9616 6467 9623 6633
rect 9636 6423 9643 6693
rect 9676 6648 9683 6934
rect 9696 6667 9703 7353
rect 9736 7287 9743 7423
rect 9776 7267 9783 7423
rect 9796 7267 9803 7313
rect 9856 7287 9863 7333
rect 9776 7187 9783 7253
rect 9736 7120 9743 7123
rect 9776 7120 9783 7123
rect 9733 7107 9747 7120
rect 9773 7107 9787 7120
rect 9716 6707 9723 7093
rect 9736 7067 9743 7093
rect 9816 6987 9823 7213
rect 9776 6936 9783 6973
rect 9856 6927 9863 7173
rect 9876 6947 9883 7373
rect 9896 7287 9903 7436
rect 9987 7443 10000 7447
rect 9987 7436 10003 7443
rect 9987 7433 10000 7436
rect 10136 7387 10143 7632
rect 10196 7607 10203 7713
rect 10216 7463 10223 7533
rect 10256 7487 10263 7693
rect 10316 7676 10323 7793
rect 10353 7680 10367 7693
rect 10356 7676 10363 7680
rect 10296 7587 10303 7643
rect 10296 7467 10303 7513
rect 10173 7440 10187 7453
rect 10196 7456 10223 7463
rect 10176 7436 10183 7440
rect 10196 7307 10203 7456
rect 10236 7436 10263 7443
rect 10256 7387 10263 7436
rect 10256 7347 10263 7373
rect 9900 7266 9920 7267
rect 9907 7253 9913 7266
rect 9916 7107 9923 7173
rect 9933 7167 9947 7173
rect 9953 7160 9967 7173
rect 9993 7160 10007 7173
rect 10036 7167 10043 7213
rect 9956 7156 9963 7160
rect 9996 7156 10003 7160
rect 10096 7143 10103 7293
rect 10376 7283 10383 7533
rect 10396 7367 10403 7673
rect 10456 7567 10463 7693
rect 10476 7647 10483 7793
rect 10516 7683 10523 8133
rect 10596 8027 10603 8273
rect 10636 8263 10643 8313
rect 10696 8287 10703 8353
rect 10616 8256 10643 8263
rect 10556 7967 10563 8013
rect 10560 7703 10573 7707
rect 10496 7676 10523 7683
rect 10556 7693 10573 7703
rect 10556 7676 10563 7693
rect 10596 7687 10603 7813
rect 10616 7687 10623 8256
rect 10636 7867 10643 8233
rect 10656 7967 10663 8273
rect 10676 8127 10683 8213
rect 10713 8208 10727 8213
rect 10756 8196 10763 8273
rect 10796 8196 10803 8253
rect 10876 8247 10883 8436
rect 10936 8363 10943 8694
rect 10916 8356 10943 8363
rect 10496 7547 10503 7676
rect 10536 7587 10543 7643
rect 10536 7487 10543 7573
rect 10576 7567 10583 7643
rect 10616 7627 10623 7652
rect 10556 7556 10573 7563
rect 10453 7460 10467 7473
rect 10456 7456 10463 7460
rect 10376 7276 10403 7283
rect 10156 7143 10163 7193
rect 9976 7027 9983 7123
rect 10056 7087 10063 7143
rect 10096 7136 10123 7143
rect 10136 7136 10163 7143
rect 10296 7136 10303 7213
rect 10136 6987 10143 7136
rect 9876 6916 9903 6923
rect 9756 6847 9763 6903
rect 9756 6683 9763 6833
rect 9756 6676 9783 6683
rect 9716 6636 9723 6672
rect 9656 6527 9663 6592
rect 9696 6567 9703 6603
rect 9616 6416 9663 6423
rect 9616 6367 9623 6416
rect 9716 6427 9723 6473
rect 9676 6367 9683 6383
rect 9676 6356 9693 6367
rect 9680 6353 9693 6356
rect 9636 6116 9643 6153
rect 9673 6120 9687 6133
rect 9716 6127 9723 6153
rect 9676 6116 9683 6120
rect 9736 6087 9743 6333
rect 9613 6067 9627 6072
rect 9713 6063 9727 6073
rect 9696 6060 9727 6063
rect 9693 6056 9723 6060
rect 9693 6047 9707 6056
rect 9706 6040 9707 6047
rect 9656 5896 9663 6033
rect 9713 6023 9727 6033
rect 9696 6020 9727 6023
rect 9696 6016 9723 6020
rect 9676 5947 9683 6013
rect 9696 5927 9703 6016
rect 9636 5827 9643 5863
rect 9596 5547 9603 5673
rect 9636 5667 9643 5813
rect 9676 5527 9683 5563
rect 9716 5527 9723 5653
rect 9756 5463 9763 6653
rect 9776 6327 9783 6676
rect 9796 6648 9803 6903
rect 9816 6607 9823 6813
rect 9836 6747 9843 6883
rect 9856 6667 9863 6873
rect 9896 6823 9903 6916
rect 9876 6816 9903 6823
rect 9876 6767 9883 6816
rect 9913 6667 9927 6673
rect 9827 6596 9843 6603
rect 9796 6427 9803 6473
rect 9816 6327 9823 6413
rect 9776 6287 9783 6313
rect 9776 5876 9783 6093
rect 9756 5456 9783 5463
rect 9376 5247 9383 5343
rect 9536 5327 9543 5413
rect 9116 5056 9143 5063
rect 8973 5027 8987 5033
rect 9136 5027 9143 5056
rect 8993 4840 9007 4853
rect 8996 4836 9003 4840
rect 8956 4807 8963 4823
rect 8956 4703 8963 4793
rect 9036 4783 9043 4913
rect 9036 4776 9063 4783
rect 8956 4696 8983 4703
rect 8896 4507 8903 4673
rect 8936 4547 8943 4673
rect 8976 4667 8983 4696
rect 8996 4556 9003 4593
rect 8936 4336 8943 4393
rect 8976 4348 8983 4523
rect 9016 4447 9023 4523
rect 8876 3816 8883 3972
rect 8576 3776 8603 3783
rect 8596 3543 8603 3776
rect 8816 3747 8823 3772
rect 8836 3727 8843 3783
rect 8836 3647 8843 3713
rect 8596 3536 8623 3543
rect 8556 3503 8563 3533
rect 8556 3496 8583 3503
rect 8456 3480 8463 3483
rect 8453 3467 8467 3480
rect 8496 3367 8503 3393
rect 8416 3296 8423 3333
rect 8453 3300 8467 3313
rect 8456 3296 8463 3300
rect 8516 3288 8523 3413
rect 8556 3327 8563 3393
rect 8576 3283 8583 3496
rect 8596 3287 8603 3494
rect 8556 3276 8583 3283
rect 8416 3067 8423 3233
rect 8436 3187 8443 3263
rect 8356 2996 8363 3053
rect 8456 2983 8463 3113
rect 8456 2976 8483 2983
rect 8356 2887 8363 2913
rect 8456 2867 8463 2953
rect 8293 2780 8307 2793
rect 8296 2776 8303 2780
rect 8336 2776 8343 2853
rect 8476 2847 8483 2976
rect 8516 2883 8523 3213
rect 8556 3127 8563 3276
rect 8616 3127 8623 3536
rect 8856 3327 8863 3693
rect 8896 3547 8903 4233
rect 8916 4227 8923 4303
rect 8956 4063 8963 4193
rect 8976 4187 8983 4334
rect 8956 4056 8983 4063
rect 8976 4048 8983 4056
rect 8916 3707 8923 3993
rect 8936 3747 8943 3853
rect 8916 3536 8923 3633
rect 8760 3283 8773 3287
rect 8756 3276 8773 3283
rect 8760 3273 8773 3276
rect 8856 3276 8883 3283
rect 8756 2887 8763 3253
rect 8856 3127 8863 3276
rect 8956 3267 8963 3533
rect 8976 3527 8983 3893
rect 8973 3447 8987 3453
rect 8976 3243 8983 3313
rect 8996 3247 9003 3993
rect 9016 3607 9023 3673
rect 9016 3467 9023 3572
rect 8916 3236 8943 3243
rect 8816 3016 8823 3053
rect 8856 2987 8863 3113
rect 8896 2907 8903 3233
rect 8916 2887 8923 3113
rect 8936 3107 8943 3236
rect 8956 3236 8983 3243
rect 8956 3167 8963 3236
rect 8980 3203 8993 3207
rect 8976 3200 8993 3203
rect 8973 3193 8993 3200
rect 8973 3187 8987 3193
rect 8496 2876 8523 2883
rect 8456 2787 8463 2813
rect 8256 2667 8263 2693
rect 8256 2503 8263 2653
rect 8316 2567 8323 2732
rect 8356 2687 8363 2743
rect 8256 2496 8283 2503
rect 7996 2327 8003 2353
rect 8000 2306 8013 2307
rect 8007 2293 8013 2306
rect 7996 2187 8003 2253
rect 8016 2227 8023 2272
rect 8036 2267 8043 2313
rect 8053 2260 8067 2273
rect 8056 2256 8063 2260
rect 8096 2256 8103 2313
rect 8176 2236 8183 2293
rect 8236 2236 8243 2333
rect 8256 2247 8263 2373
rect 8076 2027 8083 2223
rect 8053 1960 8067 1973
rect 8056 1956 8063 1960
rect 8096 1956 8103 1993
rect 8036 1920 8043 1923
rect 8033 1907 8047 1920
rect 7956 1796 7973 1803
rect 7516 1507 7523 1734
rect 7696 1716 7723 1723
rect 7556 1607 7563 1653
rect 7656 1647 7663 1683
rect 7576 1487 7583 1633
rect 7716 1567 7723 1716
rect 7496 1407 7503 1453
rect 7796 1448 7803 1553
rect 7876 1436 7883 1493
rect 7456 1216 7503 1223
rect 7496 1186 7503 1216
rect 7196 327 7203 393
rect 7236 188 7243 753
rect 7296 696 7303 793
rect 7316 767 7323 933
rect 7456 916 7463 1033
rect 7436 827 7443 883
rect 7316 487 7323 663
rect 7356 660 7363 663
rect 7353 647 7367 660
rect 7436 627 7443 813
rect 7516 727 7523 1153
rect 7536 886 7543 913
rect 7556 696 7563 1073
rect 7636 923 7643 1172
rect 7636 916 7663 923
rect 7696 916 7703 973
rect 7456 627 7463 694
rect 7576 527 7583 663
rect 7356 487 7363 513
rect 7536 396 7543 493
rect 7396 366 7403 393
rect 7616 367 7623 513
rect 7316 227 7323 363
rect 7356 327 7363 363
rect 7676 366 7683 872
rect 7756 567 7763 1434
rect 7776 767 7783 1053
rect 7796 987 7803 1434
rect 7956 1406 7963 1796
rect 7996 1716 8003 1833
rect 8056 1716 8063 1753
rect 8076 1468 8083 1923
rect 8116 1867 8123 1893
rect 8136 1687 8143 2013
rect 8156 1627 8163 1933
rect 7856 1327 7863 1403
rect 8016 1367 8023 1433
rect 7816 1183 7823 1253
rect 7876 1216 7903 1223
rect 7816 1176 7843 1183
rect 7816 887 7823 1013
rect 7876 928 7883 993
rect 7896 967 7903 1216
rect 7956 963 7963 1213
rect 7956 956 7983 963
rect 7913 920 7927 933
rect 7916 916 7923 920
rect 7956 887 7963 933
rect 7856 827 7863 883
rect 7856 727 7863 813
rect 7896 807 7903 883
rect 7976 867 7983 956
rect 7896 696 7903 753
rect 7796 627 7803 663
rect 7856 660 7863 663
rect 7853 647 7867 660
rect 7816 366 7823 433
rect 7676 327 7683 352
rect 7316 187 7323 213
rect 7436 176 7443 253
rect 7856 188 7863 313
rect 7896 188 7903 553
rect 7916 367 7923 653
rect 7936 647 7943 793
rect 7996 787 8003 1213
rect 8016 1186 8023 1353
rect 8036 1228 8043 1453
rect 8116 1448 8123 1473
rect 8096 1287 8103 1403
rect 8133 1387 8147 1392
rect 8056 1216 8063 1273
rect 8036 807 8043 953
rect 8076 923 8083 1183
rect 8136 1107 8143 1333
rect 8056 916 8103 923
rect 8136 916 8143 953
rect 7956 667 7963 713
rect 7936 487 7943 553
rect 7956 507 7963 593
rect 7956 396 7963 493
rect 7996 447 8003 773
rect 8056 666 8063 916
rect 8156 847 8163 873
rect 8176 727 8183 2113
rect 8216 2027 8223 2233
rect 8276 2127 8283 2413
rect 8316 2347 8323 2532
rect 8336 2387 8343 2553
rect 8356 2507 8363 2673
rect 8436 2347 8443 2553
rect 8476 2547 8483 2833
rect 8496 2747 8503 2876
rect 8536 2776 8543 2873
rect 8576 2776 8583 2873
rect 8616 2776 8623 2813
rect 8696 2756 8723 2763
rect 8556 2687 8563 2732
rect 8476 2476 8483 2512
rect 8520 2483 8533 2487
rect 8516 2476 8533 2483
rect 8520 2473 8533 2476
rect 8556 2467 8563 2593
rect 8556 2443 8563 2453
rect 8576 2447 8583 2473
rect 8496 2387 8503 2443
rect 8536 2436 8563 2443
rect 8416 2187 8423 2243
rect 8516 2147 8523 2413
rect 8536 2236 8543 2436
rect 8596 2427 8603 2743
rect 8656 2667 8663 2723
rect 8556 2067 8563 2113
rect 8216 1987 8223 2013
rect 8216 1748 8223 1973
rect 8236 1926 8243 1993
rect 8496 1956 8503 2013
rect 8576 2007 8583 2033
rect 8516 1867 8523 1923
rect 8556 1887 8563 1973
rect 8527 1856 8543 1863
rect 8296 1736 8303 1853
rect 8536 1736 8543 1856
rect 8196 827 8203 1613
rect 8216 967 8223 1593
rect 8276 1567 8283 1703
rect 8236 1187 8243 1473
rect 8376 1436 8403 1443
rect 8336 1400 8343 1403
rect 8276 1287 8283 1392
rect 8333 1387 8347 1400
rect 8396 1287 8403 1436
rect 8276 1216 8283 1273
rect 8396 1167 8403 1273
rect 8376 916 8383 1013
rect 8316 880 8323 883
rect 8313 867 8327 880
rect 7916 227 7923 293
rect 7456 67 7463 143
rect 7516 27 7523 174
rect 7936 147 7943 233
rect 7676 27 7683 143
rect 7836 47 7843 133
rect 8036 107 8043 613
rect 8056 547 8063 652
rect 8073 547 8087 553
rect 8096 247 8103 593
rect 8116 366 8123 433
rect 8116 267 8123 352
rect 8136 307 8143 663
rect 8176 607 8183 673
rect 8176 423 8183 493
rect 8196 447 8203 813
rect 8313 700 8327 713
rect 8316 696 8323 700
rect 8416 707 8423 1673
rect 8476 1527 8483 1703
rect 8576 1667 8583 1773
rect 8416 666 8423 693
rect 8436 687 8443 1513
rect 8553 1440 8567 1453
rect 8556 1436 8563 1440
rect 8596 1436 8603 1733
rect 8616 1607 8623 2474
rect 8636 2167 8643 2553
rect 8656 2206 8663 2653
rect 8716 2607 8723 2756
rect 8747 2593 8753 2607
rect 8796 2507 8803 2533
rect 8733 2480 8747 2493
rect 8736 2476 8743 2480
rect 8716 2440 8723 2443
rect 8656 2067 8663 2192
rect 8676 2027 8683 2433
rect 8713 2427 8727 2440
rect 8696 2127 8703 2273
rect 8636 1567 8643 2013
rect 8736 1956 8743 2313
rect 8776 2256 8783 2493
rect 8796 2287 8803 2493
rect 8816 2407 8823 2763
rect 8876 2227 8883 2613
rect 8916 2476 8923 2573
rect 8956 2508 8963 3132
rect 9016 3067 9023 3432
rect 9036 3187 9043 4253
rect 9056 4007 9063 4776
rect 9096 4407 9103 5013
rect 9176 5007 9183 5054
rect 9416 4927 9423 5293
rect 9476 5287 9483 5323
rect 9616 5303 9623 5353
rect 9636 5327 9643 5363
rect 9616 5296 9643 5303
rect 9476 5108 9483 5273
rect 9636 5207 9643 5296
rect 9516 5067 9523 5193
rect 9656 5043 9663 5233
rect 9713 5080 9727 5094
rect 9716 5076 9723 5080
rect 9656 5036 9683 5043
rect 9236 4707 9243 4843
rect 9336 4836 9363 4843
rect 9136 4526 9143 4653
rect 9196 4556 9203 4693
rect 9276 4527 9283 4693
rect 9336 4687 9343 4836
rect 9396 4767 9403 4803
rect 9396 4567 9403 4753
rect 9436 4583 9443 4873
rect 9456 4807 9463 4834
rect 9476 4827 9483 4933
rect 9656 4863 9663 5036
rect 9636 4856 9663 4863
rect 9596 4767 9603 4823
rect 9416 4576 9443 4583
rect 9116 4336 9123 4373
rect 9156 3927 9163 4003
rect 9196 3967 9203 4003
rect 9176 3816 9183 3873
rect 9076 3707 9083 3783
rect 9096 3683 9103 3753
rect 9076 3676 9103 3683
rect 9056 3507 9063 3633
rect 9056 3247 9063 3393
rect 9076 3247 9083 3676
rect 9093 3527 9107 3533
rect 9136 3516 9143 3733
rect 9196 3536 9203 3773
rect 9236 3567 9243 4433
rect 9256 3707 9263 4034
rect 9276 4007 9283 4073
rect 9276 3767 9283 3813
rect 9296 3767 9303 4554
rect 9416 4556 9423 4576
rect 9456 4556 9463 4593
rect 9316 3787 9323 4553
rect 9436 4487 9443 4523
rect 9336 4247 9343 4303
rect 9336 4007 9343 4233
rect 9416 4227 9423 4373
rect 9476 4348 9483 4373
rect 9396 4036 9403 4073
rect 9416 3887 9423 4003
rect 9476 3867 9483 4334
rect 9516 4307 9523 4653
rect 9556 4336 9563 4433
rect 9596 4407 9603 4593
rect 9616 4527 9623 4713
rect 9656 4607 9663 4856
rect 9696 4556 9703 4673
rect 9776 4583 9783 5456
rect 9796 5387 9803 5773
rect 9816 5767 9823 6133
rect 9836 6127 9843 6596
rect 9856 6427 9863 6653
rect 9913 6640 9927 6653
rect 9916 6636 9923 6640
rect 10016 6607 10023 6653
rect 10036 6606 10043 6793
rect 10136 6747 10143 6973
rect 10176 6916 10183 6953
rect 10256 6807 10263 7013
rect 10276 6867 10283 6953
rect 10296 6847 10303 6913
rect 10316 6827 10323 7013
rect 10396 6987 10403 7276
rect 10436 7187 10443 7423
rect 10476 7416 10503 7423
rect 10496 7387 10503 7416
rect 10453 7180 10467 7193
rect 10456 7176 10463 7180
rect 10416 7087 10423 7143
rect 10156 6636 10163 6773
rect 10276 6668 10283 6733
rect 10193 6640 10207 6653
rect 10196 6636 10203 6640
rect 9896 6416 9903 6453
rect 9976 6396 9983 6473
rect 9876 6380 9883 6383
rect 9916 6380 9923 6383
rect 9873 6367 9887 6380
rect 9913 6367 9927 6380
rect 9856 6116 9863 6173
rect 9896 6167 9903 6313
rect 9896 6116 9903 6153
rect 9876 6063 9883 6083
rect 9933 6063 9947 6073
rect 9876 6060 9947 6063
rect 9876 6056 9943 6060
rect 9976 6047 9983 6133
rect 10016 6047 10023 6453
rect 10036 6396 10043 6553
rect 10076 6207 10083 6613
rect 10176 6547 10183 6603
rect 10276 6547 10283 6614
rect 10296 6547 10303 6623
rect 10336 6423 10343 6973
rect 10436 6967 10443 7133
rect 10496 7127 10503 7373
rect 10556 7143 10563 7556
rect 10636 7487 10643 7674
rect 10656 7456 10663 7913
rect 10676 7607 10683 8113
rect 10696 8107 10703 8152
rect 10776 8107 10783 8163
rect 10856 8087 10863 8173
rect 10696 7827 10703 8013
rect 10696 7646 10703 7753
rect 10716 7687 10723 8073
rect 10876 8047 10883 8233
rect 10916 8227 10923 8356
rect 10956 8323 10963 8973
rect 11076 8980 11083 8983
rect 11073 8967 11087 8980
rect 11116 8887 11123 8983
rect 11156 8967 11163 9493
rect 11176 8847 11183 9013
rect 11216 8763 11223 9813
rect 11276 9747 11283 10023
rect 11276 9536 11283 9593
rect 11256 9467 11263 9503
rect 11256 9207 11263 9353
rect 11276 9236 11283 9333
rect 11316 9147 11323 9203
rect 11196 8756 11223 8763
rect 11056 8508 11063 8573
rect 11136 8496 11143 8593
rect 11056 8463 11063 8494
rect 11056 8456 11083 8463
rect 10936 8316 10963 8323
rect 10896 8127 10903 8183
rect 10916 8107 10923 8173
rect 10936 8147 10943 8316
rect 11076 8227 11083 8456
rect 11116 8327 11123 8463
rect 11196 8243 11203 8756
rect 11296 8687 11303 8734
rect 11316 8707 11323 8833
rect 11236 8247 11243 8673
rect 11336 8667 11343 10532
rect 11176 8236 11203 8243
rect 10773 7980 10787 7993
rect 10776 7976 10783 7980
rect 10836 7940 10843 7943
rect 10833 7927 10847 7940
rect 10773 7680 10787 7693
rect 10816 7687 10823 7833
rect 10876 7807 10883 7993
rect 10896 7783 10903 8073
rect 10876 7776 10903 7783
rect 10776 7676 10783 7680
rect 10676 7527 10683 7593
rect 10636 7387 10643 7423
rect 10676 7367 10683 7423
rect 10716 7367 10723 7633
rect 10736 7407 10743 7613
rect 10756 7327 10763 7632
rect 10596 7187 10603 7313
rect 10796 7287 10803 7643
rect 10836 7527 10843 7652
rect 10876 7567 10883 7776
rect 10896 7607 10903 7663
rect 10896 7547 10903 7593
rect 10853 7460 10867 7473
rect 10856 7456 10863 7460
rect 10896 7456 10903 7512
rect 10916 7487 10923 7654
rect 10876 7420 10883 7423
rect 10873 7407 10887 7420
rect 10516 7136 10563 7143
rect 10396 6906 10403 6952
rect 10456 6936 10463 6973
rect 10496 6936 10503 7013
rect 10536 6927 10543 7113
rect 10476 6707 10483 6903
rect 10576 6867 10583 7143
rect 10596 7007 10603 7133
rect 10596 6906 10603 6972
rect 10576 6523 10583 6773
rect 10616 6747 10623 7253
rect 10756 7136 10763 7273
rect 10856 7007 10863 7393
rect 10936 7183 10943 8033
rect 11053 7980 11067 7993
rect 11056 7976 11063 7980
rect 11036 7887 11043 7943
rect 11076 7847 11083 7943
rect 10916 7176 10943 7183
rect 10876 7083 10883 7143
rect 10876 7076 10893 7083
rect 10716 6936 10723 6993
rect 10696 6787 10703 6903
rect 10676 6627 10683 6753
rect 10556 6516 10583 6523
rect 10316 6416 10343 6423
rect 10133 6120 10147 6133
rect 10176 6127 10183 6273
rect 10136 6116 10143 6120
rect 10056 6087 10063 6114
rect 10036 5983 10043 6073
rect 10036 5976 10063 5983
rect 10056 5908 10063 5976
rect 10116 5927 10123 6083
rect 10156 6047 10163 6083
rect 10056 5876 10083 5883
rect 9876 5596 9883 5633
rect 9913 5600 9927 5613
rect 9916 5596 9923 5600
rect 9856 5427 9863 5563
rect 9896 5560 9903 5563
rect 9893 5547 9907 5560
rect 9816 5356 9843 5363
rect 9756 4576 9783 4583
rect 9596 4336 9603 4372
rect 9576 4247 9583 4303
rect 9616 4283 9623 4292
rect 9596 4276 9623 4283
rect 9416 3816 9423 3852
rect 9336 3787 9343 3814
rect 9396 3780 9403 3783
rect 9356 3687 9363 3773
rect 9393 3767 9407 3780
rect 9436 3727 9443 3783
rect 9256 3503 9263 3633
rect 9336 3507 9343 3553
rect 9236 3496 9263 3503
rect 9356 3496 9363 3573
rect 9096 3476 9123 3483
rect 9096 3447 9103 3476
rect 9113 3427 9127 3433
rect 9156 3427 9163 3483
rect 9216 3327 9223 3493
rect 9116 3260 9123 3263
rect 9156 3260 9163 3263
rect 9113 3247 9127 3260
rect 9153 3247 9167 3260
rect 8976 2767 8983 2993
rect 9056 2867 9063 2952
rect 8996 2756 9003 2833
rect 9016 2747 9023 2813
rect 9053 2768 9067 2773
rect 9036 2547 9043 2713
rect 9076 2523 9083 3153
rect 9096 2547 9103 3053
rect 9056 2516 9083 2523
rect 8796 1987 8803 2223
rect 8836 2220 8843 2223
rect 8833 2207 8847 2220
rect 8896 2187 8903 2433
rect 8936 2407 8943 2443
rect 9016 2367 9023 2493
rect 9036 2467 9043 2493
rect 8696 1920 8703 1923
rect 8656 1767 8663 1913
rect 8693 1907 8707 1920
rect 8736 1748 8743 1893
rect 8756 1847 8763 1954
rect 8716 1647 8723 1703
rect 8756 1700 8763 1703
rect 8753 1687 8767 1700
rect 8796 1627 8803 1733
rect 8816 1687 8823 2013
rect 8533 1220 8547 1233
rect 8536 1216 8543 1220
rect 8476 1180 8483 1183
rect 8473 1167 8487 1180
rect 8576 1127 8583 1403
rect 8656 1367 8663 1413
rect 8676 1407 8683 1453
rect 8616 1167 8623 1233
rect 8676 1228 8683 1353
rect 8716 1248 8723 1273
rect 8736 1243 8743 1533
rect 8756 1267 8763 1613
rect 8796 1487 8803 1573
rect 8816 1487 8823 1673
rect 8836 1507 8843 1954
rect 8856 1887 8863 1973
rect 8916 1968 8923 2133
rect 8936 2047 8943 2313
rect 9016 2287 9023 2353
rect 8956 2107 8963 2253
rect 8976 2226 8983 2273
rect 9036 2256 9043 2453
rect 9056 2327 9063 2516
rect 9116 2427 9123 3173
rect 9136 2967 9143 3013
rect 9136 2807 9143 2893
rect 9156 2783 9163 3212
rect 9176 2927 9183 3233
rect 9216 3227 9223 3292
rect 9256 3266 9263 3453
rect 9196 3007 9203 3193
rect 9233 3000 9247 3013
rect 9276 3007 9283 3333
rect 9296 3247 9303 3293
rect 9316 3023 9323 3313
rect 9413 3300 9427 3313
rect 9416 3296 9423 3300
rect 9396 3247 9403 3263
rect 9376 3236 9393 3243
rect 9376 3047 9383 3236
rect 9496 3167 9503 3673
rect 9536 3500 9543 3503
rect 9516 3267 9523 3493
rect 9533 3487 9547 3500
rect 9496 3107 9503 3153
rect 9516 3087 9523 3133
rect 9536 3047 9543 3473
rect 9556 3247 9563 4093
rect 9596 3967 9603 4276
rect 9636 4227 9643 4253
rect 9613 4040 9627 4054
rect 9616 4036 9623 4040
rect 9676 4003 9683 4393
rect 9656 3996 9683 4003
rect 9656 3987 9663 3996
rect 9647 3976 9663 3987
rect 9647 3973 9660 3976
rect 9616 3780 9623 3783
rect 9613 3767 9627 3780
rect 9616 3528 9623 3713
rect 9616 3503 9623 3514
rect 9596 3496 9623 3503
rect 9636 3487 9643 3513
rect 9576 3327 9583 3373
rect 9636 3367 9643 3413
rect 9656 3296 9663 3333
rect 9676 3307 9683 3413
rect 9556 3107 9563 3153
rect 9596 3127 9603 3252
rect 9616 3183 9623 3213
rect 9636 3207 9643 3263
rect 9616 3176 9643 3183
rect 9316 3016 9343 3023
rect 9236 2996 9243 3000
rect 9296 2947 9303 2983
rect 9136 2776 9163 2783
rect 9136 2627 9143 2776
rect 9156 2476 9163 2753
rect 9176 2567 9183 2853
rect 9196 2476 9203 2573
rect 9216 2527 9223 2873
rect 9276 2776 9283 2913
rect 9316 2907 9323 2973
rect 9256 2740 9263 2743
rect 9253 2727 9267 2740
rect 9236 2476 9243 2713
rect 9296 2687 9303 2743
rect 9276 2467 9283 2553
rect 9296 2446 9303 2573
rect 9336 2446 9343 3016
rect 9396 2627 9403 2974
rect 9636 2927 9643 3176
rect 9676 3167 9683 3253
rect 9676 3023 9683 3093
rect 9696 3067 9703 4413
rect 9716 4227 9723 4523
rect 9716 3507 9723 4033
rect 9736 3427 9743 4353
rect 9716 3027 9723 3293
rect 9676 3016 9703 3023
rect 9416 2647 9423 2853
rect 9436 2440 9443 2443
rect 9076 2256 9083 2333
rect 9176 2307 9183 2353
rect 9196 2267 9203 2373
rect 9396 2367 9403 2432
rect 9433 2427 9447 2440
rect 9176 2236 9203 2243
rect 8956 1968 8963 1993
rect 8856 1707 8863 1873
rect 8896 1763 8903 1913
rect 8973 1907 8987 1913
rect 8876 1756 8903 1763
rect 8796 1436 8803 1473
rect 8833 1440 8847 1453
rect 8836 1436 8843 1440
rect 8816 1347 8823 1403
rect 8853 1387 8867 1393
rect 8736 1236 8763 1243
rect 8756 1216 8763 1236
rect 8793 1220 8807 1233
rect 8796 1216 8803 1220
rect 8336 627 8343 663
rect 8456 647 8463 953
rect 8476 887 8483 993
rect 8176 416 8203 423
rect 8196 396 8203 416
rect 8216 247 8223 363
rect 8296 207 8303 493
rect 8376 307 8383 363
rect 8100 203 8113 207
rect 8096 193 8113 203
rect 8096 176 8103 193
rect 8293 180 8307 193
rect 8296 176 8303 180
rect 8076 140 8083 143
rect 8073 127 8087 140
rect 8116 47 8123 143
rect 8156 127 8163 174
rect 8320 143 8333 147
rect 8316 136 8333 143
rect 8320 133 8333 136
rect 8416 127 8423 363
rect 8436 107 8443 253
rect 8456 143 8463 413
rect 8496 247 8503 673
rect 8516 307 8523 1053
rect 8556 916 8563 1013
rect 8656 928 8663 1172
rect 8736 1167 8743 1183
rect 8727 1156 8743 1167
rect 8727 1153 8740 1156
rect 8776 1147 8783 1183
rect 8596 767 8603 793
rect 8596 696 8603 753
rect 8556 547 8563 663
rect 8616 627 8623 853
rect 8636 707 8643 793
rect 8576 427 8583 473
rect 8616 427 8623 613
rect 8573 400 8587 413
rect 8613 400 8627 413
rect 8656 407 8663 914
rect 8576 396 8583 400
rect 8616 396 8623 400
rect 8596 267 8603 363
rect 8456 136 8473 143
rect 8487 143 8500 147
rect 8487 136 8503 143
rect 8487 133 8500 136
rect 8536 67 8543 143
rect 8576 47 8583 132
rect 8596 27 8603 253
rect 8616 67 8623 293
rect 8636 87 8643 352
rect 8676 327 8683 914
rect 8696 708 8703 1033
rect 8716 207 8723 973
rect 8736 887 8743 1133
rect 8836 1047 8843 1253
rect 8876 1247 8883 1756
rect 8896 1547 8903 1734
rect 8996 1647 9003 2213
rect 9056 2207 9063 2223
rect 9047 2196 9063 2207
rect 9047 2193 9060 2196
rect 9016 1927 9023 2173
rect 9036 1907 9043 1954
rect 9076 1927 9083 2193
rect 9096 2167 9103 2223
rect 9136 2067 9143 2203
rect 9196 2087 9203 2236
rect 9296 2107 9303 2243
rect 9196 2076 9213 2087
rect 9200 2073 9213 2076
rect 9116 2007 9123 2033
rect 9316 2027 9323 2073
rect 9193 1960 9207 1973
rect 9196 1956 9203 1960
rect 9096 1687 9103 1954
rect 9176 1920 9183 1923
rect 9173 1907 9187 1920
rect 9136 1736 9143 1853
rect 9193 1747 9207 1753
rect 9216 1747 9223 1773
rect 9236 1707 9243 1893
rect 9256 1807 9263 1993
rect 9396 1956 9403 1993
rect 9436 1867 9443 2353
rect 9456 2307 9463 2373
rect 9473 2240 9487 2253
rect 9476 2236 9483 2240
rect 9153 1687 9167 1692
rect 9107 1533 9113 1547
rect 8856 1187 8863 1213
rect 8856 1067 8863 1133
rect 8896 1067 8903 1473
rect 8916 1467 8923 1533
rect 8916 1287 8923 1413
rect 8956 1367 8963 1493
rect 9073 1440 9087 1453
rect 9076 1436 9083 1440
rect 8976 1347 8983 1434
rect 8996 1347 9003 1393
rect 9016 1367 9023 1403
rect 9076 1347 9083 1373
rect 9016 1247 9023 1273
rect 8973 1220 8987 1233
rect 9013 1220 9027 1233
rect 8976 1216 8983 1220
rect 9016 1216 9023 1220
rect 8796 916 8803 993
rect 8896 967 8903 1053
rect 8996 1027 9003 1183
rect 8833 928 8847 933
rect 9016 916 9023 953
rect 9056 916 9063 1253
rect 9116 1247 9123 1433
rect 9136 1347 9143 1553
rect 9156 1407 9163 1533
rect 9176 1307 9183 1633
rect 9196 1363 9203 1693
rect 9276 1607 9283 1773
rect 9236 1487 9243 1533
rect 9216 1407 9223 1453
rect 9296 1448 9303 1853
rect 9196 1356 9223 1363
rect 8736 347 8743 773
rect 8776 747 8783 883
rect 8816 880 8823 883
rect 8813 867 8827 880
rect 8816 696 8863 703
rect 8796 660 8803 663
rect 8793 647 8807 660
rect 8756 367 8763 553
rect 8856 507 8863 696
rect 8876 587 8883 693
rect 8936 627 8943 893
rect 8956 847 8963 913
rect 8996 767 9003 833
rect 9036 767 9043 883
rect 9096 867 9103 913
rect 9076 666 9083 713
rect 9116 667 9123 993
rect 8996 627 9003 663
rect 8996 396 9003 433
rect 8813 347 8827 352
rect 8856 267 8863 333
rect 8716 176 8723 193
rect 8876 146 8883 393
rect 8956 307 8963 394
rect 9136 287 9143 1293
rect 9216 1228 9223 1356
rect 9156 407 9163 1214
rect 9236 1127 9243 1173
rect 9176 807 9183 1013
rect 9236 916 9243 1033
rect 9256 963 9263 1353
rect 9276 987 9283 1403
rect 9296 1147 9303 1214
rect 9256 956 9283 963
rect 9216 880 9223 883
rect 9196 767 9203 873
rect 9213 867 9227 880
rect 9276 807 9283 956
rect 9196 703 9203 753
rect 9236 727 9243 753
rect 9227 716 9243 727
rect 9227 713 9240 716
rect 9196 696 9223 703
rect 9176 507 9183 694
rect 9236 527 9243 663
rect 9316 627 9323 1793
rect 9333 1767 9347 1773
rect 9376 1627 9383 1692
rect 9416 1607 9423 1703
rect 9256 503 9263 533
rect 9236 496 9263 503
rect 9176 307 9183 493
rect 9236 396 9243 496
rect 9296 427 9303 493
rect 9336 487 9343 1172
rect 9356 887 9363 1493
rect 9376 1247 9383 1592
rect 9456 1567 9463 2033
rect 9496 1947 9503 2293
rect 9516 2243 9523 2373
rect 9536 2267 9543 2833
rect 9556 2667 9563 2774
rect 9556 2307 9563 2473
rect 9576 2307 9583 2873
rect 9736 2867 9743 3373
rect 9756 3047 9763 4576
rect 9776 4527 9783 4554
rect 9796 4427 9803 4893
rect 9816 4867 9823 5273
rect 9836 5067 9843 5356
rect 9836 5027 9843 5053
rect 9816 4816 9833 4823
rect 9796 4336 9803 4392
rect 9816 4367 9823 4816
rect 9856 4603 9863 5233
rect 9916 5187 9923 5513
rect 9936 5287 9943 5374
rect 9956 5127 9963 5693
rect 9976 5307 9983 5753
rect 9916 5076 9923 5113
rect 9896 4967 9903 5043
rect 9916 4826 9923 4933
rect 9956 4820 9963 4823
rect 9953 4807 9967 4820
rect 9996 4807 10003 5733
rect 10056 5727 10063 5876
rect 10016 5247 10023 5693
rect 10096 5596 10103 5633
rect 10156 5627 10163 6033
rect 10176 5643 10183 5893
rect 10196 5866 10203 6153
rect 10176 5636 10203 5643
rect 10147 5623 10163 5627
rect 10147 5616 10183 5623
rect 10147 5613 10160 5616
rect 10156 5566 10163 5593
rect 10036 5347 10043 5552
rect 10113 5547 10127 5552
rect 10156 5447 10163 5552
rect 10093 5388 10107 5393
rect 10176 5387 10183 5616
rect 10196 5566 10203 5636
rect 10116 5307 10123 5343
rect 10156 5287 10163 5343
rect 10016 5046 10023 5093
rect 10016 4827 10023 4853
rect 9847 4596 9863 4603
rect 9836 4336 9843 4593
rect 9936 4556 9943 4733
rect 9856 4447 9863 4554
rect 9867 4436 9883 4443
rect 9876 4347 9883 4436
rect 9816 4267 9823 4292
rect 9896 4006 9903 4393
rect 9916 4307 9923 4523
rect 9776 3527 9783 3913
rect 9856 3816 9863 3971
rect 9896 3816 9903 3873
rect 9936 3827 9943 4333
rect 9956 3987 9963 4512
rect 10016 4467 10023 4633
rect 10036 4443 10043 5253
rect 10056 4927 10063 5173
rect 10076 4747 10083 5273
rect 10196 5207 10203 5373
rect 10216 5267 10223 6313
rect 10133 5080 10147 5093
rect 10136 5076 10143 5080
rect 10096 5007 10103 5073
rect 10196 5043 10203 5063
rect 10156 5036 10203 5043
rect 10236 4907 10243 6133
rect 10256 5827 10263 6113
rect 10256 5127 10263 5713
rect 10276 5707 10283 6253
rect 10316 6148 10323 6416
rect 10376 6247 10383 6352
rect 10436 6227 10443 6393
rect 10476 6167 10483 6473
rect 10353 5900 10367 5913
rect 10396 5907 10403 6113
rect 10356 5896 10363 5900
rect 10376 5643 10383 5852
rect 10356 5636 10383 5643
rect 10356 5607 10363 5636
rect 10416 5583 10423 6133
rect 10456 6087 10463 6113
rect 10456 5683 10463 5993
rect 10476 5866 10483 6153
rect 10476 5707 10483 5793
rect 10496 5727 10503 6513
rect 10556 6487 10563 6516
rect 10576 6416 10583 6493
rect 10596 6447 10603 6553
rect 10696 6507 10703 6733
rect 10516 6327 10523 6373
rect 10536 6307 10543 6413
rect 10696 6407 10703 6453
rect 10716 6396 10723 6613
rect 10736 6527 10743 6893
rect 10756 6503 10763 6993
rect 10896 6767 10903 7073
rect 10916 6867 10923 6903
rect 10836 6567 10843 6603
rect 10916 6547 10923 6853
rect 10936 6606 10943 6633
rect 10956 6527 10963 7553
rect 10976 6867 10983 7513
rect 11016 7426 11023 7473
rect 11056 7468 11063 7493
rect 11127 7483 11140 7487
rect 11127 7473 11143 7483
rect 11136 7456 11143 7473
rect 11116 7420 11123 7423
rect 10736 6496 10763 6503
rect 10736 6467 10743 6496
rect 10596 6363 10603 6383
rect 10576 6356 10603 6363
rect 10536 6147 10543 6293
rect 10533 6120 10547 6133
rect 10536 6116 10543 6120
rect 10576 6116 10583 6356
rect 10616 6116 10623 6253
rect 10636 6127 10643 6383
rect 10516 5827 10523 5913
rect 10556 5896 10563 6013
rect 10596 6007 10603 6083
rect 10656 5927 10663 6193
rect 10616 5827 10623 5863
rect 10656 5727 10663 5892
rect 10676 5767 10683 6033
rect 10456 5676 10483 5683
rect 10396 5576 10423 5583
rect 10336 5527 10343 5563
rect 10276 5347 10283 5513
rect 10336 5407 10343 5473
rect 10333 5380 10347 5393
rect 10396 5387 10403 5576
rect 10436 5387 10443 5583
rect 10476 5487 10483 5676
rect 10616 5576 10623 5713
rect 10716 5667 10723 6313
rect 10736 6067 10743 6414
rect 10836 6287 10843 6403
rect 10813 6120 10827 6133
rect 10816 6116 10823 6120
rect 10776 6076 10803 6083
rect 10736 5643 10743 5953
rect 10716 5636 10743 5643
rect 10716 5407 10723 5636
rect 10756 5627 10763 6073
rect 10776 6047 10783 6076
rect 10796 5896 10803 6053
rect 10876 5947 10883 6273
rect 10916 6086 10923 6113
rect 10916 6047 10923 6072
rect 10833 5900 10847 5913
rect 10836 5896 10843 5900
rect 10776 5747 10783 5832
rect 10816 5807 10823 5863
rect 10776 5616 10783 5733
rect 10856 5627 10863 5831
rect 10896 5763 10903 5913
rect 10876 5756 10903 5763
rect 10816 5583 10823 5613
rect 10336 5376 10343 5380
rect 10736 5383 10743 5583
rect 10816 5576 10843 5583
rect 10856 5427 10863 5573
rect 10716 5376 10743 5383
rect 10433 5360 10447 5373
rect 10436 5356 10443 5360
rect 10296 5267 10303 5333
rect 10356 5307 10363 5333
rect 10416 5207 10423 5354
rect 10476 5227 10483 5373
rect 10616 5327 10623 5363
rect 10427 5196 10443 5203
rect 10436 5147 10443 5196
rect 10253 5047 10267 5052
rect 10296 4947 10303 5113
rect 10433 5060 10447 5073
rect 10436 5056 10443 5060
rect 10536 5047 10543 5213
rect 10616 5207 10623 5253
rect 10716 5207 10723 5376
rect 10736 5356 10743 5376
rect 10816 5327 10823 5393
rect 10756 5227 10763 5313
rect 10776 5247 10783 5323
rect 10636 5067 10643 5193
rect 10776 5167 10783 5233
rect 10716 5108 10723 5153
rect 10116 4527 10123 4854
rect 10136 4563 10143 4673
rect 10156 4647 10163 4823
rect 10236 4667 10243 4812
rect 10216 4568 10223 4633
rect 10276 4627 10283 4854
rect 10296 4647 10303 4933
rect 10476 4856 10483 4913
rect 10456 4727 10463 4823
rect 10536 4687 10543 5033
rect 10656 4856 10663 5033
rect 10676 4727 10683 4823
rect 10136 4556 10163 4563
rect 10016 4436 10043 4443
rect 9976 3963 9983 4193
rect 9996 3987 10003 4033
rect 10016 3983 10023 4436
rect 10076 4336 10083 4393
rect 10096 4267 10103 4303
rect 10036 4036 10043 4253
rect 10116 4247 10123 4373
rect 10136 4267 10143 4556
rect 10176 4287 10183 4523
rect 10176 4227 10183 4273
rect 10096 4036 10103 4173
rect 10196 4083 10203 4393
rect 10236 4187 10243 4613
rect 10716 4587 10723 5094
rect 10256 4507 10263 4543
rect 10276 4336 10283 4453
rect 10316 4407 10323 4532
rect 10356 4443 10363 4534
rect 10356 4436 10383 4443
rect 10296 4267 10303 4303
rect 10336 4207 10343 4303
rect 10376 4127 10383 4436
rect 10596 4427 10603 4574
rect 10456 4247 10463 4333
rect 10476 4207 10483 4413
rect 10576 4348 10583 4373
rect 10656 4316 10663 4513
rect 10756 4427 10763 5093
rect 10793 5080 10807 5093
rect 10796 5076 10803 5080
rect 10816 5040 10823 5043
rect 10813 5027 10827 5040
rect 10856 4947 10863 5273
rect 10876 5047 10883 5756
rect 10916 5627 10923 5853
rect 10896 5387 10903 5583
rect 10893 5360 10907 5373
rect 10916 5368 10923 5573
rect 10936 5447 10943 6193
rect 10976 6127 10983 6633
rect 10996 6587 11003 6813
rect 11076 6667 11083 7412
rect 11113 7407 11127 7420
rect 11116 7156 11123 7293
rect 11156 6907 11163 7154
rect 11036 6600 11043 6603
rect 11033 6587 11047 6600
rect 11016 6396 11023 6533
rect 11036 6187 11043 6513
rect 11096 6403 11103 6553
rect 11076 6396 11103 6403
rect 11096 6267 11103 6396
rect 10956 6027 10963 6114
rect 11033 6120 11047 6133
rect 11036 6116 11043 6120
rect 10976 5967 10983 6033
rect 10956 5867 10963 5894
rect 10976 5847 10983 5932
rect 10996 5847 11003 5973
rect 11056 5947 11063 6083
rect 11096 6027 11103 6173
rect 11116 5987 11123 6653
rect 11076 5896 11083 5973
rect 11096 5907 11103 5933
rect 11076 5747 11083 5833
rect 11076 5607 11083 5712
rect 11096 5707 11103 5853
rect 11116 5727 11123 5893
rect 11136 5747 11143 6733
rect 11156 5727 11163 6633
rect 11096 5583 11103 5633
rect 11076 5576 11103 5583
rect 10896 5356 10903 5360
rect 10896 5007 10903 5093
rect 10916 4983 10923 5313
rect 10936 5007 10943 5433
rect 11176 5387 11183 8236
rect 11233 8220 11247 8233
rect 11236 8216 11243 8220
rect 11296 8147 11303 8652
rect 11316 8187 11323 8313
rect 11196 7907 11203 8133
rect 11216 7923 11223 8033
rect 11256 7976 11263 8113
rect 11296 7984 11303 8053
rect 11296 7977 11343 7984
rect 11276 7923 11283 7943
rect 11216 7916 11243 7923
rect 11236 7696 11243 7916
rect 11256 7916 11283 7923
rect 11256 7867 11263 7916
rect 11276 7643 11283 7893
rect 11296 7667 11303 7773
rect 11276 7636 11303 7643
rect 11196 6747 11203 7453
rect 11216 6936 11243 6943
rect 11196 6047 11203 6712
rect 11216 6587 11223 6936
rect 11296 6727 11303 7636
rect 11316 7467 11323 7943
rect 11316 6647 11323 7353
rect 11236 6327 11243 6593
rect 11256 6587 11263 6603
rect 11236 6116 11243 6213
rect 11256 6207 11263 6573
rect 11296 6567 11303 6603
rect 11336 6587 11343 7977
rect 11196 5827 11203 6012
rect 11196 5647 11203 5713
rect 11216 5667 11223 6013
rect 11296 5896 11303 6013
rect 11316 5860 11323 5863
rect 11313 5847 11327 5860
rect 11236 5628 11243 5833
rect 11276 5647 11283 5813
rect 11300 5723 11313 5727
rect 11296 5713 11313 5723
rect 11296 5667 11303 5713
rect 11256 5367 11263 5533
rect 11176 5356 11203 5363
rect 10956 5047 10963 5213
rect 11176 5207 11183 5356
rect 10996 5076 11003 5193
rect 10916 4976 10943 4983
rect 10873 4860 10887 4873
rect 10876 4856 10883 4860
rect 10856 4467 10863 4823
rect 10556 4267 10563 4303
rect 10616 4207 10623 4283
rect 10176 4076 10203 4083
rect 10176 4023 10183 4076
rect 10136 4020 10143 4023
rect 10133 4007 10147 4020
rect 10056 4000 10063 4003
rect 10053 3987 10067 4000
rect 10176 4016 10203 4023
rect 10016 3976 10043 3983
rect 9976 3956 10003 3963
rect 9816 3567 9823 3813
rect 9916 3567 9923 3772
rect 9776 3387 9783 3413
rect 9776 3247 9783 3352
rect 9796 3307 9803 3453
rect 9816 3367 9823 3483
rect 9836 3296 9843 3433
rect 9856 3347 9863 3483
rect 9873 3300 9887 3313
rect 9896 3307 9903 3553
rect 9956 3543 9963 3573
rect 9936 3536 9963 3543
rect 9916 3467 9923 3514
rect 9936 3447 9943 3536
rect 9876 3296 9883 3300
rect 9816 3260 9823 3263
rect 9796 3207 9803 3253
rect 9813 3247 9827 3260
rect 9856 3243 9863 3263
rect 9916 3247 9923 3313
rect 9836 3236 9863 3243
rect 9596 2487 9603 2853
rect 9616 2476 9623 2573
rect 9636 2507 9643 2793
rect 9673 2780 9687 2793
rect 9756 2787 9763 3012
rect 9720 2783 9733 2787
rect 9676 2776 9683 2780
rect 9716 2776 9733 2783
rect 9720 2773 9733 2776
rect 9516 2236 9543 2243
rect 9476 1667 9483 1912
rect 9496 1467 9503 1933
rect 9516 1707 9523 2193
rect 9556 2127 9563 2253
rect 9536 1847 9543 1993
rect 9576 1956 9583 2053
rect 9596 2047 9603 2413
rect 9616 2007 9623 2293
rect 9636 2227 9643 2443
rect 9656 2207 9663 2433
rect 9676 2147 9683 2513
rect 9696 2347 9703 2732
rect 9716 2267 9723 2713
rect 9756 2707 9763 2752
rect 9736 2347 9743 2653
rect 9736 2256 9743 2293
rect 9756 2287 9763 2493
rect 9776 2447 9783 3013
rect 9687 2136 9703 2143
rect 9656 1967 9663 2093
rect 9676 1927 9683 1954
rect 9640 1923 9653 1927
rect 9496 1436 9503 1453
rect 9416 1367 9423 1434
rect 9416 1216 9423 1313
rect 9387 1113 9393 1127
rect 9436 1087 9443 1183
rect 9476 1047 9483 1353
rect 9536 1007 9543 1734
rect 9556 1706 9563 1873
rect 9596 1827 9603 1923
rect 9636 1916 9653 1923
rect 9640 1913 9653 1916
rect 9616 1736 9623 1873
rect 9656 1736 9663 1833
rect 9496 907 9503 993
rect 9456 807 9463 883
rect 9476 727 9483 853
rect 9516 727 9523 933
rect 9336 247 9343 413
rect 9396 387 9403 713
rect 9433 700 9447 713
rect 9436 696 9443 700
rect 9476 696 9483 713
rect 9456 507 9463 663
rect 9436 360 9443 363
rect 9433 347 9447 360
rect 9476 343 9483 363
rect 9456 336 9483 343
rect 9396 267 9403 293
rect 9456 267 9463 336
rect 8736 67 8743 132
rect 8876 87 8883 132
rect 8896 47 8903 173
rect 8916 146 8923 193
rect 8996 107 9003 143
rect 9136 87 9143 173
rect 9336 147 9343 233
rect 9433 180 9447 193
rect 9436 176 9443 180
rect 9220 143 9233 147
rect 9176 140 9183 143
rect 9173 127 9187 140
rect 9216 136 9233 143
rect 9220 133 9233 136
rect 9227 126 9240 127
rect 9227 113 9233 126
rect 9316 87 9323 132
rect 9333 107 9347 112
rect 8976 27 8983 73
rect 9536 67 9543 793
rect 9556 507 9563 1653
rect 9576 1407 9583 1693
rect 9636 1683 9643 1703
rect 9616 1676 9643 1683
rect 9596 1447 9603 1533
rect 9616 1327 9623 1676
rect 9636 1567 9643 1593
rect 9636 1307 9643 1473
rect 9696 1468 9703 2136
rect 9716 1927 9723 2013
rect 9796 1988 9803 3033
rect 9816 2987 9823 3113
rect 9836 3027 9843 3236
rect 9876 3063 9883 3113
rect 9876 3056 9903 3063
rect 9836 2927 9843 2992
rect 9836 2727 9843 2833
rect 9816 2567 9823 2693
rect 9816 2476 9823 2553
rect 9856 2507 9863 3053
rect 9896 2996 9903 3056
rect 9936 3003 9943 3293
rect 9956 3107 9963 3513
rect 9976 3247 9983 3733
rect 9996 3527 10003 3956
rect 10016 3808 10023 3913
rect 10036 3863 10043 3976
rect 10056 3887 10063 3973
rect 10176 3927 10183 4016
rect 10236 4007 10243 4113
rect 10536 4107 10543 4193
rect 10536 4068 10543 4093
rect 10496 4016 10523 4023
rect 10036 3856 10063 3863
rect 10056 3747 10063 3856
rect 10296 3803 10303 3913
rect 10476 3847 10483 4014
rect 10173 3647 10187 3653
rect 10036 3516 10043 3553
rect 10073 3520 10087 3533
rect 10076 3516 10083 3520
rect 9936 2996 9963 3003
rect 9916 2960 9923 2963
rect 9913 2947 9927 2960
rect 9956 2827 9963 2996
rect 9836 2087 9843 2273
rect 9856 2127 9863 2432
rect 9716 1748 9723 1773
rect 9736 1487 9743 1953
rect 9756 1443 9763 1973
rect 9836 1956 9843 1993
rect 9776 1707 9783 1813
rect 9856 1736 9863 1913
rect 9876 1867 9883 2813
rect 9896 2627 9903 2743
rect 9896 2187 9903 2493
rect 9956 2387 9963 2743
rect 9976 2607 9983 3153
rect 9996 3127 10003 3293
rect 10016 3267 10023 3373
rect 10036 3307 10043 3413
rect 10096 3347 10103 3483
rect 10136 3387 10143 3553
rect 10156 3427 10163 3613
rect 10176 3447 10183 3493
rect 10196 3447 10203 3803
rect 10296 3796 10323 3803
rect 10296 3667 10303 3796
rect 10356 3687 10363 3763
rect 10216 3487 10223 3514
rect 10236 3487 10243 3633
rect 10316 3516 10323 3593
rect 10356 3527 10363 3553
rect 10056 3296 10063 3333
rect 10156 3276 10163 3413
rect 10236 3407 10243 3433
rect 9996 2727 10003 3092
rect 9976 2307 9983 2533
rect 9896 1927 9903 1953
rect 9916 1807 9923 2213
rect 9936 2147 9943 2193
rect 9956 2167 9963 2223
rect 10016 2207 10023 3232
rect 10036 2747 10043 2893
rect 10056 2788 10063 3233
rect 10076 3207 10083 3263
rect 10076 3047 10083 3113
rect 10096 2747 10103 2933
rect 10116 2907 10123 2963
rect 10156 2776 10163 2983
rect 10196 2947 10203 3393
rect 10216 3276 10223 3353
rect 10256 3347 10263 3453
rect 10296 3447 10303 3483
rect 10336 3480 10343 3483
rect 10333 3467 10347 3480
rect 10336 3427 10343 3453
rect 10376 3407 10383 3453
rect 10396 3427 10403 3493
rect 10416 3447 10423 3593
rect 10456 3547 10463 3833
rect 10476 3503 10483 3793
rect 10496 3747 10503 3993
rect 10516 3947 10523 4016
rect 10576 3907 10583 4133
rect 10676 4067 10683 4413
rect 10776 4247 10783 4323
rect 10916 4163 10923 4873
rect 10936 4767 10943 4976
rect 10956 4316 10963 4553
rect 10976 4306 10983 5013
rect 11016 4967 11023 5043
rect 11016 4807 11023 4953
rect 11056 4856 11063 4933
rect 11096 4856 11103 4993
rect 11136 4863 11143 5093
rect 11156 5046 11163 5133
rect 11136 4856 11163 4863
rect 11156 4826 11163 4856
rect 11116 4820 11123 4823
rect 11113 4807 11127 4820
rect 11176 4787 11183 5172
rect 11216 5083 11223 5313
rect 11236 5247 11243 5323
rect 11256 5123 11263 5313
rect 11276 5247 11283 5612
rect 11296 5587 11303 5613
rect 11296 5187 11303 5552
rect 11236 5120 11263 5123
rect 11233 5116 11263 5120
rect 11233 5107 11247 5116
rect 11196 5076 11223 5083
rect 10996 4556 11003 4633
rect 11056 4547 11063 4673
rect 11013 4320 11027 4333
rect 11016 4316 11023 4320
rect 10976 4207 10983 4292
rect 10916 4156 10943 4163
rect 10596 4020 10603 4023
rect 10593 4007 10607 4020
rect 10516 3786 10523 3893
rect 10636 3843 10643 4053
rect 10573 3820 10587 3833
rect 10616 3836 10643 3843
rect 10576 3816 10583 3820
rect 10616 3816 10623 3836
rect 10656 3827 10663 4023
rect 10596 3747 10603 3783
rect 10636 3747 10643 3783
rect 10696 3643 10703 4093
rect 10816 3816 10823 3873
rect 10853 3820 10867 3833
rect 10856 3816 10863 3820
rect 10836 3763 10843 3783
rect 10836 3756 10863 3763
rect 10696 3636 10723 3643
rect 10436 3496 10483 3503
rect 10436 3427 10443 3496
rect 10436 3387 10443 3413
rect 10456 3407 10463 3473
rect 10476 3403 10483 3433
rect 10476 3396 10503 3403
rect 10256 3247 10263 3333
rect 10076 2476 10083 2573
rect 9936 1907 9943 2053
rect 9956 1847 9963 1973
rect 9976 1923 9983 2193
rect 10036 2187 10043 2373
rect 9996 1967 10003 2173
rect 10016 2087 10023 2133
rect 10096 2107 10103 2712
rect 10016 1983 10023 2073
rect 10016 1976 10043 1983
rect 10036 1956 10043 1976
rect 10116 1927 10123 2693
rect 10136 2467 10143 2732
rect 10176 2303 10183 2593
rect 10196 2427 10203 2873
rect 10216 2827 10223 2983
rect 10236 2887 10243 2974
rect 10256 2587 10263 3233
rect 10396 3167 10403 3283
rect 10496 3223 10503 3396
rect 10516 3276 10523 3393
rect 10556 3240 10563 3243
rect 10553 3227 10567 3240
rect 10496 3216 10523 3223
rect 10416 2987 10423 3033
rect 10316 2740 10323 2743
rect 10313 2727 10327 2740
rect 10256 2476 10263 2513
rect 10176 2300 10203 2303
rect 10176 2296 10207 2300
rect 10193 2287 10207 2296
rect 10156 2220 10163 2223
rect 10153 2207 10167 2220
rect 10236 2223 10243 2443
rect 10276 2440 10283 2443
rect 10273 2427 10287 2440
rect 10356 2427 10363 2513
rect 10256 2226 10263 2293
rect 10216 2216 10243 2223
rect 9976 1916 10003 1923
rect 9916 1767 9923 1793
rect 9756 1436 9783 1443
rect 9576 447 9583 1233
rect 9656 1228 9663 1333
rect 9636 1147 9643 1183
rect 9596 947 9603 1073
rect 9596 886 9603 933
rect 9656 916 9663 993
rect 9696 767 9703 1333
rect 9716 847 9723 1293
rect 9736 886 9743 1053
rect 9653 700 9667 713
rect 9656 696 9663 700
rect 9696 696 9703 753
rect 9653 400 9667 413
rect 9656 396 9663 400
rect 9676 360 9683 363
rect 9673 347 9687 360
rect 9556 87 9563 193
rect 9576 187 9583 293
rect 9596 167 9603 233
rect 9656 176 9663 273
rect 9716 147 9723 613
rect 9736 347 9743 872
rect 9756 427 9763 1353
rect 9636 27 9643 132
rect 9676 87 9683 143
rect 9696 67 9703 113
rect 9736 47 9743 253
rect 9776 47 9783 1436
rect 9796 927 9803 1434
rect 9816 1406 9823 1613
rect 9836 1567 9843 1703
rect 9856 1587 9863 1653
rect 9836 1267 9843 1453
rect 9856 1406 9863 1573
rect 9876 1507 9883 1703
rect 9976 1547 9983 1734
rect 9936 1436 9943 1473
rect 9856 947 9863 993
rect 9916 967 9923 1253
rect 9956 1228 9963 1392
rect 9936 1047 9943 1093
rect 9856 916 9863 933
rect 9796 587 9803 913
rect 9916 886 9923 953
rect 9956 927 9963 1214
rect 9976 1027 9983 1253
rect 9856 667 9863 753
rect 9916 696 9923 833
rect 9976 666 9983 1013
rect 9796 146 9803 493
rect 9916 396 9923 493
rect 9816 366 9823 393
rect 9896 360 9903 363
rect 9893 347 9907 360
rect 9856 176 9863 313
rect 9836 140 9843 143
rect 9833 127 9847 140
rect 9936 107 9943 353
rect 9996 347 10003 1916
rect 10016 1847 10023 1923
rect 10056 1920 10063 1923
rect 10053 1907 10067 1920
rect 10016 1407 10023 1833
rect 10036 1223 10043 1853
rect 10096 1807 10103 1873
rect 10073 1740 10087 1753
rect 10076 1736 10083 1740
rect 10136 1743 10143 1873
rect 10127 1736 10143 1743
rect 10016 1216 10043 1223
rect 10056 1216 10063 1693
rect 10096 1687 10103 1703
rect 10096 1676 10113 1687
rect 10100 1673 10113 1676
rect 10076 1367 10083 1533
rect 10096 1267 10103 1553
rect 10156 1507 10163 1913
rect 10147 1480 10183 1483
rect 10147 1476 10187 1480
rect 10173 1467 10187 1476
rect 10196 1467 10203 2173
rect 10216 1667 10223 2216
rect 10276 1956 10283 2333
rect 10376 2287 10383 2813
rect 10496 2807 10503 3173
rect 10516 3067 10523 3216
rect 10556 3016 10563 3213
rect 10596 3027 10603 3393
rect 10716 3367 10723 3636
rect 10776 3536 10783 3673
rect 10796 3547 10803 3753
rect 10736 3500 10743 3503
rect 10733 3487 10747 3500
rect 10616 3227 10623 3313
rect 10616 3016 10623 3213
rect 10596 2887 10603 2973
rect 10616 2867 10623 2933
rect 10636 2907 10643 2974
rect 10436 2447 10443 2474
rect 10456 2387 10463 2793
rect 10476 2587 10483 2793
rect 10533 2780 10547 2793
rect 10536 2776 10543 2780
rect 10516 2740 10523 2743
rect 10513 2727 10527 2740
rect 10596 2736 10623 2743
rect 10533 2480 10547 2493
rect 10536 2476 10543 2480
rect 10516 2440 10523 2443
rect 10296 1987 10303 2273
rect 10316 2147 10323 2173
rect 10336 2007 10343 2273
rect 10433 2260 10447 2273
rect 10436 2256 10443 2260
rect 10256 1767 10263 1923
rect 10296 1887 10303 1923
rect 10236 1756 10253 1763
rect 10153 1440 10167 1453
rect 10216 1443 10223 1613
rect 10236 1483 10243 1756
rect 10276 1736 10283 1793
rect 10336 1767 10343 1972
rect 10356 1907 10363 2213
rect 10376 2127 10383 2223
rect 10416 2187 10423 2223
rect 10476 2207 10483 2433
rect 10513 2427 10527 2440
rect 10320 1746 10340 1747
rect 10320 1743 10333 1746
rect 10316 1736 10333 1743
rect 10320 1733 10333 1736
rect 10273 1667 10287 1673
rect 10236 1476 10263 1483
rect 10156 1436 10163 1440
rect 10196 1436 10223 1443
rect 10016 487 10023 1216
rect 10136 1227 10143 1403
rect 10176 1400 10183 1403
rect 10173 1387 10187 1400
rect 10156 1376 10173 1383
rect 10087 1133 10093 1147
rect 10116 1107 10123 1183
rect 10136 1067 10143 1173
rect 10136 1007 10143 1053
rect 10056 916 10063 993
rect 10136 883 10143 914
rect 10116 876 10143 883
rect 10016 146 10023 433
rect 10056 347 10063 733
rect 10116 696 10123 876
rect 10156 666 10163 1376
rect 10176 1127 10183 1214
rect 10076 656 10093 663
rect 10076 447 10083 656
rect 10076 367 10083 433
rect 10156 396 10163 573
rect 10076 176 10083 332
rect 10176 168 10183 993
rect 10196 827 10203 1293
rect 10216 1186 10223 1213
rect 10196 627 10203 694
rect 10216 666 10223 973
rect 10196 156 10203 293
rect 10216 166 10223 473
rect 10096 140 10103 143
rect 10093 127 10107 140
rect 10236 127 10243 1453
rect 10256 1406 10263 1476
rect 10256 1347 10263 1392
rect 10296 1247 10303 1493
rect 10316 1216 10323 1673
rect 10333 1467 10347 1473
rect 10356 1443 10363 1893
rect 10376 1527 10383 1953
rect 10396 1927 10403 2133
rect 10416 1867 10423 1954
rect 10396 1507 10403 1753
rect 10416 1707 10423 1813
rect 10336 1436 10363 1443
rect 10336 1387 10343 1436
rect 10336 1180 10343 1183
rect 10333 1167 10347 1180
rect 10253 1127 10267 1133
rect 10296 916 10303 1073
rect 10276 807 10283 872
rect 10336 787 10343 914
rect 10356 696 10363 1133
rect 10376 703 10383 1273
rect 10396 747 10403 1373
rect 10416 1186 10423 1233
rect 10416 847 10423 1073
rect 10436 803 10443 2193
rect 10496 2147 10503 2273
rect 10516 2207 10523 2373
rect 10536 2167 10543 2233
rect 10556 2226 10563 2433
rect 10556 1967 10563 2212
rect 10456 1787 10463 1913
rect 10496 1887 10503 1923
rect 10536 1920 10543 1923
rect 10533 1907 10547 1920
rect 10536 1736 10543 1893
rect 10556 1827 10563 1913
rect 10476 1667 10483 1703
rect 10516 1683 10523 1703
rect 10496 1676 10523 1683
rect 10456 967 10463 1433
rect 10476 1287 10483 1533
rect 10496 1307 10503 1676
rect 10516 1387 10523 1613
rect 10536 1247 10543 1493
rect 10576 1467 10583 2593
rect 10596 2347 10603 2493
rect 10616 2447 10623 2736
rect 10636 2447 10643 2872
rect 10656 2587 10663 2983
rect 10676 2607 10683 3353
rect 10756 3296 10763 3494
rect 10796 3407 10803 3493
rect 10796 3296 10803 3333
rect 10816 3327 10823 3673
rect 10836 3567 10843 3733
rect 10856 3563 10863 3756
rect 10876 3563 10883 3751
rect 10896 3567 10903 3773
rect 10856 3556 10883 3563
rect 10836 3467 10843 3503
rect 10836 3308 10843 3453
rect 10736 3127 10743 3263
rect 10776 3243 10783 3263
rect 10756 3236 10783 3243
rect 10756 3187 10763 3236
rect 10856 3207 10863 3493
rect 10876 3247 10883 3556
rect 10916 3547 10923 3733
rect 10896 3496 10923 3503
rect 10896 3227 10903 3473
rect 10916 3407 10923 3496
rect 10916 3207 10923 3393
rect 10776 3027 10783 3193
rect 10716 2667 10723 2853
rect 10776 2776 10783 2833
rect 10813 2780 10827 2793
rect 10816 2776 10823 2780
rect 10736 2476 10743 2774
rect 10796 2707 10803 2743
rect 10696 2227 10703 2433
rect 10716 2287 10723 2443
rect 10756 2407 10763 2443
rect 10596 1747 10603 1954
rect 10616 1887 10623 2173
rect 10656 2167 10663 2223
rect 10716 2207 10723 2273
rect 10756 2187 10763 2313
rect 10816 2287 10823 2474
rect 10813 2260 10827 2273
rect 10816 2256 10823 2260
rect 10856 2256 10863 2333
rect 10876 2307 10883 2873
rect 10776 2187 10783 2253
rect 10836 2207 10843 2223
rect 10836 2196 10853 2207
rect 10840 2193 10853 2196
rect 10616 1523 10623 1773
rect 10636 1547 10643 1993
rect 10656 1887 10663 2093
rect 10676 1926 10683 2013
rect 10756 1887 10763 1923
rect 10736 1736 10743 1833
rect 10796 1823 10803 1913
rect 10816 1847 10823 2193
rect 10796 1816 10823 1823
rect 10676 1706 10683 1733
rect 10756 1683 10763 1703
rect 10736 1676 10763 1683
rect 10736 1647 10743 1676
rect 10616 1516 10643 1523
rect 10596 1436 10603 1473
rect 10636 1448 10643 1516
rect 10576 1347 10583 1403
rect 10476 1176 10503 1183
rect 10476 1087 10483 1176
rect 10536 1127 10543 1183
rect 10496 947 10503 1093
rect 10616 1067 10623 1403
rect 10556 916 10563 953
rect 10536 847 10543 883
rect 10436 796 10453 803
rect 10376 696 10403 703
rect 10336 660 10343 663
rect 10333 647 10347 660
rect 10276 307 10283 453
rect 10336 427 10343 553
rect 10356 427 10363 493
rect 10396 467 10403 696
rect 10436 687 10443 713
rect 10296 327 10303 413
rect 10353 400 10367 413
rect 10356 396 10363 400
rect 10456 366 10463 793
rect 10596 703 10603 973
rect 10576 696 10603 703
rect 10496 447 10503 694
rect 10556 660 10563 663
rect 10553 647 10567 660
rect 10636 607 10643 1233
rect 10656 1147 10663 1393
rect 10536 407 10543 513
rect 10336 307 10343 363
rect 10476 267 10483 394
rect 10596 396 10603 433
rect 10636 396 10643 572
rect 10496 156 10503 393
rect 10676 126 10683 1453
rect 10716 1367 10723 1593
rect 10736 1407 10743 1633
rect 10756 1407 10763 1653
rect 10816 1607 10823 1816
rect 10836 1627 10843 2153
rect 10856 1667 10863 1893
rect 10876 1687 10883 2213
rect 10833 1440 10847 1453
rect 10836 1436 10843 1440
rect 10896 1443 10903 2773
rect 10916 2747 10923 3153
rect 10936 3027 10943 4156
rect 10996 4056 11003 4093
rect 11036 4007 11043 4053
rect 11056 4047 11063 4273
rect 10956 3867 10963 3973
rect 10956 3747 10963 3772
rect 10996 3767 11003 3913
rect 11016 3787 11023 3953
rect 11056 3816 11063 4033
rect 11076 3927 11083 4253
rect 11096 3967 11103 4753
rect 11116 4147 11123 4553
rect 11136 4003 11143 4773
rect 11196 4607 11203 5076
rect 11236 4967 11243 5043
rect 11156 4087 11163 4593
rect 11236 4567 11243 4953
rect 11316 4807 11323 5653
rect 11216 4520 11223 4523
rect 11213 4507 11227 4520
rect 11236 4027 11243 4133
rect 11136 3996 11163 4003
rect 11096 3816 11103 3853
rect 11076 3780 11083 3783
rect 11073 3767 11087 3780
rect 11116 3707 11123 3783
rect 11156 3767 11163 3996
rect 11076 3563 11083 3693
rect 11076 3556 11103 3563
rect 11096 3507 11103 3556
rect 11236 3536 11243 3673
rect 11256 3547 11263 4073
rect 10936 2727 10943 2913
rect 10956 2827 10963 2972
rect 10976 2787 10983 3013
rect 10996 2803 11003 2893
rect 11016 2827 11023 2983
rect 11036 2887 11043 3393
rect 11076 3307 11083 3393
rect 11096 3267 11103 3293
rect 10996 2796 11023 2803
rect 11016 2776 11023 2796
rect 11056 2788 11063 3133
rect 11076 2986 11083 3193
rect 10996 2687 11003 2743
rect 11036 2740 11043 2743
rect 11033 2727 11047 2740
rect 10956 2476 10963 2653
rect 10996 2587 11003 2633
rect 10916 2436 10943 2443
rect 10916 2327 10923 2436
rect 10916 1807 10923 2292
rect 10936 1883 10943 2373
rect 10956 2167 10963 2413
rect 10976 2347 10983 2443
rect 11016 2427 11023 2613
rect 11036 2387 11043 2473
rect 11056 2256 11063 2673
rect 11076 2587 11083 2733
rect 11076 2427 11083 2573
rect 11096 2327 11103 3053
rect 11116 2443 11123 3393
rect 11136 2487 11143 3333
rect 11176 3327 11183 3533
rect 11196 3407 11203 3453
rect 11216 3347 11223 3493
rect 11276 3483 11283 4673
rect 11296 3507 11303 4553
rect 11336 4443 11343 5733
rect 11316 4436 11343 4443
rect 11316 3507 11323 4436
rect 11276 3476 11323 3483
rect 11167 3303 11180 3307
rect 11167 3296 11183 3303
rect 11167 3293 11180 3296
rect 11196 3247 11203 3263
rect 11236 3260 11243 3263
rect 11233 3247 11247 3260
rect 11207 3236 11223 3243
rect 11156 2627 11163 3213
rect 11176 2547 11183 3013
rect 11216 3003 11223 3236
rect 11256 3027 11263 3253
rect 11196 2996 11223 3003
rect 11196 2927 11203 2996
rect 11196 2527 11203 2873
rect 11256 2807 11263 2963
rect 11276 2887 11283 3447
rect 11296 3287 11303 3413
rect 11213 2787 11227 2793
rect 11276 2783 11283 2813
rect 11256 2776 11283 2783
rect 11116 2436 11143 2443
rect 10976 2207 10983 2254
rect 10996 1968 11003 2212
rect 11076 2187 11083 2223
rect 11016 1926 11023 1993
rect 10936 1876 10963 1883
rect 10916 1683 10923 1734
rect 10936 1703 10943 1853
rect 10956 1787 10963 1876
rect 10936 1696 10963 1703
rect 11016 1696 11043 1703
rect 10916 1676 10943 1683
rect 10896 1436 10923 1443
rect 10776 1403 10783 1434
rect 10776 1396 10803 1403
rect 10736 1216 10743 1293
rect 10756 1176 10783 1183
rect 10736 916 10743 1133
rect 10716 787 10723 883
rect 10696 387 10703 613
rect 10716 547 10723 773
rect 10776 763 10783 1176
rect 10796 1147 10803 1396
rect 10816 1187 10823 1353
rect 10856 1347 10863 1403
rect 10836 807 10843 913
rect 10856 847 10863 973
rect 10767 756 10783 763
rect 10756 696 10763 753
rect 10876 687 10883 1373
rect 10896 1167 10903 1333
rect 10916 1007 10923 1436
rect 10936 1387 10943 1676
rect 10956 1347 10963 1453
rect 10973 920 10987 933
rect 10976 916 10983 920
rect 10916 847 10923 883
rect 10956 807 10963 883
rect 10996 696 11003 873
rect 11016 867 11023 1673
rect 11036 1647 11043 1696
rect 11056 1436 11063 1734
rect 11076 1706 11083 1993
rect 11076 1567 11083 1692
rect 11096 1587 11103 2193
rect 11116 1867 11123 1893
rect 11136 1887 11143 2436
rect 11156 2367 11163 2443
rect 11196 2423 11203 2443
rect 11196 2416 11223 2423
rect 11156 2207 11163 2313
rect 11176 2268 11183 2413
rect 11176 2007 11183 2254
rect 11196 2167 11203 2393
rect 11216 2367 11223 2416
rect 11216 1968 11223 2273
rect 11236 2227 11243 2433
rect 11256 2287 11263 2533
rect 11276 2307 11283 2513
rect 11296 2407 11303 3233
rect 11256 2007 11263 2223
rect 11076 1307 11083 1403
rect 11036 887 11043 1214
rect 11056 1187 11063 1213
rect 11056 947 11063 1152
rect 11056 747 11063 933
rect 10736 146 10743 593
rect 10756 367 10763 394
rect 10776 367 10783 453
rect 10813 400 10827 413
rect 10976 408 10983 652
rect 11016 507 11023 663
rect 11056 467 11063 694
rect 11076 666 11083 1173
rect 11116 923 11123 1773
rect 11136 1187 11143 1693
rect 11156 1667 11163 1913
rect 11196 1887 11203 1923
rect 11236 1867 11243 1923
rect 11216 1736 11223 1793
rect 11236 1667 11243 1703
rect 11296 1627 11303 2153
rect 11216 1387 11223 1613
rect 11256 1436 11263 1573
rect 11276 1396 11303 1403
rect 11196 1216 11203 1293
rect 11216 1180 11223 1183
rect 11213 1167 11227 1180
rect 11276 1127 11283 1373
rect 11096 916 11123 923
rect 11096 427 11103 916
rect 10816 396 10823 400
rect 11116 396 11123 733
rect 11136 627 11143 883
rect 10976 366 10983 394
rect 11076 343 11083 363
rect 11056 336 11083 343
rect 11056 247 11063 336
rect 11076 176 11083 313
rect 11136 203 11143 413
rect 11156 327 11163 853
rect 11216 696 11223 1113
rect 11296 987 11303 1396
rect 11236 627 11243 663
rect 11116 196 11143 203
rect 11116 176 11123 196
rect 10756 107 10763 143
rect 11096 47 11103 143
rect 11316 107 11323 3476
rect 11336 2367 11343 4193
rect 11336 146 11343 2293
<< m3contact >>
rect 13 11094 27 11108
rect 193 11094 207 11108
rect 333 11073 347 11087
rect 13 10893 27 10907
rect 93 10753 107 10767
rect 33 10673 47 10687
rect 153 11052 167 11066
rect 1353 11113 1367 11127
rect 853 11093 867 11107
rect 1073 11094 1087 11108
rect 1213 11093 1227 11107
rect 1313 11094 1327 11108
rect 493 11074 507 11088
rect 413 11052 427 11066
rect 273 10774 287 10788
rect 433 10814 447 10828
rect 793 11074 807 11088
rect 913 11074 927 11088
rect 613 10993 627 11007
rect 793 10993 807 11007
rect 453 10813 467 10827
rect 493 10814 507 10828
rect 173 10673 187 10687
rect 373 10673 387 10687
rect 133 10574 147 10588
rect 273 10633 287 10647
rect 193 10532 207 10546
rect 173 10274 187 10288
rect 253 10273 267 10287
rect 253 10232 267 10246
rect 213 10093 227 10107
rect 173 10054 187 10068
rect 253 10054 267 10068
rect 193 9853 207 9867
rect 133 9833 147 9847
rect 233 9793 247 9807
rect 133 9754 147 9768
rect 193 9754 207 9768
rect 253 9753 267 9767
rect 173 9712 187 9726
rect 213 9712 227 9726
rect 133 9534 147 9548
rect 173 9534 187 9548
rect 213 9534 227 9548
rect 253 9534 267 9548
rect 93 9433 107 9447
rect 73 5993 87 6007
rect 13 5793 27 5807
rect 113 9213 127 9227
rect 173 9253 187 9267
rect 213 9153 227 9167
rect 153 9014 167 9028
rect 213 9013 227 9027
rect 413 10774 427 10788
rect 473 10673 487 10687
rect 413 10633 427 10647
rect 333 10593 347 10607
rect 393 10593 407 10607
rect 313 10113 327 10127
rect 293 9853 307 9867
rect 373 10574 387 10588
rect 393 10532 407 10546
rect 433 10532 447 10546
rect 473 10532 487 10546
rect 553 10774 567 10788
rect 653 10774 667 10788
rect 553 10673 567 10687
rect 633 10673 647 10687
rect 573 10613 587 10627
rect 833 10753 847 10767
rect 833 10653 847 10667
rect 573 10532 587 10546
rect 613 10532 627 10546
rect 713 10533 727 10547
rect 533 10393 547 10407
rect 633 10393 647 10407
rect 393 10313 407 10327
rect 633 10313 647 10327
rect 493 10274 507 10288
rect 593 10274 607 10288
rect 373 10232 387 10246
rect 453 10113 467 10127
rect 413 10054 427 10068
rect 613 10232 627 10246
rect 713 10274 727 10288
rect 713 10233 727 10247
rect 673 10193 687 10207
rect 493 10093 507 10107
rect 513 10054 527 10068
rect 573 10054 587 10068
rect 653 10054 667 10068
rect 353 9713 367 9727
rect 313 9693 327 9707
rect 293 9553 307 9567
rect 433 10012 447 10026
rect 493 10012 507 10026
rect 513 9993 527 10007
rect 553 9873 567 9887
rect 413 9833 427 9847
rect 513 9833 527 9847
rect 473 9712 487 9726
rect 433 9693 447 9707
rect 393 9553 407 9567
rect 373 9533 387 9547
rect 433 9534 447 9548
rect 493 9533 507 9547
rect 333 9493 347 9507
rect 453 9492 467 9506
rect 513 9492 527 9506
rect 413 9234 427 9248
rect 453 9234 467 9248
rect 493 9234 507 9248
rect 333 9192 347 9206
rect 393 9192 407 9206
rect 313 9093 327 9107
rect 433 9093 447 9107
rect 233 8993 247 9007
rect 113 8973 127 8987
rect 113 8433 127 8447
rect 173 8972 187 8986
rect 233 8953 247 8967
rect 213 8913 227 8927
rect 173 8753 187 8767
rect 153 8714 167 8728
rect 213 8713 227 8727
rect 193 8573 207 8587
rect 233 8493 247 8507
rect 233 8333 247 8347
rect 273 8994 287 9008
rect 313 8992 327 9006
rect 453 8992 467 9006
rect 293 8953 307 8967
rect 633 9993 647 10007
rect 853 10613 867 10627
rect 1113 11052 1127 11066
rect 1053 11033 1067 11047
rect 1093 10993 1107 11007
rect 1033 10814 1047 10828
rect 1513 11093 1527 11107
rect 1553 11094 1567 11108
rect 1293 11052 1307 11066
rect 1333 11052 1347 11066
rect 1393 11053 1407 11067
rect 1213 10873 1227 10887
rect 1153 10814 1167 10828
rect 1053 10773 1067 10787
rect 1193 10772 1207 10786
rect 1313 10774 1327 10788
rect 1593 11052 1607 11066
rect 1533 11033 1547 11047
rect 1793 11133 1807 11147
rect 1913 11133 1927 11147
rect 1833 11113 1847 11127
rect 1873 11113 1887 11127
rect 1773 11052 1787 11066
rect 1733 10993 1747 11007
rect 1813 10993 1827 11007
rect 1733 10953 1747 10967
rect 1733 10893 1747 10907
rect 1533 10853 1547 10867
rect 1113 10733 1127 10747
rect 1213 10733 1227 10747
rect 1033 10693 1047 10707
rect 1213 10693 1227 10707
rect 913 10653 927 10667
rect 893 10573 907 10587
rect 833 10532 847 10546
rect 873 10532 887 10546
rect 913 10473 927 10487
rect 873 10433 887 10447
rect 833 10333 847 10347
rect 793 10274 807 10288
rect 893 10232 907 10246
rect 853 10193 867 10207
rect 813 10113 827 10127
rect 853 10054 867 10068
rect 833 9873 847 9887
rect 773 9813 787 9827
rect 573 9793 587 9807
rect 593 9774 607 9788
rect 753 9774 767 9788
rect 1513 10772 1527 10786
rect 1553 10772 1567 10786
rect 1673 10753 1687 10767
rect 1793 10813 1807 10827
rect 1273 10653 1287 10667
rect 1493 10653 1507 10667
rect 1213 10473 1227 10487
rect 1213 10433 1227 10447
rect 1073 10353 1087 10367
rect 1073 10313 1087 10327
rect 1113 10274 1127 10288
rect 1193 10274 1207 10288
rect 1093 10232 1107 10246
rect 1133 10232 1147 10246
rect 1193 10233 1207 10247
rect 1033 10093 1047 10107
rect 1113 10213 1127 10227
rect 1093 10113 1107 10127
rect 1233 10413 1247 10427
rect 1213 10173 1227 10187
rect 1233 10113 1247 10127
rect 1113 10093 1127 10107
rect 1193 10093 1207 10107
rect 1173 10054 1187 10068
rect 1213 9993 1227 10007
rect 1113 9813 1127 9827
rect 573 9613 587 9627
rect 573 9353 587 9367
rect 913 9773 927 9787
rect 713 9754 727 9768
rect 893 9753 907 9767
rect 633 9713 647 9727
rect 653 9693 667 9707
rect 693 9693 707 9707
rect 773 9534 787 9548
rect 633 9433 647 9447
rect 673 9393 687 9407
rect 773 9393 787 9407
rect 1093 9713 1107 9727
rect 953 9633 967 9647
rect 873 9613 887 9627
rect 833 9534 847 9548
rect 893 9492 907 9506
rect 853 9453 867 9467
rect 1053 9534 1067 9548
rect 973 9453 987 9467
rect 953 9433 967 9447
rect 813 9353 827 9367
rect 853 9273 867 9287
rect 633 9231 647 9245
rect 773 9233 787 9247
rect 893 9234 907 9248
rect 593 9133 607 9147
rect 653 9133 667 9147
rect 673 9113 687 9127
rect 753 9053 767 9067
rect 733 9014 747 9028
rect 613 8952 627 8966
rect 653 8953 667 8967
rect 513 8833 527 8847
rect 553 8833 567 8847
rect 333 8753 347 8767
rect 453 8753 467 8767
rect 293 8633 307 8647
rect 373 8714 387 8728
rect 353 8593 367 8607
rect 413 8593 427 8607
rect 333 8533 347 8547
rect 133 8073 147 8087
rect 213 8152 227 8166
rect 173 8053 187 8067
rect 213 8033 227 8047
rect 173 7932 187 7946
rect 113 7813 127 7827
rect 453 8533 467 8547
rect 413 8494 427 8508
rect 313 8313 327 8327
rect 353 8313 367 8327
rect 293 8152 307 8166
rect 273 7773 287 7787
rect 193 7733 207 7747
rect 253 7673 267 7687
rect 213 7632 227 7646
rect 253 7632 267 7646
rect 173 7454 187 7468
rect 253 7454 267 7468
rect 193 7412 207 7426
rect 153 7154 167 7168
rect 193 7154 207 7168
rect 133 6953 147 6967
rect 173 6953 187 6967
rect 193 6934 207 6948
rect 233 6933 247 6947
rect 273 7273 287 7287
rect 273 7154 287 7168
rect 293 6993 307 7007
rect 273 6953 287 6967
rect 253 6913 267 6927
rect 213 6893 227 6907
rect 213 6773 227 6787
rect 133 6634 147 6648
rect 233 6634 247 6648
rect 213 6592 227 6606
rect 173 6553 187 6567
rect 253 6553 267 6567
rect 433 8433 447 8447
rect 493 8293 507 8307
rect 373 8273 387 8287
rect 413 8273 427 8287
rect 433 8194 447 8208
rect 453 8152 467 8166
rect 413 8133 427 8147
rect 393 8073 407 8087
rect 353 7974 367 7988
rect 433 7974 447 7988
rect 333 7632 347 7646
rect 733 8913 747 8927
rect 613 8753 627 8767
rect 913 9192 927 9206
rect 873 9153 887 9167
rect 813 9014 827 9028
rect 833 8972 847 8986
rect 773 8733 787 8747
rect 813 8733 827 8747
rect 613 8694 627 8708
rect 753 8694 767 8708
rect 793 8633 807 8647
rect 673 8573 687 8587
rect 633 8533 647 8547
rect 773 8533 787 8547
rect 773 8473 787 8487
rect 653 8413 667 8427
rect 693 8313 707 8327
rect 533 8293 547 8307
rect 513 7953 527 7967
rect 653 8194 667 8208
rect 693 8194 707 8208
rect 553 8152 567 8166
rect 673 8133 687 8147
rect 633 8053 647 8067
rect 553 8033 567 8047
rect 413 7932 427 7946
rect 413 7753 427 7767
rect 493 7893 507 7907
rect 493 7753 507 7767
rect 453 7733 467 7747
rect 433 7674 447 7688
rect 413 7632 427 7646
rect 353 7593 367 7607
rect 393 7493 407 7507
rect 413 7493 427 7507
rect 473 7593 487 7607
rect 453 7454 467 7468
rect 333 7413 347 7427
rect 373 7412 387 7426
rect 413 7412 427 7426
rect 653 7952 667 7966
rect 853 8673 867 8687
rect 873 8613 887 8627
rect 893 8452 907 8466
rect 1013 9393 1027 9407
rect 1013 9333 1027 9347
rect 993 9313 1007 9327
rect 1133 9533 1147 9547
rect 1133 9492 1147 9506
rect 1113 9473 1127 9487
rect 1153 9393 1167 9407
rect 1113 9273 1127 9287
rect 1013 9192 1027 9206
rect 1053 9192 1067 9206
rect 1093 9192 1107 9206
rect 1153 9193 1167 9207
rect 1133 9093 1147 9107
rect 1093 9053 1107 9067
rect 1053 9014 1067 9028
rect 1133 9033 1147 9047
rect 1073 8972 1087 8986
rect 1033 8933 1047 8947
rect 1073 8933 1087 8947
rect 1133 8933 1147 8947
rect 1033 8713 1047 8727
rect 1073 8672 1087 8686
rect 993 8593 1007 8607
rect 1073 8553 1087 8567
rect 993 8494 1007 8508
rect 1073 8494 1087 8508
rect 1113 8494 1127 8508
rect 1213 9753 1227 9767
rect 1373 10473 1387 10487
rect 1333 10433 1347 10447
rect 1533 10552 1547 10566
rect 1533 10353 1547 10367
rect 1293 10274 1307 10288
rect 1353 10193 1367 10207
rect 1353 10172 1367 10186
rect 1513 10213 1527 10227
rect 1473 10193 1487 10207
rect 1413 10133 1427 10147
rect 1473 10013 1487 10027
rect 1273 9713 1287 9727
rect 1373 9753 1387 9767
rect 1413 9754 1427 9768
rect 1453 9754 1467 9768
rect 1313 9712 1327 9726
rect 1353 9712 1367 9726
rect 1233 9673 1247 9687
rect 1293 9653 1307 9667
rect 1253 9534 1267 9548
rect 1453 9713 1467 9727
rect 1393 9673 1407 9687
rect 1353 9613 1367 9627
rect 1453 9573 1467 9587
rect 1213 9453 1227 9467
rect 1173 8633 1187 8647
rect 993 8453 1007 8467
rect 1093 8452 1107 8466
rect 1153 8453 1167 8467
rect 1313 9492 1327 9506
rect 1353 9473 1367 9487
rect 1233 9413 1247 9427
rect 1273 9413 1287 9427
rect 1353 9234 1367 9248
rect 1273 9193 1287 9207
rect 1433 9254 1447 9268
rect 1373 9192 1387 9206
rect 1413 9192 1427 9206
rect 1333 9113 1347 9127
rect 1313 9093 1327 9107
rect 1273 9033 1287 9047
rect 1333 9053 1347 9067
rect 1413 9013 1427 9027
rect 1233 8833 1247 8847
rect 1333 8933 1347 8947
rect 1373 8873 1387 8887
rect 1313 8853 1327 8867
rect 1293 8773 1307 8787
rect 1633 10274 1647 10288
rect 1713 10653 1727 10667
rect 1693 10613 1707 10627
rect 1693 10552 1707 10566
rect 1793 10493 1807 10507
rect 1773 10433 1787 10447
rect 1873 10333 1887 10347
rect 1773 10293 1787 10307
rect 1813 10293 1827 10307
rect 1673 10273 1687 10287
rect 1573 10213 1587 10227
rect 1533 10193 1547 10207
rect 1613 10193 1627 10207
rect 1553 10173 1567 10187
rect 1573 10012 1587 10026
rect 1613 9754 1627 9768
rect 2053 11094 2067 11108
rect 2093 11094 2107 11108
rect 1933 10853 1947 10867
rect 1973 10853 1987 10867
rect 2013 10794 2027 10808
rect 1993 10633 2007 10647
rect 2073 10633 2087 10647
rect 1993 10612 2007 10626
rect 2033 10613 2047 10627
rect 1953 10574 1967 10588
rect 1973 10532 1987 10546
rect 2013 10532 2027 10546
rect 2073 10532 2087 10546
rect 2033 10274 2047 10288
rect 1833 10232 1847 10246
rect 1913 10232 1927 10246
rect 2053 10232 2067 10246
rect 1773 10173 1787 10187
rect 2053 10153 2067 10167
rect 1793 10133 1807 10147
rect 1713 10054 1727 10068
rect 1753 10054 1767 10068
rect 1853 10093 1867 10107
rect 2053 10093 2067 10107
rect 1993 10073 2007 10087
rect 1913 10053 1927 10067
rect 1993 10054 2007 10068
rect 1853 10033 1867 10047
rect 1713 10013 1727 10027
rect 1773 9993 1787 10007
rect 1813 9993 1827 10007
rect 1873 9933 1887 9947
rect 1713 9853 1727 9867
rect 1593 9712 1607 9726
rect 1633 9653 1647 9667
rect 1513 9633 1527 9647
rect 1553 9573 1567 9587
rect 1513 9534 1527 9548
rect 1633 9533 1647 9547
rect 1753 9754 1767 9768
rect 1833 9754 1847 9768
rect 1773 9712 1787 9726
rect 1813 9712 1827 9726
rect 1753 9593 1767 9607
rect 1733 9573 1747 9587
rect 1693 9492 1707 9506
rect 1793 9492 1807 9506
rect 1873 9473 1887 9487
rect 1533 9453 1547 9467
rect 1753 9453 1767 9467
rect 1473 9393 1487 9407
rect 1553 9333 1567 9347
rect 2053 10033 2067 10047
rect 1973 9993 1987 10007
rect 1933 9753 1947 9767
rect 1933 9712 1947 9726
rect 2033 9793 2047 9807
rect 2033 9754 2047 9768
rect 2013 9712 2027 9726
rect 2093 9713 2107 9727
rect 2053 9673 2067 9687
rect 2013 9534 2027 9548
rect 2093 9534 2107 9548
rect 1993 9333 2007 9347
rect 1913 9313 1927 9327
rect 2073 9453 2087 9467
rect 1913 9273 1927 9287
rect 2033 9273 2047 9287
rect 1613 9254 1627 9268
rect 1513 9213 1527 9227
rect 1653 9212 1667 9226
rect 1773 9214 1787 9228
rect 1913 9214 1927 9228
rect 1473 9173 1487 9187
rect 1573 9173 1587 9187
rect 1673 9173 1687 9187
rect 1573 9133 1587 9147
rect 1553 9053 1567 9067
rect 1453 9013 1467 9027
rect 1533 8972 1547 8986
rect 1433 8853 1447 8867
rect 1373 8773 1387 8787
rect 1233 8734 1247 8748
rect 1313 8734 1327 8748
rect 1353 8692 1367 8706
rect 1273 8653 1287 8667
rect 1473 8733 1487 8747
rect 1773 9073 1787 9087
rect 1873 9033 1887 9047
rect 1853 9014 1867 9028
rect 1753 8972 1767 8986
rect 1833 8933 1847 8947
rect 1793 8853 1807 8867
rect 1693 8733 1707 8747
rect 1773 8733 1787 8747
rect 1633 8653 1647 8667
rect 1353 8573 1367 8587
rect 1313 8494 1327 8508
rect 973 8433 987 8447
rect 1213 8433 1227 8447
rect 813 8413 827 8427
rect 1533 8573 1547 8587
rect 1433 8533 1447 8547
rect 1453 8494 1467 8508
rect 1573 8494 1587 8508
rect 1433 8473 1447 8487
rect 1373 8433 1387 8447
rect 1293 8393 1307 8407
rect 1293 8353 1307 8367
rect 1333 8353 1347 8367
rect 953 8333 967 8347
rect 813 8233 827 8247
rect 893 8194 907 8208
rect 933 8193 947 8207
rect 873 8093 887 8107
rect 893 8093 907 8107
rect 853 8073 867 8087
rect 853 7973 867 7987
rect 1093 8313 1107 8327
rect 1293 8194 1307 8208
rect 1073 8152 1087 8166
rect 1313 8152 1327 8166
rect 953 8113 967 8127
rect 1273 8113 1287 8127
rect 1353 8073 1367 8087
rect 1253 7993 1267 8007
rect 793 7913 807 7927
rect 853 7913 867 7927
rect 893 7813 907 7827
rect 953 7893 967 7907
rect 913 7793 927 7807
rect 633 7753 647 7767
rect 893 7753 907 7767
rect 673 7733 687 7747
rect 873 7674 887 7688
rect 553 7593 567 7607
rect 853 7632 867 7646
rect 653 7553 667 7567
rect 773 7513 787 7527
rect 573 7493 587 7507
rect 593 7454 607 7468
rect 633 7454 647 7468
rect 493 7412 507 7426
rect 613 7412 627 7426
rect 473 7353 487 7367
rect 333 7313 347 7327
rect 313 6913 327 6927
rect 373 7213 387 7227
rect 413 7053 427 7067
rect 593 7393 607 7407
rect 653 7273 667 7287
rect 593 7193 607 7207
rect 653 7193 667 7207
rect 613 7154 627 7168
rect 673 7154 687 7168
rect 493 7033 507 7047
rect 633 7112 647 7126
rect 673 7033 687 7047
rect 593 6953 607 6967
rect 333 6893 347 6907
rect 473 6893 487 6907
rect 313 6873 327 6887
rect 213 6433 227 6447
rect 493 6773 507 6787
rect 373 6633 387 6647
rect 433 6634 447 6648
rect 333 6613 347 6627
rect 353 6473 367 6487
rect 333 6453 347 6467
rect 313 6433 327 6447
rect 253 6373 267 6387
rect 173 6313 187 6327
rect 233 6253 247 6267
rect 173 6114 187 6128
rect 333 6313 347 6327
rect 313 6213 327 6227
rect 633 6733 647 6747
rect 753 7013 767 7027
rect 693 6993 707 7007
rect 813 7493 827 7507
rect 853 7454 867 7468
rect 893 7454 907 7468
rect 833 7412 847 7426
rect 1113 7952 1127 7966
rect 1313 7913 1327 7927
rect 1313 7833 1327 7847
rect 1273 7713 1287 7727
rect 973 7674 987 7688
rect 973 7633 987 7647
rect 973 7553 987 7567
rect 953 7413 967 7427
rect 973 7373 987 7387
rect 893 7333 907 7347
rect 793 7153 807 7167
rect 793 7113 807 7127
rect 853 7112 867 7126
rect 893 7113 907 7127
rect 793 7053 807 7067
rect 793 6993 807 7007
rect 773 6934 787 6948
rect 833 6934 847 6948
rect 693 6853 707 6867
rect 533 6633 547 6647
rect 633 6634 647 6648
rect 693 6634 707 6648
rect 413 6592 427 6606
rect 453 6592 467 6606
rect 493 6593 507 6607
rect 413 6473 427 6487
rect 373 6414 387 6428
rect 453 6414 467 6428
rect 393 6372 407 6386
rect 513 6372 527 6386
rect 433 6153 447 6167
rect 353 6114 367 6128
rect 393 6114 407 6128
rect 853 6892 867 6906
rect 973 7033 987 7047
rect 973 6893 987 6907
rect 1033 7674 1047 7688
rect 1313 7674 1327 7688
rect 1033 7513 1047 7527
rect 1333 7632 1347 7646
rect 1293 7593 1307 7607
rect 1393 8412 1407 8426
rect 1093 7573 1107 7587
rect 1373 7573 1387 7587
rect 1353 7533 1367 7547
rect 1053 7493 1067 7507
rect 1233 7493 1247 7507
rect 1033 7473 1047 7487
rect 1073 7454 1087 7468
rect 1113 7454 1127 7468
rect 1293 7413 1307 7427
rect 1113 7393 1127 7407
rect 1253 7393 1267 7407
rect 1053 7353 1067 7367
rect 1233 7213 1247 7227
rect 1133 7153 1147 7167
rect 1613 8493 1627 8507
rect 1553 8452 1567 8466
rect 1713 8653 1727 8667
rect 1653 8633 1667 8647
rect 1733 8494 1747 8508
rect 1793 8573 1807 8587
rect 1753 8452 1767 8466
rect 1633 8413 1647 8427
rect 1613 8393 1627 8407
rect 1453 8353 1467 8367
rect 1433 8233 1447 8247
rect 1413 8194 1427 8208
rect 1413 7873 1427 7887
rect 1953 9173 1967 9187
rect 2053 9133 2067 9147
rect 2013 9113 2027 9127
rect 1993 9033 2007 9047
rect 2053 9033 2067 9047
rect 2033 9014 2047 9028
rect 2013 8972 2027 8986
rect 2073 8973 2087 8987
rect 1913 8933 1927 8947
rect 1973 8933 1987 8947
rect 1913 8853 1927 8867
rect 1933 8653 1947 8667
rect 1873 8633 1887 8647
rect 1833 8393 1847 8407
rect 1653 8273 1667 8287
rect 1793 8273 1807 8287
rect 1473 8233 1487 8247
rect 1473 8192 1487 8206
rect 1513 8194 1527 8208
rect 1853 8233 1867 8247
rect 1753 8194 1767 8208
rect 1793 8194 1807 8208
rect 1473 8113 1487 8127
rect 1753 8133 1767 8147
rect 1793 8133 1807 8147
rect 1653 8113 1667 8127
rect 1733 8113 1747 8127
rect 1533 8073 1547 8087
rect 1513 8033 1527 8047
rect 1473 7974 1487 7988
rect 1453 7913 1467 7927
rect 1433 7674 1447 7688
rect 1693 8053 1707 8067
rect 1593 7993 1607 8007
rect 1653 7993 1667 8007
rect 1553 7974 1567 7988
rect 1613 7932 1627 7946
rect 1573 7913 1587 7927
rect 1553 7753 1567 7767
rect 1573 7693 1587 7707
rect 1613 7693 1627 7707
rect 1433 7533 1447 7547
rect 1573 7632 1587 7646
rect 1573 7513 1587 7527
rect 1533 7493 1547 7507
rect 1393 7473 1407 7487
rect 1373 7293 1387 7307
rect 1313 7273 1327 7287
rect 1353 7273 1367 7287
rect 1313 7233 1327 7247
rect 1293 7174 1307 7188
rect 1353 7174 1367 7188
rect 1253 7132 1267 7146
rect 1253 7073 1267 7087
rect 1233 7033 1247 7047
rect 1033 6953 1047 6967
rect 1313 7053 1327 7067
rect 1273 7033 1287 7047
rect 1073 6934 1087 6948
rect 1113 6934 1127 6948
rect 1253 6934 1267 6948
rect 1013 6893 1027 6907
rect 833 6853 847 6867
rect 953 6853 967 6867
rect 993 6853 1007 6867
rect 973 6753 987 6767
rect 1013 6753 1027 6767
rect 653 6592 667 6606
rect 653 6533 667 6547
rect 733 6513 747 6527
rect 653 6453 667 6467
rect 573 6414 587 6428
rect 613 6414 627 6428
rect 633 6372 647 6386
rect 573 6313 587 6327
rect 573 6253 587 6267
rect 633 6153 647 6167
rect 733 6193 747 6207
rect 693 6133 707 6147
rect 453 6053 467 6067
rect 513 6053 527 6067
rect 593 5993 607 6007
rect 93 5733 107 5747
rect 33 5473 47 5487
rect 313 5973 327 5987
rect 413 5973 427 5987
rect 213 5933 227 5947
rect 293 5893 307 5907
rect 553 5893 567 5907
rect 313 5872 327 5886
rect 413 5872 427 5886
rect 173 5852 187 5866
rect 253 5832 267 5846
rect 413 5833 427 5847
rect 373 5733 387 5747
rect 273 5613 287 5627
rect 173 5473 187 5487
rect 353 5374 367 5388
rect 693 6053 707 6067
rect 653 5874 667 5888
rect 593 5793 607 5807
rect 393 5572 407 5586
rect 553 5573 567 5587
rect 413 5533 427 5547
rect 633 5613 647 5627
rect 653 5533 667 5547
rect 673 5413 687 5427
rect 453 5374 467 5388
rect 593 5374 607 5388
rect 673 5374 687 5388
rect 213 5332 227 5346
rect 153 5313 167 5327
rect 193 5173 207 5187
rect 253 5093 267 5107
rect 333 5093 347 5107
rect 293 5032 307 5046
rect 133 4973 147 4987
rect 173 4933 187 4947
rect 293 4873 307 4887
rect 193 4812 207 4826
rect 293 4812 307 4826
rect 233 4673 247 4687
rect 273 4633 287 4647
rect 193 4573 207 4587
rect 133 4512 147 4526
rect 173 4512 187 4526
rect 73 3772 87 3786
rect 213 4413 227 4427
rect 213 4373 227 4387
rect 213 4253 227 4267
rect 153 4233 167 4247
rect 193 4233 207 4247
rect 213 3933 227 3947
rect 233 3814 247 3828
rect 213 3772 227 3786
rect 273 3773 287 3787
rect 173 3713 187 3727
rect 273 3633 287 3647
rect 233 3593 247 3607
rect 193 3514 207 3528
rect 133 3473 147 3487
rect 173 3472 187 3486
rect 253 3473 267 3487
rect 213 3373 227 3387
rect 173 3294 187 3308
rect 213 3294 227 3308
rect 273 3294 287 3308
rect 193 3252 207 3266
rect 253 3253 267 3267
rect 173 3233 187 3247
rect 233 3113 247 3127
rect 193 2893 207 2907
rect 133 2833 147 2847
rect 113 2433 127 2447
rect 173 2793 187 2807
rect 233 2793 247 2807
rect 213 2774 227 2788
rect 233 2732 247 2746
rect 273 2633 287 2647
rect 173 2474 187 2488
rect 193 2432 207 2446
rect 193 2293 207 2307
rect 173 2273 187 2287
rect 213 2254 227 2268
rect 253 2254 267 2268
rect 133 2213 147 2227
rect 193 2212 207 2226
rect 273 2093 287 2107
rect 193 2073 207 2087
rect 253 2073 267 2087
rect 173 1912 187 1926
rect 253 1912 267 1926
rect 193 1773 207 1787
rect 213 1692 227 1706
rect 313 4713 327 4727
rect 393 5332 407 5346
rect 433 5293 447 5307
rect 453 5113 467 5127
rect 513 5074 527 5088
rect 553 5074 567 5088
rect 533 5032 547 5046
rect 493 4973 507 4987
rect 573 4893 587 4907
rect 413 4812 427 4826
rect 573 4812 587 4826
rect 353 4773 367 4787
rect 413 4773 427 4787
rect 633 5313 647 5327
rect 693 5313 707 5327
rect 633 5273 647 5287
rect 613 5074 627 5088
rect 613 4953 627 4967
rect 693 5133 707 5147
rect 633 4854 647 4868
rect 653 4812 667 4826
rect 593 4713 607 4727
rect 413 4593 427 4607
rect 373 4573 387 4587
rect 533 4554 547 4568
rect 613 4554 627 4568
rect 793 6612 807 6626
rect 833 6613 847 6627
rect 773 6513 787 6527
rect 753 5793 767 5807
rect 853 6513 867 6527
rect 993 6513 1007 6527
rect 793 6453 807 6467
rect 973 6493 987 6507
rect 1093 6873 1107 6887
rect 1293 6873 1307 6887
rect 1173 6853 1187 6867
rect 1133 6733 1147 6747
rect 1133 6654 1147 6668
rect 1093 6612 1107 6626
rect 1093 6533 1107 6547
rect 1073 6493 1087 6507
rect 1033 6433 1047 6447
rect 1193 6653 1207 6667
rect 1173 6513 1187 6527
rect 1173 6394 1187 6408
rect 1053 6372 1067 6386
rect 1333 6654 1347 6668
rect 1373 7133 1387 7147
rect 1493 7454 1507 7468
rect 1433 7393 1447 7407
rect 1473 7373 1487 7387
rect 1513 7373 1527 7387
rect 1413 7293 1427 7307
rect 1393 7112 1407 7126
rect 1273 6613 1287 6627
rect 1433 7273 1447 7287
rect 1533 7253 1547 7267
rect 1553 7233 1567 7247
rect 1513 7193 1527 7207
rect 1493 7112 1507 7126
rect 1533 7073 1547 7087
rect 1493 7013 1507 7027
rect 1453 6993 1467 7007
rect 1453 6933 1467 6947
rect 1533 6934 1547 6948
rect 1433 6873 1447 6887
rect 1373 6592 1387 6606
rect 1413 6592 1427 6606
rect 1272 6393 1286 6407
rect 1133 6352 1147 6366
rect 1193 6352 1207 6366
rect 1293 6392 1307 6406
rect 1033 6313 1047 6327
rect 1093 6313 1107 6327
rect 993 6293 1007 6307
rect 833 6193 847 6207
rect 973 6193 987 6207
rect 813 6153 827 6167
rect 793 5993 807 6007
rect 833 6133 847 6147
rect 893 6114 907 6128
rect 1013 6114 1027 6128
rect 813 5973 827 5987
rect 853 5953 867 5967
rect 913 5953 927 5967
rect 793 5894 807 5908
rect 873 5894 887 5908
rect 953 5894 967 5908
rect 773 5594 787 5608
rect 753 5533 767 5547
rect 853 5852 867 5866
rect 833 5594 847 5608
rect 973 5813 987 5827
rect 893 5552 907 5566
rect 953 5553 967 5567
rect 813 5473 827 5487
rect 853 5473 867 5487
rect 753 5433 767 5447
rect 873 5453 887 5467
rect 813 5333 827 5347
rect 733 5133 747 5147
rect 713 5073 727 5087
rect 853 5332 867 5346
rect 853 5213 867 5227
rect 813 5032 827 5046
rect 773 4993 787 5007
rect 733 4973 747 4987
rect 773 4953 787 4967
rect 713 4853 727 4867
rect 693 4553 707 4567
rect 433 4512 447 4526
rect 533 4513 547 4527
rect 633 4512 647 4526
rect 533 4453 547 4467
rect 673 4453 687 4467
rect 393 4413 407 4427
rect 373 4333 387 4347
rect 433 4334 447 4348
rect 513 4313 527 4327
rect 373 4293 387 4307
rect 413 4253 427 4267
rect 513 4253 527 4267
rect 453 4233 467 4247
rect 413 4193 427 4207
rect 373 4033 387 4047
rect 373 3993 387 4007
rect 333 3973 347 3987
rect 353 3513 367 3527
rect 433 3973 447 3987
rect 393 3893 407 3907
rect 513 3893 527 3907
rect 473 3833 487 3847
rect 413 3713 427 3727
rect 513 3633 527 3647
rect 673 4373 687 4387
rect 673 4334 687 4348
rect 693 4292 707 4306
rect 633 4253 647 4267
rect 593 4073 607 4087
rect 553 4034 567 4048
rect 633 4034 647 4048
rect 693 4013 707 4027
rect 553 3827 567 3828
rect 553 3814 567 3827
rect 653 3992 667 4006
rect 613 3953 627 3967
rect 593 3933 607 3947
rect 633 3933 647 3947
rect 613 3873 627 3887
rect 593 3833 607 3847
rect 573 3733 587 3747
rect 553 3673 567 3687
rect 473 3593 487 3607
rect 453 3553 467 3567
rect 413 3514 427 3528
rect 433 3472 447 3486
rect 373 3293 387 3307
rect 413 3294 427 3308
rect 453 3294 467 3308
rect 393 3233 407 3247
rect 433 3233 447 3247
rect 333 3053 347 3067
rect 313 2633 327 2647
rect 573 3553 587 3567
rect 533 3294 547 3308
rect 533 3253 547 3267
rect 513 3233 527 3247
rect 693 3933 707 3947
rect 733 4553 747 4567
rect 733 4512 747 4526
rect 753 4493 767 4507
rect 733 4334 747 4348
rect 733 4113 747 4127
rect 993 5773 1007 5787
rect 1113 6293 1127 6307
rect 1073 6114 1087 6128
rect 1273 6273 1287 6287
rect 1193 6153 1207 6167
rect 1033 6093 1047 6107
rect 1093 5953 1107 5967
rect 1113 5894 1127 5908
rect 1173 5893 1187 5907
rect 1093 5793 1107 5807
rect 1153 5733 1167 5747
rect 1153 5673 1167 5687
rect 1053 5633 1067 5647
rect 1073 5552 1087 5566
rect 1053 5533 1067 5547
rect 1133 5553 1147 5567
rect 1033 5393 1047 5407
rect 1013 5333 1027 5347
rect 993 5273 1007 5287
rect 1033 5213 1047 5227
rect 973 5173 987 5187
rect 1033 5173 1047 5187
rect 913 5113 927 5127
rect 953 5113 967 5127
rect 893 4893 907 4907
rect 993 5074 1007 5088
rect 973 5032 987 5046
rect 913 4853 927 4867
rect 793 4812 807 4826
rect 793 4773 807 4787
rect 773 4093 787 4107
rect 733 3992 747 4006
rect 713 3873 727 3887
rect 653 3833 667 3847
rect 733 3833 747 3847
rect 693 3814 707 3828
rect 613 3772 627 3786
rect 673 3772 687 3786
rect 713 3772 727 3786
rect 773 3773 787 3787
rect 753 3713 767 3727
rect 593 3514 607 3528
rect 653 3514 667 3528
rect 573 3213 587 3227
rect 533 3173 547 3187
rect 473 3093 487 3107
rect 373 2952 387 2966
rect 433 2952 447 2966
rect 353 2773 367 2787
rect 353 2732 367 2746
rect 413 2732 427 2746
rect 453 2713 467 2727
rect 393 2693 407 2707
rect 333 2474 347 2488
rect 433 2633 447 2647
rect 373 2432 387 2446
rect 313 2273 327 2287
rect 453 2553 467 2567
rect 513 2833 527 2847
rect 513 2713 527 2727
rect 553 3093 567 3107
rect 613 3294 627 3308
rect 593 3053 607 3067
rect 673 3472 687 3486
rect 673 3294 687 3308
rect 653 3252 667 3266
rect 713 3252 727 3266
rect 633 3113 647 3127
rect 653 3053 667 3067
rect 753 3473 767 3487
rect 753 3413 767 3427
rect 753 3252 767 3266
rect 873 4812 887 4826
rect 1033 4812 1047 4826
rect 853 4693 867 4707
rect 833 4673 847 4687
rect 813 4554 827 4568
rect 853 4593 867 4607
rect 853 4554 867 4568
rect 833 4533 847 4547
rect 873 4493 887 4507
rect 833 4373 847 4387
rect 893 4453 907 4467
rect 913 4373 927 4387
rect 953 4533 967 4547
rect 953 4473 967 4487
rect 933 4353 947 4367
rect 833 4293 847 4307
rect 893 4292 907 4306
rect 933 4292 947 4306
rect 833 4253 847 4267
rect 813 4193 827 4207
rect 933 4233 947 4247
rect 1153 5533 1167 5547
rect 1113 5493 1127 5507
rect 1093 5393 1107 5407
rect 1193 5832 1207 5846
rect 1213 5733 1227 5747
rect 1513 6873 1527 6887
rect 1553 6853 1567 6867
rect 1673 7973 1687 7987
rect 1673 7932 1687 7946
rect 1853 8153 1867 8167
rect 1813 8113 1827 8127
rect 1853 8053 1867 8067
rect 1893 8593 1907 8607
rect 1933 8593 1947 8607
rect 1813 7974 1827 7988
rect 1753 7893 1767 7907
rect 1793 7893 1807 7907
rect 1833 7892 1847 7906
rect 1713 7753 1727 7767
rect 1693 7613 1707 7627
rect 1773 7713 1787 7727
rect 1773 7613 1787 7627
rect 1753 7593 1767 7607
rect 1733 7533 1747 7547
rect 1713 7473 1727 7487
rect 1633 7453 1647 7467
rect 1693 7454 1707 7468
rect 1493 6813 1507 6827
rect 1593 6813 1607 6827
rect 1453 6592 1467 6606
rect 1573 6634 1587 6648
rect 1553 6592 1567 6606
rect 1593 6533 1607 6547
rect 1493 6473 1507 6487
rect 1473 6453 1487 6467
rect 1453 6233 1467 6247
rect 1293 6193 1307 6207
rect 1353 6193 1367 6207
rect 1433 6193 1447 6207
rect 1373 6072 1387 6086
rect 1293 6033 1307 6047
rect 1333 6033 1347 6047
rect 1433 6033 1447 6047
rect 1333 5973 1347 5987
rect 1433 5933 1447 5947
rect 1373 5894 1387 5908
rect 1413 5894 1427 5908
rect 1453 5894 1467 5908
rect 1533 6413 1547 6427
rect 1613 6413 1627 6427
rect 1653 7353 1667 7367
rect 1793 7413 1807 7427
rect 1773 7353 1787 7367
rect 1692 7253 1706 7267
rect 1713 7253 1727 7267
rect 1673 7233 1687 7247
rect 1673 7154 1687 7168
rect 1733 7213 1747 7227
rect 1773 7154 1787 7168
rect 1853 7773 1867 7787
rect 1933 8553 1947 8567
rect 1913 8494 1927 8508
rect 1953 8494 1967 8508
rect 1913 8453 1927 8467
rect 1973 8452 1987 8466
rect 1933 8273 1947 8287
rect 1973 8194 1987 8208
rect 1953 8152 1967 8166
rect 2893 11153 2907 11167
rect 3793 11153 3807 11167
rect 2273 11133 2287 11147
rect 2573 11133 2587 11147
rect 2193 11094 2207 11108
rect 2233 11094 2247 11108
rect 2353 11093 2367 11107
rect 2493 11094 2507 11108
rect 2573 11072 2587 11086
rect 2193 11033 2207 11047
rect 2293 11052 2307 11066
rect 2353 11052 2367 11066
rect 2513 11052 2527 11066
rect 2253 11013 2267 11027
rect 2313 11013 2327 11027
rect 2473 11013 2487 11027
rect 2173 10794 2187 10808
rect 2493 10794 2507 10808
rect 2313 10773 2327 10787
rect 2253 10713 2267 10727
rect 2173 10693 2187 10707
rect 2153 10573 2167 10587
rect 2233 10574 2247 10588
rect 2133 9593 2147 9607
rect 2113 9173 2127 9187
rect 2213 10493 2227 10507
rect 2273 10274 2287 10288
rect 2413 10613 2427 10627
rect 2373 10573 2387 10587
rect 2353 10393 2367 10407
rect 2333 10274 2347 10288
rect 2313 10213 2327 10227
rect 2253 10113 2267 10127
rect 2233 10093 2247 10107
rect 2213 10012 2227 10026
rect 2333 9953 2347 9967
rect 2273 9933 2287 9947
rect 2193 9793 2207 9807
rect 2233 9754 2247 9768
rect 2253 9712 2267 9726
rect 2193 9534 2207 9548
rect 2293 9633 2307 9647
rect 2273 9613 2287 9627
rect 2213 9273 2227 9287
rect 2553 10973 2567 10987
rect 2573 10973 2587 10987
rect 2553 10793 2567 10807
rect 2553 10752 2567 10766
rect 2553 10574 2567 10588
rect 2493 10533 2507 10547
rect 2533 10533 2547 10547
rect 2433 10453 2447 10467
rect 2413 10373 2427 10387
rect 2373 10173 2387 10187
rect 2373 10113 2387 10127
rect 2393 10093 2407 10107
rect 2373 10012 2387 10026
rect 2553 10453 2567 10467
rect 2493 10313 2507 10327
rect 2453 10274 2467 10288
rect 2473 10113 2487 10127
rect 2533 10113 2547 10127
rect 2493 10093 2507 10107
rect 2413 10053 2427 10067
rect 2453 10054 2467 10068
rect 2553 10054 2567 10068
rect 2433 10012 2447 10026
rect 2373 9913 2387 9927
rect 2393 9773 2407 9787
rect 2373 9673 2387 9687
rect 2353 9533 2367 9547
rect 2333 9493 2347 9507
rect 2293 9373 2307 9387
rect 2313 9333 2327 9347
rect 2153 9234 2167 9248
rect 2193 9234 2207 9248
rect 2253 9234 2267 9248
rect 2233 9193 2247 9207
rect 2213 9113 2227 9127
rect 2272 9173 2286 9187
rect 2293 9173 2307 9187
rect 2213 8933 2227 8947
rect 2133 8893 2147 8907
rect 2213 8853 2227 8867
rect 1913 8053 1927 8067
rect 2013 8053 2027 8067
rect 1993 7993 2007 8007
rect 1933 7793 1947 7807
rect 2173 8793 2187 8807
rect 2073 8714 2087 8728
rect 2133 8714 2147 8728
rect 2153 8672 2167 8686
rect 2113 8633 2127 8647
rect 2193 8613 2207 8627
rect 2193 8553 2207 8567
rect 2173 8494 2187 8508
rect 2273 8773 2287 8787
rect 2273 8713 2287 8727
rect 2273 8573 2287 8587
rect 2073 8453 2087 8467
rect 2153 8452 2167 8466
rect 2193 8393 2207 8407
rect 2353 9192 2367 9206
rect 2453 9873 2467 9887
rect 2553 9873 2567 9887
rect 2533 9813 2547 9827
rect 2493 9773 2507 9787
rect 2713 11072 2727 11086
rect 3213 11133 3227 11147
rect 3373 11133 3387 11147
rect 3473 11133 3487 11147
rect 3253 11094 3267 11108
rect 3313 11094 3327 11108
rect 2953 11074 2967 11088
rect 2993 11053 3007 11067
rect 2993 11013 3007 11027
rect 3013 10973 3027 10987
rect 2753 10933 2767 10947
rect 2673 10853 2687 10867
rect 2753 10853 2767 10867
rect 2713 10813 2727 10827
rect 2653 10752 2667 10766
rect 2693 10752 2707 10766
rect 2713 10693 2727 10707
rect 2673 10574 2687 10588
rect 2833 10813 2847 10827
rect 2953 10813 2967 10827
rect 3133 10933 3147 10947
rect 2913 10794 2927 10808
rect 3073 10794 3087 10808
rect 2893 10752 2907 10766
rect 2933 10752 2947 10766
rect 2833 10693 2847 10707
rect 2973 10693 2987 10707
rect 2753 10573 2767 10587
rect 2893 10574 2907 10588
rect 2953 10574 2967 10588
rect 2593 10533 2607 10547
rect 2653 10532 2667 10546
rect 2693 10532 2707 10546
rect 2593 10453 2607 10467
rect 2913 10532 2927 10546
rect 2753 10413 2767 10427
rect 2653 10373 2667 10387
rect 2953 10353 2967 10367
rect 2813 10313 2827 10327
rect 2633 10274 2647 10288
rect 2673 10274 2687 10288
rect 2713 10274 2727 10288
rect 2773 10273 2787 10287
rect 2793 10253 2807 10267
rect 2733 10232 2747 10246
rect 2773 10232 2787 10246
rect 2693 10213 2707 10227
rect 2753 10173 2767 10187
rect 2773 10133 2787 10147
rect 2753 10113 2767 10127
rect 2633 10093 2647 10107
rect 2593 10053 2607 10067
rect 2713 10054 2727 10068
rect 2913 10274 2927 10288
rect 2813 10233 2827 10247
rect 2933 10232 2947 10246
rect 3173 10774 3187 10788
rect 3073 10673 3087 10687
rect 3153 10673 3167 10687
rect 3113 10574 3127 10588
rect 3293 10613 3307 10627
rect 3213 10574 3227 10588
rect 3093 10532 3107 10546
rect 3052 10352 3066 10366
rect 3073 10353 3087 10367
rect 3133 10353 3147 10367
rect 2933 10173 2947 10187
rect 2973 10173 2987 10187
rect 2913 10093 2927 10107
rect 2853 10073 2867 10087
rect 2893 10053 2907 10067
rect 2973 10054 2987 10068
rect 3013 10054 3027 10068
rect 2873 9893 2887 9907
rect 2693 9873 2707 9887
rect 2633 9813 2647 9827
rect 2573 9774 2587 9788
rect 2433 9733 2447 9747
rect 2613 9732 2627 9746
rect 2733 9793 2747 9807
rect 2413 9693 2427 9707
rect 2473 9693 2487 9707
rect 2433 9633 2447 9647
rect 2393 9613 2407 9627
rect 2513 9633 2527 9647
rect 2453 9453 2467 9467
rect 2493 9273 2507 9287
rect 2413 9234 2427 9248
rect 2453 9234 2467 9248
rect 2473 9192 2487 9206
rect 2413 9133 2427 9147
rect 2353 9093 2367 9107
rect 2393 9093 2407 9107
rect 2333 9073 2347 9087
rect 2473 8972 2487 8986
rect 2953 9873 2967 9887
rect 2893 9793 2907 9807
rect 2933 9773 2947 9787
rect 2913 9693 2927 9707
rect 2913 9653 2927 9667
rect 2873 9553 2887 9567
rect 2673 9534 2687 9548
rect 2653 9492 2667 9506
rect 2773 9333 2787 9347
rect 2713 9234 2727 9248
rect 2733 9173 2747 9187
rect 2693 9133 2707 9147
rect 2613 9113 2627 9127
rect 2693 9112 2707 9126
rect 2573 9073 2587 9087
rect 2533 9033 2547 9047
rect 2513 8913 2527 8927
rect 2433 8873 2447 8887
rect 2553 9013 2567 9027
rect 2553 8972 2567 8986
rect 2553 8933 2567 8947
rect 2533 8853 2547 8867
rect 2493 8833 2507 8847
rect 2473 8773 2487 8787
rect 2353 8733 2367 8747
rect 2433 8733 2447 8747
rect 2393 8714 2407 8728
rect 2313 8633 2327 8647
rect 2313 8593 2327 8607
rect 2413 8653 2427 8667
rect 2373 8553 2387 8567
rect 2393 8494 2407 8508
rect 2453 8494 2467 8508
rect 2373 8473 2387 8487
rect 2313 8452 2327 8466
rect 2433 8452 2447 8466
rect 2393 8413 2407 8427
rect 2373 8373 2387 8387
rect 2293 8353 2307 8367
rect 2233 8293 2247 8307
rect 2193 8213 2207 8227
rect 2073 8194 2087 8208
rect 2153 8194 2167 8208
rect 2313 8213 2327 8227
rect 2093 8033 2107 8047
rect 2133 8033 2147 8047
rect 2073 7993 2087 8007
rect 2053 7974 2067 7988
rect 2173 7974 2187 7988
rect 2073 7932 2087 7946
rect 2133 7932 2147 7946
rect 2193 7893 2207 7907
rect 2073 7873 2087 7887
rect 2033 7773 2047 7787
rect 1993 7713 2007 7727
rect 2033 7693 2047 7707
rect 1993 7674 2007 7688
rect 2093 7773 2107 7787
rect 2193 7733 2207 7747
rect 2093 7693 2107 7707
rect 2073 7674 2087 7688
rect 2453 8333 2467 8347
rect 2393 8273 2407 8287
rect 2333 8194 2347 8208
rect 2373 8194 2387 8208
rect 2413 8194 2427 8208
rect 2313 8133 2327 8147
rect 2273 8113 2287 8127
rect 2233 7973 2247 7987
rect 2312 8073 2326 8087
rect 2333 8073 2347 8087
rect 2433 8153 2447 8167
rect 2413 8113 2427 8127
rect 2433 8093 2447 8107
rect 2413 8073 2427 8087
rect 2393 8013 2407 8027
rect 2313 7974 2327 7988
rect 2393 7973 2407 7987
rect 2393 7933 2407 7947
rect 2333 7913 2347 7927
rect 2373 7913 2387 7927
rect 2253 7893 2267 7907
rect 2373 7853 2387 7867
rect 2233 7833 2247 7847
rect 1933 7632 1947 7646
rect 1973 7632 1987 7646
rect 2013 7593 2027 7607
rect 1913 7573 1927 7587
rect 1973 7573 1987 7587
rect 1893 7553 1907 7567
rect 1853 7473 1867 7487
rect 1833 7313 1847 7327
rect 1833 7253 1847 7267
rect 1813 7153 1827 7167
rect 1913 7454 1927 7468
rect 1953 7454 1967 7468
rect 1893 7412 1907 7426
rect 1853 7233 1867 7247
rect 1893 7193 1907 7207
rect 1852 7153 1866 7167
rect 1873 7153 1887 7167
rect 1793 7112 1807 7126
rect 1833 7113 1847 7127
rect 1693 7073 1707 7087
rect 1753 7073 1767 7087
rect 1673 7053 1687 7067
rect 1773 6993 1787 7007
rect 1653 6934 1667 6948
rect 1733 6934 1747 6948
rect 1893 7112 1907 7126
rect 1873 7053 1887 7067
rect 1913 7033 1927 7047
rect 1793 6873 1807 6887
rect 1853 6873 1867 6887
rect 1753 6813 1767 6827
rect 1833 6693 1847 6707
rect 1653 6673 1667 6687
rect 1633 6273 1647 6287
rect 1613 6213 1627 6227
rect 1513 6193 1527 6207
rect 1533 6114 1547 6128
rect 1513 5993 1527 6007
rect 1513 5913 1527 5927
rect 1313 5833 1327 5847
rect 1233 5653 1247 5667
rect 1233 5393 1247 5407
rect 1073 5332 1087 5346
rect 1073 5074 1087 5088
rect 1133 5253 1147 5267
rect 1173 5173 1187 5187
rect 1213 5093 1227 5107
rect 1113 5033 1127 5047
rect 1193 5032 1207 5046
rect 1393 5852 1407 5866
rect 1493 5852 1507 5866
rect 1353 5713 1367 5727
rect 1273 5513 1287 5527
rect 1253 5013 1267 5027
rect 1173 4993 1187 5007
rect 1313 5413 1327 5427
rect 1313 5273 1327 5287
rect 1353 5473 1367 5487
rect 1353 5433 1367 5447
rect 1493 5793 1507 5807
rect 1613 6013 1627 6027
rect 1593 5993 1607 6007
rect 1793 6634 1807 6648
rect 2213 7673 2227 7687
rect 2313 7713 2327 7727
rect 2313 7633 2327 7647
rect 2533 8793 2547 8807
rect 2513 8733 2527 8747
rect 2493 8673 2507 8687
rect 2493 8553 2507 8567
rect 2493 8353 2507 8367
rect 2533 8714 2547 8728
rect 2533 8453 2547 8467
rect 2513 8113 2527 8127
rect 2653 9014 2667 9028
rect 2693 9014 2707 9028
rect 2753 9014 2767 9028
rect 2733 8973 2747 8987
rect 2713 8933 2727 8947
rect 2713 8853 2727 8867
rect 2613 8714 2627 8728
rect 2653 8714 2667 8728
rect 2673 8672 2687 8686
rect 2693 8653 2707 8667
rect 2673 8613 2687 8627
rect 2693 8593 2707 8607
rect 2673 8553 2687 8567
rect 2633 8513 2647 8527
rect 2573 8413 2587 8427
rect 2653 8452 2667 8466
rect 2693 8453 2707 8467
rect 2693 8413 2707 8427
rect 2613 8373 2627 8387
rect 2553 8293 2567 8307
rect 2613 8194 2627 8208
rect 2653 8172 2667 8186
rect 2973 9732 2987 9746
rect 3113 10313 3127 10327
rect 3153 10274 3167 10288
rect 3073 10233 3087 10247
rect 3133 10232 3147 10246
rect 3173 10213 3187 10227
rect 3233 10313 3247 10327
rect 3233 10233 3247 10247
rect 3393 11094 3407 11108
rect 3433 11094 3447 11108
rect 3533 11093 3547 11107
rect 3693 11094 3707 11108
rect 3393 11053 3407 11067
rect 3513 11052 3527 11066
rect 3493 11033 3507 11047
rect 3473 11013 3487 11027
rect 3453 10973 3467 10987
rect 3373 10813 3387 10827
rect 3433 10793 3447 10807
rect 3373 10753 3387 10767
rect 3353 10713 3367 10727
rect 3373 10613 3387 10627
rect 3313 10573 3327 10587
rect 3353 10574 3367 10588
rect 3373 10532 3387 10546
rect 3433 10573 3447 10587
rect 3353 10513 3367 10527
rect 3313 10493 3327 10507
rect 3293 10213 3307 10227
rect 3213 10193 3227 10207
rect 3133 10173 3147 10187
rect 3153 10133 3167 10147
rect 3053 9973 3067 9987
rect 3053 9873 3067 9887
rect 2953 9573 2967 9587
rect 2993 9573 3007 9587
rect 3113 9853 3127 9867
rect 3113 9813 3127 9827
rect 3113 9754 3127 9768
rect 3053 9553 3067 9567
rect 2973 9533 2987 9547
rect 2933 9333 2947 9347
rect 3213 10054 3227 10068
rect 3293 10053 3307 10067
rect 3233 9973 3247 9987
rect 3213 9953 3227 9967
rect 3253 9953 3267 9967
rect 3173 9933 3187 9947
rect 3173 9853 3187 9867
rect 3153 9833 3167 9847
rect 3173 9754 3187 9768
rect 3133 9653 3147 9667
rect 3133 9553 3147 9567
rect 3073 9492 3087 9506
rect 3113 9493 3127 9507
rect 2993 9473 3007 9487
rect 2973 9253 2987 9267
rect 2793 9053 2807 9067
rect 2813 9013 2827 9027
rect 2793 8973 2807 8987
rect 2773 8952 2787 8966
rect 2873 9233 2887 9247
rect 2953 9234 2967 9248
rect 3133 9353 3147 9367
rect 3093 9253 3107 9267
rect 3013 9234 3027 9248
rect 3013 9193 3027 9207
rect 2933 9153 2947 9167
rect 3213 9693 3227 9707
rect 3193 9293 3207 9307
rect 3393 10373 3407 10387
rect 3473 10533 3487 10547
rect 3453 10373 3467 10387
rect 3333 10232 3347 10246
rect 3313 9933 3327 9947
rect 3413 10232 3427 10246
rect 3433 10193 3447 10207
rect 3473 10054 3487 10068
rect 3753 11074 3767 11088
rect 3853 11133 3867 11147
rect 3673 11052 3687 11066
rect 3713 11052 3727 11066
rect 3533 11033 3547 11047
rect 3853 11072 3867 11086
rect 3993 11072 4007 11086
rect 3713 11013 3727 11027
rect 3713 10853 3727 10867
rect 3613 10794 3627 10808
rect 3633 10752 3647 10766
rect 3573 10574 3587 10588
rect 3713 10753 3727 10767
rect 4153 10973 4167 10987
rect 4093 10913 4107 10927
rect 4113 10873 4127 10887
rect 4073 10814 4087 10828
rect 3913 10774 3927 10788
rect 4013 10774 4027 10788
rect 3733 10733 3747 10747
rect 3773 10733 3787 10747
rect 3533 10532 3547 10546
rect 3673 10533 3687 10547
rect 3593 10493 3607 10507
rect 3673 10373 3687 10387
rect 3613 10293 3627 10307
rect 3573 10253 3587 10267
rect 3713 10252 3727 10266
rect 3533 10233 3547 10247
rect 3633 10232 3647 10246
rect 3713 10213 3727 10227
rect 3533 10153 3547 10167
rect 3713 10153 3727 10167
rect 3373 9953 3387 9967
rect 3413 9953 3427 9967
rect 3513 10013 3527 10027
rect 3633 10073 3647 10087
rect 3693 10054 3707 10068
rect 3793 10574 3807 10588
rect 3933 10573 3947 10587
rect 4033 10753 4047 10767
rect 4053 10574 4067 10588
rect 4093 10574 4107 10588
rect 3813 10532 3827 10546
rect 3773 10393 3787 10407
rect 3933 10532 3947 10546
rect 3993 10532 4007 10546
rect 4033 10532 4047 10546
rect 4093 10393 4107 10407
rect 4173 10913 4187 10927
rect 4153 10813 4167 10827
rect 4173 10753 4187 10767
rect 4193 10733 4207 10747
rect 4473 10913 4487 10927
rect 4553 10913 4567 10927
rect 4373 10774 4387 10788
rect 4773 11133 4787 11147
rect 4833 11133 4847 11147
rect 4533 10814 4547 10828
rect 4813 10814 4827 10828
rect 4673 10733 4687 10747
rect 4193 10693 4207 10707
rect 4233 10693 4247 10707
rect 4133 10613 4147 10627
rect 4233 10613 4247 10627
rect 4293 10613 4307 10627
rect 4613 10613 4627 10627
rect 4453 10574 4467 10588
rect 4573 10573 4587 10587
rect 4593 10553 4607 10567
rect 4193 10532 4207 10546
rect 3973 10333 3987 10347
rect 4113 10333 4127 10347
rect 4153 10333 4167 10347
rect 3812 10253 3826 10267
rect 3833 10254 3847 10268
rect 3873 10153 3887 10167
rect 3933 10054 3947 10068
rect 3653 10012 3667 10026
rect 3713 10013 3727 10027
rect 3733 10013 3747 10027
rect 3573 9973 3587 9987
rect 3633 9973 3647 9987
rect 3533 9933 3547 9947
rect 3453 9893 3467 9907
rect 3553 9873 3567 9887
rect 3433 9754 3447 9768
rect 3473 9754 3487 9768
rect 3333 9713 3347 9727
rect 3373 9712 3387 9726
rect 3413 9633 3427 9647
rect 3293 9573 3307 9587
rect 3353 9573 3367 9587
rect 3273 9492 3287 9506
rect 3313 9473 3327 9487
rect 3173 9253 3187 9267
rect 3213 9234 3227 9248
rect 3193 9192 3207 9206
rect 3273 9192 3287 9206
rect 3113 9173 3127 9187
rect 3153 9173 3167 9187
rect 3273 9153 3287 9167
rect 3093 9113 3107 9127
rect 3253 9093 3267 9107
rect 2893 9014 2907 9028
rect 2773 8893 2787 8907
rect 2853 8893 2867 8907
rect 2853 8872 2867 8886
rect 2773 8853 2787 8867
rect 2753 8833 2767 8847
rect 2953 8952 2967 8966
rect 2973 8893 2987 8907
rect 2913 8813 2927 8827
rect 2933 8753 2947 8767
rect 2893 8714 2907 8728
rect 2813 8693 2827 8707
rect 2913 8653 2927 8667
rect 2753 8613 2767 8627
rect 2753 8573 2767 8587
rect 2833 8593 2847 8607
rect 2793 8573 2807 8587
rect 2913 8533 2927 8547
rect 2793 8513 2807 8527
rect 2853 8494 2867 8508
rect 2873 8452 2887 8466
rect 2913 8452 2927 8466
rect 3113 8913 3127 8927
rect 3033 8853 3047 8867
rect 3133 8853 3147 8867
rect 2993 8773 3007 8787
rect 3133 8813 3147 8827
rect 3213 8813 3227 8827
rect 3173 8793 3187 8807
rect 3313 9234 3327 9248
rect 3293 9053 3307 9067
rect 3273 8993 3287 9007
rect 3293 8933 3307 8947
rect 3253 8793 3267 8807
rect 3273 8773 3287 8787
rect 3213 8753 3227 8767
rect 3253 8753 3267 8767
rect 3213 8714 3227 8728
rect 3033 8673 3047 8687
rect 3113 8672 3127 8686
rect 3153 8672 3167 8686
rect 3193 8593 3207 8607
rect 3073 8533 3087 8547
rect 3153 8493 3167 8507
rect 2833 8433 2847 8447
rect 2973 8433 2987 8447
rect 3093 8433 3107 8447
rect 3053 8393 3067 8407
rect 2773 8353 2787 8367
rect 3133 8393 3147 8407
rect 2753 8233 2767 8247
rect 2733 8213 2747 8227
rect 2733 8173 2747 8187
rect 2493 7973 2507 7987
rect 2533 7973 2547 7987
rect 2633 8113 2647 8127
rect 2693 8113 2707 8127
rect 2593 8053 2607 8067
rect 2513 7932 2527 7946
rect 2473 7833 2487 7847
rect 2453 7813 2467 7827
rect 2653 7833 2667 7847
rect 2593 7793 2607 7807
rect 2633 7793 2647 7807
rect 2433 7693 2447 7707
rect 2333 7593 2347 7607
rect 2113 7573 2127 7587
rect 2253 7573 2267 7587
rect 2012 7533 2026 7547
rect 2033 7533 2047 7547
rect 2073 7533 2087 7547
rect 2053 7473 2067 7487
rect 2233 7533 2247 7547
rect 2213 7513 2227 7527
rect 2153 7473 2167 7487
rect 2213 7473 2227 7487
rect 2213 7433 2227 7447
rect 2253 7432 2267 7446
rect 2353 7432 2367 7446
rect 2133 7412 2147 7426
rect 2053 7353 2067 7367
rect 1993 7154 2007 7168
rect 1973 7112 1987 7126
rect 1933 6993 1947 7007
rect 2013 6973 2027 6987
rect 1973 6934 1987 6948
rect 2013 6873 2027 6887
rect 1993 6853 2007 6867
rect 2093 7333 2107 7347
rect 2093 7133 2107 7147
rect 2113 7093 2127 7107
rect 2113 7072 2127 7086
rect 2093 7053 2107 7067
rect 2073 6813 2087 6827
rect 2073 6634 2087 6648
rect 1773 6592 1787 6606
rect 1913 6593 1927 6607
rect 1993 6573 2007 6587
rect 2073 6573 2087 6587
rect 1813 6533 1827 6547
rect 1673 6513 1687 6527
rect 1713 6414 1727 6428
rect 1673 6173 1687 6187
rect 1653 5953 1667 5967
rect 1633 5894 1647 5908
rect 1613 5852 1627 5866
rect 1553 5833 1567 5847
rect 1653 5753 1667 5767
rect 1533 5713 1547 5727
rect 1593 5693 1607 5707
rect 1533 5594 1547 5608
rect 1573 5594 1587 5608
rect 1473 5493 1487 5507
rect 1433 5393 1447 5407
rect 1533 5473 1547 5487
rect 1513 5374 1527 5388
rect 1413 5332 1427 5346
rect 1373 5293 1387 5307
rect 1353 5213 1367 5227
rect 1333 5093 1347 5107
rect 1273 4973 1287 4987
rect 1173 4953 1187 4967
rect 1153 4933 1167 4947
rect 1133 4893 1147 4907
rect 1413 5153 1427 5167
rect 1473 5074 1487 5088
rect 1393 5032 1407 5046
rect 1353 4873 1367 4887
rect 1293 4853 1307 4867
rect 1413 4854 1427 4868
rect 1133 4813 1147 4827
rect 1213 4753 1227 4767
rect 1093 4713 1107 4727
rect 1073 4673 1087 4687
rect 1453 4812 1467 4826
rect 1453 4613 1467 4627
rect 1293 4573 1307 4587
rect 1433 4573 1447 4587
rect 1113 4554 1127 4568
rect 1333 4554 1347 4568
rect 1373 4554 1387 4568
rect 1233 4513 1247 4527
rect 1113 4493 1127 4507
rect 1093 4473 1107 4487
rect 1213 4353 1227 4367
rect 1153 4334 1167 4348
rect 1193 4334 1207 4348
rect 1133 4292 1147 4306
rect 933 4212 947 4226
rect 1053 4213 1067 4227
rect 853 3953 867 3967
rect 853 3813 867 3827
rect 893 3814 907 3828
rect 1133 4153 1147 4167
rect 993 4034 1007 4048
rect 1033 4034 1047 4048
rect 1193 4133 1207 4147
rect 1213 4073 1227 4087
rect 1213 4033 1227 4047
rect 993 3814 1007 3828
rect 813 3753 827 3767
rect 913 3753 927 3767
rect 873 3713 887 3727
rect 853 3613 867 3627
rect 993 3673 1007 3687
rect 953 3653 967 3667
rect 993 3652 1007 3666
rect 973 3613 987 3627
rect 933 3593 947 3607
rect 873 3553 887 3567
rect 913 3553 927 3567
rect 833 3514 847 3528
rect 873 3514 887 3528
rect 933 3533 947 3547
rect 813 3173 827 3187
rect 953 3513 967 3527
rect 893 3472 907 3486
rect 973 3472 987 3486
rect 953 3413 967 3427
rect 913 3373 927 3387
rect 953 3333 967 3347
rect 833 3113 847 3127
rect 873 3113 887 3127
rect 813 3093 827 3107
rect 733 2993 747 3007
rect 653 2893 667 2907
rect 633 2793 647 2807
rect 673 2774 687 2788
rect 553 2713 567 2727
rect 533 2693 547 2707
rect 513 2613 527 2627
rect 453 2433 467 2447
rect 493 2433 507 2447
rect 373 2253 387 2267
rect 413 2212 427 2226
rect 293 1773 307 1787
rect 173 1673 187 1687
rect 253 1673 267 1687
rect 193 1493 207 1507
rect 93 1392 107 1406
rect 73 1273 87 1287
rect 213 1392 227 1406
rect 393 2053 407 2067
rect 413 1912 427 1926
rect 493 1912 507 1926
rect 373 1873 387 1887
rect 413 1734 427 1748
rect 393 1692 407 1706
rect 473 1673 487 1687
rect 413 1593 427 1607
rect 193 1353 207 1367
rect 333 1353 347 1367
rect 433 1392 447 1406
rect 413 1353 427 1367
rect 393 1313 407 1327
rect 213 1172 227 1186
rect 393 1172 407 1186
rect 133 933 147 947
rect 173 933 187 947
rect 233 914 247 928
rect 373 914 387 928
rect 413 914 427 928
rect 433 913 447 927
rect 453 914 467 928
rect 173 872 187 886
rect 233 873 247 887
rect 393 872 407 886
rect 253 753 267 767
rect 193 733 207 747
rect 133 694 147 708
rect 133 652 147 666
rect 213 652 227 666
rect 173 613 187 627
rect 393 694 407 708
rect 453 694 467 708
rect 413 652 427 666
rect 452 653 466 667
rect 673 2713 687 2727
rect 653 2613 667 2627
rect 533 2573 547 2587
rect 533 2533 547 2547
rect 593 2493 607 2507
rect 633 2474 647 2488
rect 573 2432 587 2446
rect 693 2673 707 2687
rect 673 2413 687 2427
rect 633 2353 647 2367
rect 693 2353 707 2367
rect 613 2313 627 2327
rect 573 2293 587 2307
rect 533 2273 547 2287
rect 533 1873 547 1887
rect 513 1734 527 1748
rect 493 1353 507 1367
rect 513 1313 527 1327
rect 513 873 527 887
rect 473 652 487 666
rect 253 613 267 627
rect 213 453 227 467
rect 373 433 387 447
rect 453 433 467 447
rect 113 394 127 408
rect 153 394 167 408
rect 333 407 347 408
rect 93 353 107 367
rect 333 394 347 407
rect 413 394 427 408
rect 173 352 187 366
rect 113 213 127 227
rect 173 213 187 227
rect 213 174 227 188
rect 393 352 407 366
rect 413 273 427 287
rect 413 213 427 227
rect 333 173 347 187
rect 393 132 407 146
rect 453 133 467 147
rect 713 2293 727 2307
rect 573 2212 587 2226
rect 613 2212 627 2226
rect 613 2033 627 2047
rect 693 2113 707 2127
rect 653 1953 667 1967
rect 713 1954 727 1968
rect 593 1912 607 1926
rect 633 1912 647 1926
rect 693 1912 707 1926
rect 613 1793 627 1807
rect 653 1734 667 1748
rect 633 1692 647 1706
rect 593 1653 607 1667
rect 633 1633 647 1647
rect 613 1392 627 1406
rect 553 1213 567 1227
rect 613 1214 627 1228
rect 653 1213 667 1227
rect 673 1214 687 1228
rect 633 1172 647 1186
rect 593 914 607 928
rect 573 872 587 886
rect 613 853 627 867
rect 613 753 627 767
rect 573 694 587 708
rect 793 2873 807 2887
rect 833 2913 847 2927
rect 913 3213 927 3227
rect 913 3173 927 3187
rect 953 3233 967 3247
rect 993 3233 1007 3247
rect 933 2993 947 3007
rect 893 2933 907 2947
rect 893 2853 907 2867
rect 933 2853 947 2867
rect 833 2813 847 2827
rect 873 2813 887 2827
rect 1053 3992 1067 4006
rect 1093 3992 1107 4006
rect 1133 3992 1147 4006
rect 1293 4493 1307 4507
rect 1273 4333 1287 4347
rect 1373 4493 1387 4507
rect 1313 4473 1327 4487
rect 1353 4353 1367 4367
rect 1393 4334 1407 4348
rect 1373 4292 1387 4306
rect 1433 4292 1447 4306
rect 1333 4253 1347 4267
rect 1393 4253 1407 4267
rect 1313 4233 1327 4247
rect 1373 4093 1387 4107
rect 1353 4053 1367 4067
rect 1292 4033 1306 4047
rect 1313 4034 1327 4048
rect 1053 3913 1067 3927
rect 1213 3913 1227 3927
rect 1033 3673 1047 3687
rect 1073 3893 1087 3907
rect 1133 3893 1147 3907
rect 1073 3772 1087 3786
rect 1153 3772 1167 3786
rect 1213 3773 1227 3787
rect 1113 3514 1127 3528
rect 1093 3472 1107 3486
rect 1233 3453 1247 3467
rect 1053 3294 1067 3308
rect 1293 3993 1307 4007
rect 1273 3873 1287 3887
rect 1253 3333 1267 3347
rect 1013 3213 1027 3227
rect 1153 3294 1167 3308
rect 1153 3213 1167 3227
rect 1133 3133 1147 3147
rect 973 2793 987 2807
rect 833 2732 847 2746
rect 873 2732 887 2746
rect 813 2613 827 2627
rect 893 2573 907 2587
rect 893 2533 907 2547
rect 773 2493 787 2507
rect 753 2474 767 2488
rect 853 2474 867 2488
rect 873 2432 887 2446
rect 833 2413 847 2427
rect 933 2513 947 2527
rect 933 2432 947 2446
rect 793 2373 807 2387
rect 773 2333 787 2347
rect 753 2253 767 2267
rect 753 2213 767 2227
rect 873 2313 887 2327
rect 833 2293 847 2307
rect 873 2273 887 2287
rect 913 2193 927 2207
rect 953 2273 967 2287
rect 953 2213 967 2227
rect 933 1973 947 1987
rect 793 1954 807 1968
rect 833 1954 847 1968
rect 873 1954 887 1968
rect 753 1913 767 1927
rect 813 1912 827 1926
rect 733 1873 747 1887
rect 813 1833 827 1847
rect 733 1793 747 1807
rect 713 1593 727 1607
rect 813 1773 827 1787
rect 833 1753 847 1767
rect 773 1733 787 1747
rect 873 1693 887 1707
rect 933 1613 947 1627
rect 813 1593 827 1607
rect 773 1513 787 1527
rect 733 1453 747 1467
rect 853 1453 867 1467
rect 693 853 707 867
rect 673 733 687 747
rect 593 593 607 607
rect 773 1434 787 1448
rect 813 1434 827 1448
rect 1052 2933 1066 2947
rect 1013 2893 1027 2907
rect 1033 2873 1047 2887
rect 1073 2932 1087 2946
rect 1113 2933 1127 2947
rect 1113 2893 1127 2907
rect 1073 2793 1087 2807
rect 1073 2772 1087 2786
rect 1253 3252 1267 3266
rect 1333 3992 1347 4006
rect 1373 3893 1387 3907
rect 1313 3853 1327 3867
rect 1333 3814 1347 3828
rect 1673 5552 1687 5566
rect 1633 5374 1647 5388
rect 1733 6353 1747 6367
rect 1733 6313 1747 6327
rect 1713 6253 1727 6267
rect 1833 6473 1847 6487
rect 1953 6473 1967 6487
rect 1813 6133 1827 6147
rect 1793 6114 1807 6128
rect 1873 6414 1887 6428
rect 1913 6414 1927 6428
rect 1873 6353 1887 6367
rect 1953 6353 1967 6367
rect 1953 6313 1967 6327
rect 1913 6213 1927 6227
rect 1893 6133 1907 6147
rect 1733 6072 1747 6086
rect 1733 6033 1747 6047
rect 1773 5953 1787 5967
rect 1733 5852 1747 5866
rect 1733 5733 1747 5747
rect 1853 6072 1867 6086
rect 1893 5973 1907 5987
rect 1773 5653 1787 5667
rect 1833 5894 1847 5908
rect 1953 6173 1967 6187
rect 1953 6113 1967 6127
rect 1933 6093 1947 6107
rect 1913 5833 1927 5847
rect 1813 5593 1827 5607
rect 1893 5573 1907 5587
rect 1773 5552 1787 5566
rect 1833 5552 1847 5566
rect 1873 5553 1887 5567
rect 2113 7033 2127 7047
rect 2153 7233 2167 7247
rect 2233 7313 2247 7327
rect 2193 7174 2207 7188
rect 2153 7153 2167 7167
rect 2193 7153 2207 7167
rect 2673 7812 2687 7826
rect 2593 7772 2607 7786
rect 2653 7773 2667 7787
rect 2553 7693 2567 7707
rect 2633 7674 2647 7688
rect 2533 7633 2547 7647
rect 2513 7533 2527 7547
rect 2613 7632 2627 7646
rect 2593 7593 2607 7607
rect 2593 7533 2607 7547
rect 2573 7513 2587 7527
rect 2533 7493 2547 7507
rect 2633 7473 2647 7487
rect 2613 7433 2627 7447
rect 2553 7373 2567 7387
rect 2593 7373 2607 7387
rect 2333 7293 2347 7307
rect 2493 7293 2507 7307
rect 2273 7174 2287 7188
rect 2573 7233 2587 7247
rect 2293 7133 2307 7147
rect 2213 7112 2227 7126
rect 2333 7133 2347 7147
rect 2433 7134 2447 7148
rect 2313 7093 2327 7107
rect 2173 7013 2187 7027
rect 2233 6973 2247 6987
rect 2153 6934 2167 6948
rect 2193 6934 2207 6948
rect 2293 6953 2307 6967
rect 2133 6853 2147 6867
rect 2113 6553 2127 6567
rect 2093 6513 2107 6527
rect 2253 6873 2267 6887
rect 2213 6853 2227 6867
rect 2153 6693 2167 6707
rect 2213 6693 2227 6707
rect 2233 6592 2247 6606
rect 2273 6592 2287 6606
rect 2273 6513 2287 6527
rect 2053 6493 2067 6507
rect 2133 6493 2147 6507
rect 2033 6273 2047 6287
rect 2033 6193 2047 6207
rect 2093 6413 2107 6427
rect 2133 6414 2147 6428
rect 2173 6414 2187 6428
rect 2153 6372 2167 6386
rect 2153 6353 2167 6367
rect 2553 7013 2567 7027
rect 2393 6973 2407 6987
rect 2313 6934 2327 6948
rect 2293 6414 2307 6428
rect 2273 6333 2287 6347
rect 2153 6293 2167 6307
rect 2193 6293 2207 6307
rect 2193 6233 2207 6247
rect 2153 6173 2167 6187
rect 2133 6153 2147 6167
rect 2153 6133 2167 6147
rect 2173 6092 2187 6106
rect 2033 6072 2047 6086
rect 2073 6013 2087 6027
rect 2073 5992 2087 6006
rect 2013 5913 2027 5927
rect 1953 5873 1967 5887
rect 1953 5693 1967 5707
rect 2173 5933 2187 5947
rect 2113 5894 2127 5908
rect 2153 5893 2167 5907
rect 2052 5833 2066 5847
rect 2073 5833 2087 5847
rect 2113 5713 2127 5727
rect 2013 5673 2027 5687
rect 2453 6934 2467 6948
rect 2393 6892 2407 6906
rect 2433 6892 2447 6906
rect 2473 6873 2487 6887
rect 2513 6873 2527 6887
rect 2453 6813 2467 6827
rect 2393 6753 2407 6767
rect 2353 6673 2367 6687
rect 2453 6693 2467 6707
rect 2413 6634 2427 6648
rect 2353 6592 2367 6606
rect 2393 6592 2407 6606
rect 2433 6553 2447 6567
rect 2473 6513 2487 6527
rect 2393 6493 2407 6507
rect 2453 6473 2467 6487
rect 2373 6353 2387 6367
rect 2412 6353 2426 6367
rect 2433 6353 2447 6367
rect 2313 6213 2327 6227
rect 2493 6453 2507 6467
rect 2473 6373 2487 6387
rect 2453 6133 2467 6147
rect 2293 6113 2307 6127
rect 2433 6113 2447 6127
rect 2273 6093 2287 6107
rect 2213 5993 2227 6007
rect 2353 5993 2367 6007
rect 2393 5993 2407 6007
rect 2193 5852 2207 5866
rect 2313 5973 2327 5987
rect 2393 5873 2407 5887
rect 2293 5852 2307 5866
rect 2333 5833 2347 5847
rect 2213 5733 2227 5747
rect 2093 5613 2107 5627
rect 2173 5613 2187 5627
rect 2033 5552 2047 5566
rect 2073 5552 2087 5566
rect 1893 5493 1907 5507
rect 1833 5453 1847 5467
rect 1713 5393 1727 5407
rect 1813 5393 1827 5407
rect 1573 5333 1587 5347
rect 1953 5433 1967 5447
rect 1873 5413 1887 5427
rect 1833 5373 1847 5387
rect 1913 5374 1927 5388
rect 1513 5293 1527 5307
rect 1533 5233 1547 5247
rect 1493 4753 1507 4767
rect 1553 5113 1567 5127
rect 1813 5332 1827 5346
rect 1633 5173 1647 5187
rect 1693 5173 1707 5187
rect 1593 5074 1607 5088
rect 1613 5013 1627 5027
rect 1893 5332 1907 5346
rect 1853 5153 1867 5167
rect 1873 5113 1887 5127
rect 1713 5074 1727 5088
rect 1693 4953 1707 4967
rect 1593 4913 1607 4927
rect 1653 4913 1667 4927
rect 1573 4854 1587 4868
rect 1553 4773 1567 4787
rect 1533 4613 1547 4627
rect 1653 4854 1667 4868
rect 1593 4813 1607 4827
rect 1573 4593 1587 4607
rect 1673 4812 1687 4826
rect 1713 4812 1727 4826
rect 1693 4713 1707 4727
rect 1673 4693 1687 4707
rect 1633 4673 1647 4687
rect 1693 4633 1707 4647
rect 1693 4593 1707 4607
rect 1533 4573 1547 4587
rect 1573 4554 1587 4568
rect 1473 4513 1487 4527
rect 1553 4512 1567 4526
rect 1593 4493 1607 4507
rect 1513 4334 1527 4348
rect 1493 4293 1507 4307
rect 1453 4233 1467 4247
rect 1433 4173 1447 4187
rect 1413 4093 1427 4107
rect 1393 3873 1407 3887
rect 1473 4053 1487 4067
rect 1432 3992 1446 4006
rect 1453 3992 1467 4006
rect 1413 3814 1427 3828
rect 1353 3772 1367 3786
rect 1633 4273 1647 4287
rect 1693 4453 1707 4467
rect 1693 4334 1707 4348
rect 1693 4273 1707 4287
rect 1673 4233 1687 4247
rect 1573 4193 1587 4207
rect 1613 4173 1627 4187
rect 1573 4153 1587 4167
rect 1513 4093 1527 4107
rect 1513 4034 1527 4048
rect 1573 4034 1587 4048
rect 1673 4053 1687 4067
rect 1493 3793 1507 3807
rect 1473 3753 1487 3767
rect 1453 3733 1467 3747
rect 1393 3693 1407 3707
rect 1333 3573 1347 3587
rect 1413 3533 1427 3547
rect 1393 3453 1407 3467
rect 1313 3433 1327 3447
rect 1353 3433 1367 3447
rect 1293 3253 1307 3267
rect 1193 3193 1207 3207
rect 1173 2913 1187 2927
rect 1153 2873 1167 2887
rect 1153 2774 1167 2788
rect 1053 2713 1067 2727
rect 1353 3373 1367 3387
rect 1333 3333 1347 3347
rect 1313 3213 1327 3227
rect 1313 3073 1327 3087
rect 1293 3053 1307 3067
rect 1313 3033 1327 3047
rect 1333 2993 1347 3007
rect 1213 2893 1227 2907
rect 1133 2732 1147 2746
rect 1193 2733 1207 2747
rect 1113 2713 1127 2727
rect 1173 2693 1187 2707
rect 1073 2633 1087 2647
rect 1113 2633 1127 2647
rect 1113 2533 1127 2547
rect 1053 2474 1067 2488
rect 1093 2432 1107 2446
rect 1032 2373 1046 2387
rect 1053 2373 1067 2387
rect 1093 2373 1107 2387
rect 1013 2333 1027 2347
rect 1033 2293 1047 2307
rect 1033 2253 1047 2267
rect 1093 2333 1107 2347
rect 1113 2273 1127 2287
rect 1073 2212 1087 2226
rect 973 2113 987 2127
rect 993 2093 1007 2107
rect 1073 2073 1087 2087
rect 1013 1954 1027 1968
rect 1113 1967 1127 1968
rect 1113 1954 1127 1967
rect 1053 1912 1067 1926
rect 1113 1873 1127 1887
rect 1093 1853 1107 1867
rect 993 1813 1007 1827
rect 973 1753 987 1767
rect 1033 1753 1047 1767
rect 1013 1692 1027 1706
rect 1093 1653 1107 1667
rect 1053 1633 1067 1647
rect 973 1533 987 1547
rect 1033 1453 1047 1467
rect 1073 1434 1087 1448
rect 1053 1392 1067 1406
rect 953 1353 967 1367
rect 1053 1353 1067 1367
rect 833 1313 847 1327
rect 833 1273 847 1287
rect 833 1214 847 1228
rect 773 1173 787 1187
rect 813 1172 827 1186
rect 1053 1153 1067 1167
rect 873 993 887 1007
rect 793 914 807 928
rect 813 793 827 807
rect 833 773 847 787
rect 793 652 807 666
rect 913 953 927 967
rect 933 914 947 928
rect 973 914 987 928
rect 1013 914 1027 928
rect 973 853 987 867
rect 933 653 947 667
rect 973 652 987 666
rect 813 633 827 647
rect 873 633 887 647
rect 593 533 607 547
rect 733 533 747 547
rect 753 453 767 467
rect 533 353 547 367
rect 873 612 887 626
rect 833 593 847 607
rect 753 313 767 327
rect 593 293 607 307
rect 873 352 887 366
rect 833 273 847 287
rect 753 253 767 267
rect 793 253 807 267
rect 593 174 607 188
rect 813 213 827 227
rect 913 273 927 287
rect 613 132 627 146
rect 753 133 767 147
rect 793 132 807 146
rect 193 113 207 127
rect 473 113 487 127
rect 1153 2213 1167 2227
rect 1153 2173 1167 2187
rect 1193 2653 1207 2667
rect 1173 2033 1187 2047
rect 1153 1954 1167 1968
rect 1153 1912 1167 1926
rect 1193 1913 1207 1927
rect 1133 1853 1147 1867
rect 1133 1793 1147 1807
rect 1133 1692 1147 1706
rect 1313 2953 1327 2967
rect 1273 2933 1287 2947
rect 1373 3293 1387 3307
rect 1373 3233 1387 3247
rect 1373 2994 1387 3008
rect 1373 2933 1387 2947
rect 1593 3992 1607 4006
rect 1633 3933 1647 3947
rect 1613 3814 1627 3828
rect 1513 3733 1527 3747
rect 1573 3673 1587 3687
rect 1573 3593 1587 3607
rect 1593 3533 1607 3547
rect 1553 3514 1567 3528
rect 1433 3393 1447 3407
rect 1413 3353 1427 3367
rect 1473 3294 1487 3308
rect 1453 3252 1467 3266
rect 1533 3473 1547 3487
rect 1413 3213 1427 3227
rect 1513 3213 1527 3227
rect 1393 2893 1407 2907
rect 1333 2732 1347 2746
rect 1393 2733 1407 2747
rect 1373 2633 1387 2647
rect 1233 2573 1247 2587
rect 1233 2513 1247 2527
rect 1253 2474 1267 2488
rect 1293 2474 1307 2488
rect 1333 2474 1347 2488
rect 1393 2474 1407 2488
rect 1233 2393 1247 2407
rect 1313 2432 1327 2446
rect 1353 2432 1367 2446
rect 1353 2353 1367 2367
rect 1253 2333 1267 2347
rect 1233 2212 1247 2226
rect 1293 2254 1307 2268
rect 1333 2153 1347 2167
rect 1313 2073 1327 2087
rect 1233 2053 1247 2067
rect 1313 2033 1327 2047
rect 1293 2013 1307 2027
rect 1293 1954 1307 1968
rect 1273 1912 1287 1926
rect 1153 1434 1167 1448
rect 1113 1153 1127 1167
rect 1073 953 1087 967
rect 1253 1734 1267 1748
rect 1233 1633 1247 1647
rect 1273 1633 1287 1647
rect 1273 1612 1287 1626
rect 1213 1433 1227 1447
rect 1313 1433 1327 1447
rect 1213 1393 1227 1407
rect 1373 2313 1387 2327
rect 1393 2073 1407 2087
rect 1373 1773 1387 1787
rect 1353 1493 1367 1507
rect 1253 1392 1267 1406
rect 1333 1392 1347 1406
rect 1273 1353 1287 1367
rect 1193 1133 1207 1147
rect 1233 993 1247 1007
rect 1193 953 1207 967
rect 1153 914 1167 928
rect 1273 1133 1287 1147
rect 1053 833 1067 847
rect 1093 813 1107 827
rect 1033 733 1047 747
rect 1073 652 1087 666
rect 1133 652 1147 666
rect 993 613 1007 627
rect 1253 913 1267 927
rect 1213 872 1227 886
rect 1233 833 1247 847
rect 1033 593 1047 607
rect 1153 593 1167 607
rect 1013 352 1027 366
rect 1293 993 1307 1007
rect 1353 993 1367 1007
rect 1333 914 1347 928
rect 1353 873 1367 887
rect 1573 3472 1587 3486
rect 1833 5074 1847 5088
rect 1933 5053 1947 5067
rect 1853 5032 1867 5046
rect 1893 5032 1907 5046
rect 1753 4993 1767 5007
rect 1733 4713 1747 4727
rect 1893 4933 1907 4947
rect 1773 4853 1787 4867
rect 1853 4854 1867 4868
rect 1933 4854 1947 4868
rect 1773 4773 1787 4787
rect 1773 4733 1787 4747
rect 1893 4793 1907 4807
rect 1893 4673 1907 4687
rect 1873 4592 1887 4606
rect 1753 4573 1767 4587
rect 1813 4573 1827 4587
rect 1793 4493 1807 4507
rect 1873 4513 1887 4527
rect 1753 4473 1767 4487
rect 1853 4473 1867 4487
rect 1833 4334 1847 4348
rect 1873 4292 1887 4306
rect 1773 4253 1787 4267
rect 1713 4193 1727 4207
rect 1693 3813 1707 3827
rect 1713 3793 1727 3807
rect 1693 3613 1707 3627
rect 1653 3533 1667 3547
rect 1573 3393 1587 3407
rect 1533 3193 1547 3207
rect 1573 3133 1587 3147
rect 1453 2994 1467 3008
rect 1493 2994 1507 3008
rect 1473 2952 1487 2966
rect 1513 2952 1527 2966
rect 1453 2933 1467 2947
rect 1433 2432 1447 2446
rect 1413 1773 1427 1787
rect 1413 1733 1427 1747
rect 1413 1553 1427 1567
rect 1393 1353 1407 1367
rect 1693 3473 1707 3487
rect 1833 4093 1847 4107
rect 1893 4093 1907 4107
rect 1893 4053 1907 4067
rect 1873 3992 1887 4006
rect 1853 3833 1867 3847
rect 1833 3814 1847 3828
rect 1793 3772 1807 3786
rect 1813 3733 1827 3747
rect 1773 3693 1787 3707
rect 1733 3593 1747 3607
rect 1713 3313 1727 3327
rect 1633 3293 1647 3307
rect 1753 3533 1767 3547
rect 1793 3472 1807 3486
rect 1833 3693 1847 3707
rect 1793 3353 1807 3367
rect 1853 3653 1867 3667
rect 2533 6852 2547 6866
rect 2633 7413 2647 7427
rect 2693 7673 2707 7687
rect 2693 7632 2707 7646
rect 2673 7373 2687 7387
rect 2613 7353 2627 7367
rect 2633 7333 2647 7347
rect 2593 7173 2607 7187
rect 2613 7132 2627 7146
rect 2693 7253 2707 7267
rect 2673 7073 2687 7087
rect 2673 6973 2687 6987
rect 3053 8214 3067 8228
rect 3093 8212 3107 8226
rect 2893 8174 2907 8188
rect 3033 8153 3047 8167
rect 3013 8113 3027 8127
rect 3013 8073 3027 8087
rect 2953 8053 2967 8067
rect 2833 8033 2847 8047
rect 2933 8033 2947 8047
rect 2753 8013 2767 8027
rect 2793 8013 2807 8027
rect 2733 7972 2747 7986
rect 2792 7913 2806 7927
rect 2813 7913 2827 7927
rect 2853 7913 2867 7927
rect 2753 7853 2767 7867
rect 2793 7853 2807 7867
rect 2733 7613 2747 7627
rect 2813 7793 2827 7807
rect 2773 7713 2787 7727
rect 2813 7713 2827 7727
rect 2933 7932 2947 7946
rect 2893 7893 2907 7907
rect 2893 7872 2907 7886
rect 2873 7773 2887 7787
rect 2933 7793 2947 7807
rect 2913 7773 2927 7787
rect 2913 7733 2927 7747
rect 2893 7674 2907 7688
rect 2773 7632 2787 7646
rect 2753 7593 2767 7607
rect 2833 7632 2847 7646
rect 2873 7613 2887 7627
rect 2793 7573 2807 7587
rect 2873 7573 2887 7587
rect 2853 7533 2867 7547
rect 2753 7493 2767 7507
rect 2813 7412 2827 7426
rect 2853 7413 2867 7427
rect 2833 7393 2847 7407
rect 2813 7373 2827 7387
rect 2793 7353 2807 7367
rect 2773 7154 2787 7168
rect 2753 7112 2767 7126
rect 2773 7013 2787 7027
rect 2713 6973 2727 6987
rect 2613 6933 2627 6947
rect 2633 6892 2647 6906
rect 2573 6873 2587 6887
rect 2553 6813 2567 6827
rect 2553 6753 2567 6767
rect 2553 6592 2567 6606
rect 2533 6553 2547 6567
rect 2553 6533 2567 6547
rect 2513 6253 2527 6267
rect 2693 6953 2707 6967
rect 2753 6934 2767 6948
rect 2693 6892 2707 6906
rect 2653 6812 2667 6826
rect 2633 6753 2647 6767
rect 2613 6653 2627 6667
rect 2733 6813 2747 6827
rect 2733 6792 2747 6806
rect 2633 6592 2647 6606
rect 2633 6553 2647 6567
rect 2673 6533 2687 6547
rect 2713 6473 2727 6487
rect 2633 6433 2647 6447
rect 2613 6414 2627 6428
rect 2753 6753 2767 6767
rect 2793 6653 2807 6667
rect 2793 6573 2807 6587
rect 2893 7353 2907 7367
rect 2873 7293 2887 7307
rect 2933 7253 2947 7267
rect 2973 8033 2987 8047
rect 3093 8113 3107 8127
rect 3112 8073 3126 8087
rect 3133 8073 3147 8087
rect 3073 7974 3087 7988
rect 3013 7932 3027 7946
rect 3013 7833 3027 7847
rect 2973 7713 2987 7727
rect 3133 7974 3147 7988
rect 3133 7933 3147 7947
rect 3253 8672 3267 8686
rect 3233 8613 3247 8627
rect 3193 8293 3207 8307
rect 3193 8153 3207 8167
rect 3193 8073 3207 8087
rect 3293 8653 3307 8667
rect 3333 9093 3347 9107
rect 3373 9553 3387 9567
rect 3393 9533 3407 9547
rect 3373 9492 3387 9506
rect 3413 9473 3427 9487
rect 3393 9453 3407 9467
rect 3493 9713 3507 9727
rect 3513 9534 3527 9548
rect 3653 9773 3667 9787
rect 3613 9754 3627 9768
rect 3453 9433 3467 9447
rect 3513 9473 3527 9487
rect 3493 9393 3507 9407
rect 3373 9234 3387 9248
rect 3473 9192 3487 9206
rect 3533 9453 3547 9467
rect 3533 9432 3547 9446
rect 3553 9393 3567 9407
rect 3533 9193 3547 9207
rect 3433 9153 3447 9167
rect 3633 9712 3647 9726
rect 3753 9893 3767 9907
rect 3733 9773 3747 9787
rect 3773 9793 3787 9807
rect 3893 9793 3907 9807
rect 3733 9713 3747 9727
rect 3713 9673 3727 9687
rect 3753 9573 3767 9587
rect 3733 9553 3747 9567
rect 3933 9773 3947 9787
rect 4033 10313 4047 10327
rect 3993 10254 4007 10268
rect 3993 10193 4007 10207
rect 3993 10113 4007 10127
rect 4013 10073 4027 10087
rect 4013 10013 4027 10027
rect 4093 10274 4107 10288
rect 4133 10054 4147 10068
rect 4053 10013 4067 10027
rect 4033 9893 4047 9907
rect 4033 9853 4047 9867
rect 3993 9793 4007 9807
rect 3813 9754 3827 9768
rect 3853 9754 3867 9768
rect 3893 9754 3907 9768
rect 3773 9534 3787 9548
rect 3833 9713 3847 9727
rect 3713 9492 3727 9506
rect 3813 9493 3827 9507
rect 3753 9453 3767 9467
rect 3713 9393 3727 9407
rect 3753 9393 3767 9407
rect 3733 9373 3747 9387
rect 3433 9132 3447 9146
rect 3473 9133 3487 9147
rect 3553 9133 3567 9147
rect 3413 9113 3427 9127
rect 3393 9093 3407 9107
rect 3353 9033 3367 9047
rect 3373 9013 3387 9027
rect 3373 8973 3387 8987
rect 3393 8933 3407 8947
rect 3393 8893 3407 8907
rect 3373 8733 3387 8747
rect 3353 8714 3367 8728
rect 3453 9033 3467 9047
rect 3433 8973 3447 8987
rect 3413 8773 3427 8787
rect 3433 8753 3447 8767
rect 3433 8713 3447 8727
rect 3353 8653 3367 8667
rect 3292 8533 3306 8547
rect 3313 8533 3327 8547
rect 3273 8513 3287 8527
rect 3233 8393 3247 8407
rect 3333 8353 3347 8367
rect 3253 8333 3267 8347
rect 3273 8313 3287 8327
rect 3333 8293 3347 8307
rect 3273 8273 3287 8287
rect 3253 8233 3267 8247
rect 3293 8213 3307 8227
rect 3273 8152 3287 8166
rect 3313 8152 3327 8166
rect 3293 8073 3307 8087
rect 3213 7974 3227 7988
rect 3253 7974 3267 7988
rect 3333 7993 3347 8007
rect 3193 7693 3207 7707
rect 3113 7674 3127 7688
rect 3153 7673 3167 7687
rect 3073 7613 3087 7627
rect 3013 7573 3027 7587
rect 3053 7493 3067 7507
rect 2973 7453 2987 7467
rect 3013 7412 3027 7426
rect 2993 7313 3007 7327
rect 2953 7233 2967 7247
rect 2873 7154 2887 7168
rect 2913 7154 2927 7168
rect 2973 7154 2987 7168
rect 2893 7112 2907 7126
rect 2933 7112 2947 7126
rect 2873 7073 2887 7087
rect 2953 7073 2967 7087
rect 2893 7053 2907 7067
rect 2933 7053 2947 7067
rect 2933 7032 2947 7046
rect 2913 6993 2927 7007
rect 2993 7113 3007 7127
rect 3053 7173 3067 7187
rect 3053 7152 3067 7166
rect 2973 6993 2987 7007
rect 3053 7073 3067 7087
rect 2933 6973 2947 6987
rect 3033 6973 3047 6987
rect 3013 6953 3027 6967
rect 2913 6933 2927 6947
rect 2953 6934 2967 6948
rect 2833 6793 2847 6807
rect 2833 6673 2847 6687
rect 2773 6533 2787 6547
rect 2813 6533 2827 6547
rect 2993 6914 3007 6928
rect 3173 7613 3187 7627
rect 3153 7592 3167 7606
rect 3173 7513 3187 7527
rect 3093 7213 3107 7227
rect 3113 7154 3127 7168
rect 3273 7932 3287 7946
rect 3413 8672 3427 8686
rect 3373 8613 3387 8627
rect 3413 8513 3427 8527
rect 3373 8433 3387 8447
rect 3413 8433 3427 8447
rect 3353 7853 3367 7867
rect 3393 8233 3407 8247
rect 3653 9313 3667 9327
rect 3593 9293 3607 9307
rect 3573 9113 3587 9127
rect 3513 9013 3527 9027
rect 3573 9014 3587 9028
rect 3613 9273 3627 9287
rect 3693 9234 3707 9248
rect 3753 9234 3767 9248
rect 3633 9193 3647 9207
rect 3613 9153 3627 9167
rect 3493 8853 3507 8867
rect 3493 8773 3507 8787
rect 3493 8733 3507 8747
rect 3553 8972 3567 8986
rect 3613 8972 3627 8986
rect 3553 8933 3567 8947
rect 3533 8733 3547 8747
rect 3533 8673 3547 8687
rect 3513 8653 3527 8667
rect 3453 8513 3467 8527
rect 3713 9192 3727 9206
rect 3753 9193 3767 9207
rect 3673 9153 3687 9167
rect 3713 9153 3727 9167
rect 3653 9113 3667 9127
rect 3633 8873 3647 8887
rect 3593 8833 3607 8847
rect 3573 8813 3587 8827
rect 3593 8753 3607 8767
rect 3673 9073 3687 9087
rect 3693 9033 3707 9047
rect 3673 8953 3687 8967
rect 3693 8933 3707 8947
rect 3673 8853 3687 8867
rect 3653 8733 3667 8747
rect 3633 8714 3647 8728
rect 3613 8672 3627 8686
rect 3653 8653 3667 8667
rect 3793 9313 3807 9327
rect 3913 9693 3927 9707
rect 3973 9753 3987 9767
rect 3973 9693 3987 9707
rect 3873 9633 3887 9647
rect 3953 9633 3967 9647
rect 3913 9573 3927 9587
rect 3973 9573 3987 9587
rect 3853 9533 3867 9547
rect 3833 9393 3847 9407
rect 3833 9333 3847 9347
rect 3813 9233 3827 9247
rect 3793 9173 3807 9187
rect 3773 9113 3787 9127
rect 3773 9033 3787 9047
rect 3833 9033 3847 9047
rect 3733 9014 3747 9028
rect 3813 9014 3827 9028
rect 3973 9534 3987 9548
rect 3973 9473 3987 9487
rect 3913 9373 3927 9387
rect 3913 9273 3927 9287
rect 4013 9313 4027 9327
rect 3913 9173 3927 9187
rect 3893 9113 3907 9127
rect 3753 8933 3767 8947
rect 3833 8972 3847 8986
rect 3793 8893 3807 8907
rect 3733 8873 3747 8887
rect 3773 8873 3787 8887
rect 3633 8633 3647 8647
rect 3713 8633 3727 8647
rect 3553 8513 3567 8527
rect 3593 8473 3607 8487
rect 3453 8452 3467 8466
rect 3493 8452 3507 8466
rect 3393 8152 3407 8166
rect 3433 8152 3447 8166
rect 3413 8113 3427 8127
rect 3333 7833 3347 7847
rect 3353 7693 3367 7707
rect 3393 7694 3407 7708
rect 3533 8433 3547 8447
rect 3513 8194 3527 8208
rect 3493 8152 3507 8166
rect 3533 8152 3547 8166
rect 3493 8113 3507 8127
rect 3493 8053 3507 8067
rect 3453 8013 3467 8027
rect 3533 8013 3547 8027
rect 3513 7932 3527 7946
rect 3613 8373 3627 8387
rect 3613 8153 3627 8167
rect 3733 8613 3747 8627
rect 3733 8513 3747 8527
rect 3893 9013 3907 9027
rect 3893 8933 3907 8947
rect 3933 9133 3947 9147
rect 4133 9973 4147 9987
rect 4173 10153 4187 10167
rect 4153 9953 4167 9967
rect 4113 9873 4127 9887
rect 4073 9753 4087 9767
rect 4093 9712 4107 9726
rect 4173 9713 4187 9727
rect 4293 10532 4307 10546
rect 4433 10532 4447 10546
rect 4573 10532 4587 10546
rect 4313 10373 4327 10387
rect 4253 10313 4267 10327
rect 4273 10274 4287 10288
rect 4353 10274 4367 10288
rect 4293 10232 4307 10246
rect 4353 10233 4367 10247
rect 4453 10373 4467 10387
rect 4513 10333 4527 10347
rect 4453 10293 4467 10307
rect 4473 10274 4487 10288
rect 4493 10213 4507 10227
rect 4413 10193 4427 10207
rect 4253 10133 4267 10147
rect 4373 10133 4387 10147
rect 4273 10054 4287 10068
rect 4253 10013 4267 10027
rect 4313 10012 4327 10026
rect 4353 9992 4367 10006
rect 4393 9953 4407 9967
rect 4233 9933 4247 9947
rect 4133 9633 4147 9647
rect 4193 9633 4207 9647
rect 4073 9533 4087 9547
rect 4053 9273 4067 9287
rect 3953 9093 3967 9107
rect 4012 9093 4026 9107
rect 4033 9093 4047 9107
rect 3913 8873 3927 8887
rect 3813 8813 3827 8827
rect 3873 8813 3887 8827
rect 3793 8733 3807 8747
rect 3793 8673 3807 8687
rect 3773 8494 3787 8508
rect 4013 9014 4027 9028
rect 4053 9013 4067 9027
rect 3993 8972 4007 8986
rect 4033 8953 4047 8967
rect 3853 8773 3867 8787
rect 3893 8714 3907 8728
rect 4093 9473 4107 9487
rect 4173 9573 4187 9587
rect 4213 9573 4227 9587
rect 4333 9853 4347 9867
rect 4253 9793 4267 9807
rect 4293 9754 4307 9768
rect 4273 9713 4287 9727
rect 4253 9693 4267 9707
rect 4313 9712 4327 9726
rect 4353 9693 4367 9707
rect 4393 9673 4407 9687
rect 4713 10574 4727 10588
rect 4653 10532 4667 10546
rect 4793 10574 4807 10588
rect 4653 10453 4667 10467
rect 4613 10193 4627 10207
rect 4533 10133 4547 10147
rect 4513 9933 4527 9947
rect 4493 9913 4507 9927
rect 4433 9773 4447 9787
rect 4313 9633 4327 9647
rect 4413 9633 4427 9647
rect 4273 9553 4287 9567
rect 4253 9534 4267 9548
rect 4293 9513 4307 9527
rect 4233 9492 4247 9506
rect 4273 9492 4287 9506
rect 4193 9473 4207 9487
rect 4193 9433 4207 9447
rect 4273 9393 4287 9407
rect 4253 9373 4267 9387
rect 4173 9333 4187 9347
rect 4133 9233 4147 9247
rect 4153 9192 4167 9206
rect 4193 9192 4207 9206
rect 4233 9192 4247 9206
rect 4173 9093 4187 9107
rect 4113 8973 4127 8987
rect 4153 8972 4167 8986
rect 4093 8953 4107 8967
rect 3953 8714 3967 8728
rect 3873 8672 3887 8686
rect 3893 8653 3907 8667
rect 3873 8613 3887 8627
rect 3833 8533 3847 8547
rect 3813 8493 3827 8507
rect 3853 8493 3867 8507
rect 3753 8353 3767 8367
rect 3833 8333 3847 8347
rect 3793 8313 3807 8327
rect 3813 8293 3827 8307
rect 3693 8253 3707 8267
rect 3833 8233 3847 8247
rect 3753 8194 3767 8208
rect 3693 8152 3707 8166
rect 3733 8152 3747 8166
rect 3633 8053 3647 8067
rect 3713 8073 3727 8087
rect 3713 8033 3727 8047
rect 3753 8033 3767 8047
rect 3713 7993 3727 8007
rect 3873 8473 3887 8487
rect 3993 8713 4007 8727
rect 3953 8653 3967 8667
rect 3913 8613 3927 8627
rect 3973 8593 3987 8607
rect 4073 8713 4087 8727
rect 4113 8714 4127 8728
rect 4013 8613 4027 8627
rect 3993 8573 4007 8587
rect 3973 8533 3987 8547
rect 4133 8672 4147 8686
rect 4093 8653 4107 8667
rect 4133 8633 4147 8647
rect 4073 8613 4087 8627
rect 3913 8494 3927 8508
rect 3973 8494 3987 8508
rect 4013 8493 4027 8507
rect 3913 8413 3927 8427
rect 3933 8293 3947 8307
rect 3893 8273 3907 8287
rect 4033 8452 4047 8466
rect 4033 8373 4047 8387
rect 3892 8213 3906 8227
rect 3913 8213 3927 8227
rect 3873 8113 3887 8127
rect 3853 8053 3867 8067
rect 3813 8033 3827 8047
rect 3773 7993 3787 8007
rect 3693 7932 3707 7946
rect 3733 7932 3747 7946
rect 3593 7893 3607 7907
rect 3473 7833 3487 7847
rect 3473 7793 3487 7807
rect 3453 7694 3467 7708
rect 3253 7653 3267 7667
rect 3433 7652 3447 7666
rect 3233 7633 3247 7647
rect 3233 7453 3247 7467
rect 3213 7393 3227 7407
rect 3193 7273 3207 7287
rect 3213 7193 3227 7207
rect 3193 7112 3207 7126
rect 3133 7073 3147 7087
rect 3333 7632 3347 7646
rect 3433 7613 3447 7627
rect 3293 7573 3307 7587
rect 3433 7513 3447 7527
rect 3553 7654 3567 7668
rect 3753 7853 3767 7867
rect 3853 8013 3867 8027
rect 3833 7993 3847 8007
rect 3813 7892 3827 7906
rect 3793 7813 3807 7827
rect 3753 7773 3767 7787
rect 3693 7633 3707 7647
rect 3493 7553 3507 7567
rect 3293 7454 3307 7468
rect 3333 7454 3347 7468
rect 3273 7412 3287 7426
rect 3293 7393 3307 7407
rect 3353 7373 3367 7387
rect 3393 7333 3407 7347
rect 3393 7253 3407 7267
rect 3353 7154 3367 7168
rect 3333 7112 3347 7126
rect 3373 7112 3387 7126
rect 3212 7053 3226 7067
rect 3233 7053 3247 7067
rect 3133 7033 3147 7047
rect 3313 7033 3327 7047
rect 3193 7013 3207 7027
rect 3333 6993 3347 7007
rect 3373 6973 3387 6987
rect 3333 6933 3347 6947
rect 3373 6933 3387 6947
rect 2973 6893 2987 6907
rect 2933 6873 2947 6887
rect 2913 6753 2927 6767
rect 2873 6634 2887 6648
rect 2953 6634 2967 6648
rect 2833 6493 2847 6507
rect 2873 6493 2887 6507
rect 2753 6414 2767 6428
rect 2733 6393 2747 6407
rect 2633 6372 2647 6386
rect 2673 6372 2687 6386
rect 2713 6373 2727 6387
rect 2913 6573 2927 6587
rect 2893 6473 2907 6487
rect 2973 6592 2987 6606
rect 2973 6493 2987 6507
rect 2793 6393 2807 6407
rect 2593 6333 2607 6347
rect 2593 6312 2607 6326
rect 2533 6193 2547 6207
rect 2533 6073 2547 6087
rect 2493 6013 2507 6027
rect 2533 6013 2547 6027
rect 2473 5893 2487 5907
rect 2453 5733 2467 5747
rect 2333 5693 2347 5707
rect 2433 5693 2447 5707
rect 2233 5594 2247 5608
rect 2293 5594 2307 5608
rect 2453 5673 2467 5687
rect 2213 5573 2227 5587
rect 2053 5473 2067 5487
rect 2173 5473 2187 5487
rect 2213 5453 2227 5467
rect 2093 5374 2107 5388
rect 2133 5374 2147 5388
rect 2193 5374 2207 5388
rect 2053 5332 2067 5346
rect 2113 5332 2127 5346
rect 2153 5332 2167 5346
rect 2133 5293 2147 5307
rect 2113 5273 2127 5287
rect 2193 5293 2207 5307
rect 2153 5173 2167 5187
rect 2093 5113 2107 5127
rect 2013 5093 2027 5107
rect 1993 5033 2007 5047
rect 1973 4993 1987 5007
rect 1953 4793 1967 4807
rect 1973 4773 1987 4787
rect 1933 4733 1947 4747
rect 1933 4653 1947 4667
rect 1973 4653 1987 4667
rect 2433 5593 2447 5607
rect 2273 5552 2287 5566
rect 2313 5533 2327 5547
rect 2273 5473 2287 5487
rect 2393 5473 2407 5487
rect 2233 5433 2247 5447
rect 2353 5413 2367 5427
rect 2293 5393 2307 5407
rect 2253 5293 2267 5307
rect 2313 5373 2327 5387
rect 2413 5373 2427 5387
rect 2413 5332 2427 5346
rect 2373 5273 2387 5287
rect 2233 5253 2247 5267
rect 2213 5233 2227 5247
rect 2253 5233 2267 5247
rect 2213 5193 2227 5207
rect 2213 5053 2227 5067
rect 2033 5033 2047 5047
rect 2013 4753 2027 4767
rect 2073 5032 2087 5046
rect 2073 4993 2087 5007
rect 2133 4913 2147 4927
rect 2093 4854 2107 4868
rect 2193 5033 2207 5047
rect 2213 4973 2227 4987
rect 2193 4853 2207 4867
rect 2113 4812 2127 4826
rect 2133 4793 2147 4807
rect 2033 4613 2047 4627
rect 1993 4593 2007 4607
rect 2113 4753 2127 4767
rect 2093 4593 2107 4607
rect 2053 4554 2067 4568
rect 1993 4512 2007 4526
rect 2033 4473 2047 4487
rect 2073 4393 2087 4407
rect 2093 4353 2107 4367
rect 2013 4334 2027 4348
rect 2073 4334 2087 4348
rect 2133 4713 2147 4727
rect 2133 4692 2147 4706
rect 2133 4473 2147 4487
rect 2153 4453 2167 4467
rect 1993 4313 2007 4327
rect 2013 4253 2027 4267
rect 2093 4292 2107 4306
rect 2053 4193 2067 4207
rect 1973 4073 1987 4087
rect 1913 3933 1927 3947
rect 1953 3933 1967 3947
rect 1933 3633 1947 3647
rect 1893 3593 1907 3607
rect 1853 3573 1867 3587
rect 1873 3552 1887 3566
rect 1913 3553 1927 3567
rect 1853 3433 1867 3447
rect 1853 3373 1867 3387
rect 1813 3313 1827 3327
rect 1793 3273 1807 3287
rect 1633 3253 1647 3267
rect 1713 3233 1727 3247
rect 1773 3233 1787 3247
rect 1653 3193 1667 3207
rect 1633 3033 1647 3047
rect 1633 2952 1647 2966
rect 1493 2893 1507 2907
rect 1613 2893 1627 2907
rect 1473 2533 1487 2547
rect 1593 2774 1607 2788
rect 1633 2774 1647 2788
rect 1533 2513 1547 2527
rect 1493 2473 1507 2487
rect 1633 2733 1647 2747
rect 1633 2513 1647 2527
rect 1573 2473 1587 2487
rect 1613 2473 1627 2487
rect 1473 2433 1487 2447
rect 1453 2353 1467 2367
rect 1553 2432 1567 2446
rect 1593 2432 1607 2446
rect 1493 2313 1507 2327
rect 1553 2293 1567 2307
rect 1513 2254 1527 2268
rect 1473 2093 1487 2107
rect 1573 2212 1587 2226
rect 1633 2273 1647 2287
rect 1613 2153 1627 2167
rect 1493 2013 1507 2027
rect 1473 1973 1487 1987
rect 1593 1993 1607 2007
rect 1533 1954 1547 1968
rect 1473 1912 1487 1926
rect 1513 1873 1527 1887
rect 1453 1813 1467 1827
rect 1453 1734 1467 1748
rect 1533 1692 1547 1706
rect 1493 1673 1507 1687
rect 1493 1473 1507 1487
rect 1573 1573 1587 1587
rect 1553 1553 1567 1567
rect 1533 1413 1547 1427
rect 1473 1392 1487 1406
rect 1513 1273 1527 1287
rect 1453 1253 1467 1267
rect 1453 1013 1467 1027
rect 1413 933 1427 947
rect 1453 914 1467 928
rect 1373 793 1387 807
rect 1333 773 1347 787
rect 1333 713 1347 727
rect 1473 872 1487 886
rect 1473 833 1487 847
rect 1373 694 1387 708
rect 1433 693 1447 707
rect 1273 653 1287 667
rect 1353 652 1367 666
rect 1393 652 1407 666
rect 1473 713 1487 727
rect 1452 652 1466 666
rect 1473 653 1487 667
rect 1553 1392 1567 1406
rect 1593 1473 1607 1487
rect 1572 1313 1586 1327
rect 1593 1313 1607 1327
rect 1593 1153 1607 1167
rect 1673 3173 1687 3187
rect 1713 3133 1727 3147
rect 1753 3093 1767 3107
rect 1713 2994 1727 3008
rect 1833 3253 1847 3267
rect 1833 3173 1847 3187
rect 1813 3133 1827 3147
rect 1813 3093 1827 3107
rect 1793 3053 1807 3067
rect 1693 2952 1707 2966
rect 1733 2833 1747 2847
rect 1833 3053 1847 3067
rect 1833 2933 1847 2947
rect 1733 2753 1747 2767
rect 1773 2732 1787 2746
rect 1793 2613 1807 2627
rect 1793 2553 1807 2567
rect 1773 2533 1787 2547
rect 1873 3293 1887 3307
rect 1913 3514 1927 3528
rect 1913 3473 1927 3487
rect 2113 4153 2127 4167
rect 1993 3992 2007 4006
rect 2093 3992 2107 4006
rect 2093 3953 2107 3967
rect 1993 3893 2007 3907
rect 2013 3814 2027 3828
rect 2053 3713 2067 3727
rect 2073 3693 2087 3707
rect 2053 3653 2067 3667
rect 1993 3514 2007 3528
rect 1933 3453 1947 3467
rect 1913 3373 1927 3387
rect 1913 3332 1927 3346
rect 1893 3213 1907 3227
rect 1873 3193 1887 3207
rect 1873 2993 1887 3007
rect 1873 2732 1887 2746
rect 1853 2493 1867 2507
rect 1813 2474 1827 2488
rect 1753 2393 1767 2407
rect 1713 2254 1727 2268
rect 1753 2254 1767 2268
rect 1793 2254 1807 2268
rect 1833 2313 1847 2327
rect 1833 2254 1847 2268
rect 1653 2213 1667 2227
rect 1793 2153 1807 2167
rect 1813 2013 1827 2027
rect 1693 1893 1707 1907
rect 1792 1954 1806 1968
rect 1813 1954 1827 1968
rect 1813 1833 1827 1847
rect 1873 2293 1887 2307
rect 1873 2133 1887 2147
rect 1853 2033 1867 2047
rect 1853 2012 1867 2026
rect 1833 1793 1847 1807
rect 1773 1773 1787 1787
rect 1953 3353 1967 3367
rect 1993 3453 2007 3467
rect 1973 3333 1987 3347
rect 1953 3293 1967 3307
rect 2033 3333 2047 3347
rect 2013 3313 2027 3327
rect 2073 3613 2087 3627
rect 2073 3333 2087 3347
rect 2053 3313 2067 3327
rect 1953 3113 1967 3127
rect 2073 3253 2087 3267
rect 2013 3213 2027 3227
rect 2073 3193 2087 3207
rect 2013 3133 2027 3147
rect 1933 3093 1947 3107
rect 1973 3093 1987 3107
rect 2012 3053 2026 3067
rect 2033 3053 2047 3067
rect 1933 3013 1947 3027
rect 1933 2933 1947 2947
rect 1993 2952 2007 2966
rect 2053 2973 2067 2987
rect 1953 2893 1967 2907
rect 2033 2893 2047 2907
rect 1953 2853 1967 2867
rect 2073 2953 2087 2967
rect 2093 2913 2107 2927
rect 2093 2892 2107 2906
rect 2073 2853 2087 2867
rect 2053 2833 2067 2847
rect 1973 2813 1987 2827
rect 1953 2793 1967 2807
rect 1933 2633 1947 2647
rect 1913 2573 1927 2587
rect 1913 2293 1927 2307
rect 1913 2193 1927 2207
rect 1993 2774 2007 2788
rect 1993 2693 2007 2707
rect 2013 2533 2027 2547
rect 2073 2733 2087 2747
rect 2093 2693 2107 2707
rect 2093 2633 2107 2647
rect 2033 2513 2047 2527
rect 2073 2513 2087 2527
rect 1973 2474 1987 2488
rect 1953 2353 1967 2367
rect 1993 2293 2007 2307
rect 2013 2273 2027 2287
rect 2013 2212 2027 2226
rect 1973 2153 1987 2167
rect 1893 2093 1907 2107
rect 1993 2053 2007 2067
rect 1893 1993 1907 2007
rect 1993 1993 2007 2007
rect 1953 1954 1967 1968
rect 1873 1933 1887 1947
rect 1993 1893 2007 1907
rect 1933 1873 1947 1887
rect 2013 1873 2027 1887
rect 2013 1813 2027 1827
rect 1913 1793 1927 1807
rect 1793 1753 1807 1767
rect 1713 1734 1727 1748
rect 1773 1733 1787 1747
rect 1673 1692 1687 1706
rect 1753 1673 1767 1687
rect 1633 1613 1647 1627
rect 1693 1473 1707 1487
rect 1773 1633 1787 1647
rect 1753 1453 1767 1467
rect 1673 1392 1687 1406
rect 1733 1392 1747 1406
rect 1633 1333 1647 1347
rect 1733 1333 1747 1347
rect 1713 1293 1727 1307
rect 1633 1253 1647 1267
rect 1673 1253 1687 1267
rect 1653 1213 1667 1227
rect 1873 1734 1887 1748
rect 2013 1773 2027 1787
rect 1893 1673 1907 1687
rect 1833 1653 1847 1667
rect 1893 1652 1907 1666
rect 1833 1473 1847 1487
rect 1813 1433 1827 1447
rect 1793 1333 1807 1347
rect 1753 1214 1767 1228
rect 1793 1213 1807 1227
rect 1613 1113 1627 1127
rect 1733 1172 1747 1186
rect 1693 1153 1707 1167
rect 1673 1053 1687 1067
rect 1713 933 1727 947
rect 1933 1593 1947 1607
rect 2073 2353 2087 2367
rect 2073 2213 2087 2227
rect 2053 2053 2067 2067
rect 2053 1954 2067 1968
rect 2133 4133 2147 4147
rect 2153 4053 2167 4067
rect 2193 4812 2207 4826
rect 2293 5074 2307 5088
rect 2353 5073 2367 5087
rect 2313 5032 2327 5046
rect 2333 4973 2347 4987
rect 2273 4953 2287 4967
rect 2313 4953 2327 4967
rect 2353 4953 2367 4967
rect 2273 4913 2287 4927
rect 2293 4893 2307 4907
rect 2253 4853 2267 4867
rect 2233 4653 2247 4667
rect 2193 4573 2207 4587
rect 2133 4013 2147 4027
rect 2133 3833 2147 3847
rect 2133 3773 2147 3787
rect 2173 3793 2187 3807
rect 2393 5153 2407 5167
rect 2373 4893 2387 4907
rect 2313 4873 2327 4887
rect 2333 4854 2347 4868
rect 2313 4812 2327 4826
rect 2353 4812 2367 4826
rect 2373 4773 2387 4787
rect 2273 4673 2287 4687
rect 2253 4573 2267 4587
rect 2293 4573 2307 4587
rect 2333 4573 2347 4587
rect 2273 4554 2287 4568
rect 2213 4512 2227 4526
rect 2253 4512 2267 4526
rect 2313 4513 2327 4527
rect 2293 4473 2307 4487
rect 2253 4334 2267 4348
rect 2333 4473 2347 4487
rect 2353 4393 2367 4407
rect 2393 4713 2407 4727
rect 2393 4613 2407 4627
rect 2373 4333 2387 4347
rect 2453 5533 2467 5547
rect 2533 5953 2547 5967
rect 2573 5993 2587 6007
rect 2573 5953 2587 5967
rect 2553 5933 2567 5947
rect 2573 5913 2587 5927
rect 2553 5733 2567 5747
rect 2533 5713 2547 5727
rect 2493 5613 2507 5627
rect 2573 5613 2587 5627
rect 2593 5593 2607 5607
rect 2473 5473 2487 5487
rect 2453 5374 2467 5388
rect 2433 5193 2447 5207
rect 2433 5074 2447 5088
rect 2472 5333 2486 5347
rect 2553 5552 2567 5566
rect 2753 6353 2767 6367
rect 2633 6333 2647 6347
rect 2673 6213 2687 6227
rect 2653 6073 2667 6087
rect 2833 6273 2847 6287
rect 2893 6372 2907 6386
rect 2873 6353 2887 6367
rect 2853 6253 2867 6267
rect 2733 6193 2747 6207
rect 2833 6193 2847 6207
rect 2733 6153 2747 6167
rect 2853 6153 2867 6167
rect 2773 6114 2787 6128
rect 2813 6114 2827 6128
rect 2693 6072 2707 6086
rect 2673 6033 2687 6047
rect 2653 5993 2667 6007
rect 2633 5813 2647 5827
rect 2653 5693 2667 5707
rect 2633 5673 2647 5687
rect 2633 5633 2647 5647
rect 2653 5613 2667 5627
rect 2633 5552 2647 5566
rect 2533 5513 2547 5527
rect 2613 5513 2627 5527
rect 2493 5332 2507 5346
rect 2553 5493 2567 5507
rect 2613 5492 2627 5506
rect 2553 5413 2567 5427
rect 2653 5473 2667 5487
rect 2693 5852 2707 5866
rect 2693 5813 2707 5827
rect 2693 5753 2707 5767
rect 2753 6072 2767 6086
rect 2793 6033 2807 6047
rect 2813 5973 2827 5987
rect 2753 5913 2767 5927
rect 2773 5894 2787 5908
rect 2853 5933 2867 5947
rect 2753 5852 2767 5866
rect 2793 5733 2807 5747
rect 2793 5673 2807 5687
rect 2813 5653 2827 5667
rect 2813 5594 2827 5608
rect 2673 5453 2687 5467
rect 2633 5413 2647 5427
rect 2593 5374 2607 5388
rect 2793 5552 2807 5566
rect 2753 5473 2767 5487
rect 2853 5473 2867 5487
rect 2733 5374 2747 5388
rect 2793 5453 2807 5467
rect 2813 5374 2827 5388
rect 2573 5332 2587 5346
rect 2613 5332 2627 5346
rect 2653 5332 2667 5346
rect 2653 5293 2667 5307
rect 2533 5273 2547 5287
rect 2573 5233 2587 5247
rect 2653 5233 2667 5247
rect 2593 5213 2607 5227
rect 2573 5133 2587 5147
rect 2553 5113 2567 5127
rect 2533 5074 2547 5088
rect 2613 5133 2627 5147
rect 2593 5113 2607 5127
rect 2433 5013 2447 5027
rect 2433 4953 2447 4967
rect 2433 4812 2447 4826
rect 2513 5032 2527 5046
rect 2493 5013 2507 5027
rect 2473 4733 2487 4747
rect 2713 5213 2727 5227
rect 2653 5073 2667 5087
rect 2733 5074 2747 5088
rect 2773 5073 2787 5087
rect 2713 5032 2727 5046
rect 2753 5032 2767 5046
rect 2553 4973 2567 4987
rect 2613 4973 2627 4987
rect 2673 4973 2687 4987
rect 2653 4953 2667 4967
rect 2593 4913 2607 4927
rect 2553 4874 2567 4888
rect 2513 4853 2527 4867
rect 2553 4853 2567 4867
rect 2573 4812 2587 4826
rect 2533 4793 2547 4807
rect 2513 4773 2527 4787
rect 2513 4733 2527 4747
rect 2493 4713 2507 4727
rect 2453 4653 2467 4667
rect 2493 4633 2507 4647
rect 2493 4573 2507 4587
rect 2433 4554 2447 4568
rect 2253 4233 2267 4247
rect 2233 4213 2247 4227
rect 2253 4173 2267 4187
rect 2233 3953 2247 3967
rect 2313 4133 2327 4147
rect 2373 4293 2387 4307
rect 2413 4293 2427 4307
rect 2433 4273 2447 4287
rect 2373 4193 2387 4207
rect 2353 4093 2367 4107
rect 2333 4073 2347 4087
rect 2333 4052 2347 4066
rect 2273 3893 2287 3907
rect 2313 3873 2327 3887
rect 2213 3753 2227 3767
rect 2273 3753 2287 3767
rect 2213 3653 2227 3667
rect 2193 3613 2207 3627
rect 2173 3593 2187 3607
rect 2253 3573 2267 3587
rect 2233 3514 2247 3528
rect 2273 3513 2287 3527
rect 2193 3472 2207 3486
rect 2213 3453 2227 3467
rect 2173 3333 2187 3347
rect 2153 3233 2167 3247
rect 2213 3213 2227 3227
rect 2233 3193 2247 3207
rect 2213 3153 2227 3167
rect 2193 3133 2207 3147
rect 2273 3132 2287 3146
rect 2253 3093 2267 3107
rect 2153 3013 2167 3027
rect 2173 2952 2187 2966
rect 2213 2913 2227 2927
rect 2313 3753 2327 3767
rect 2313 3732 2327 3746
rect 2333 3633 2347 3647
rect 2313 3453 2327 3467
rect 2313 3313 2327 3327
rect 2313 3252 2327 3266
rect 2413 4073 2427 4087
rect 2393 3933 2407 3947
rect 2433 4013 2447 4027
rect 2473 4473 2487 4487
rect 2573 4773 2587 4787
rect 2593 4673 2607 4687
rect 2553 4653 2567 4667
rect 2553 4473 2567 4487
rect 2533 4413 2547 4427
rect 2633 4812 2647 4826
rect 2633 4713 2647 4727
rect 2613 4613 2627 4627
rect 2633 4554 2647 4568
rect 2633 4513 2647 4527
rect 2633 4473 2647 4487
rect 2593 4353 2607 4367
rect 2533 4334 2547 4348
rect 2573 4334 2587 4348
rect 2513 4293 2527 4307
rect 2493 4133 2507 4147
rect 2473 4033 2487 4047
rect 2533 4093 2547 4107
rect 2453 3993 2467 4007
rect 2513 3992 2527 4006
rect 2453 3953 2467 3967
rect 2553 3953 2567 3967
rect 2433 3933 2447 3947
rect 2493 3893 2507 3907
rect 2493 3853 2507 3867
rect 2533 3853 2547 3867
rect 2513 3833 2527 3847
rect 2473 3814 2487 3828
rect 2533 3813 2547 3827
rect 2413 3793 2427 3807
rect 2453 3733 2467 3747
rect 2413 3693 2427 3707
rect 2393 3553 2407 3567
rect 2493 3653 2507 3667
rect 2493 3632 2507 3646
rect 2513 3613 2527 3627
rect 2453 3514 2467 3528
rect 2493 3514 2507 3528
rect 2353 3353 2367 3367
rect 2373 3333 2387 3347
rect 2353 3294 2367 3308
rect 2313 3213 2327 3227
rect 2313 3173 2327 3187
rect 2313 2993 2327 3007
rect 2313 2952 2327 2966
rect 2293 2893 2307 2907
rect 2293 2853 2307 2867
rect 2233 2774 2247 2788
rect 2273 2774 2287 2788
rect 2193 2732 2207 2746
rect 2253 2733 2267 2747
rect 2173 2713 2187 2727
rect 2153 2613 2167 2627
rect 2133 2513 2147 2527
rect 2173 2573 2187 2587
rect 2193 2533 2207 2547
rect 2253 2493 2267 2507
rect 2433 3472 2447 3486
rect 2473 3413 2487 3427
rect 2433 3333 2447 3347
rect 2393 3313 2407 3327
rect 2433 3312 2447 3326
rect 2453 3252 2467 3266
rect 2413 3113 2427 3127
rect 2373 3073 2387 3087
rect 2453 3073 2467 3087
rect 2413 3053 2427 3067
rect 2353 2993 2367 3007
rect 2333 2893 2347 2907
rect 2353 2793 2367 2807
rect 2353 2732 2367 2746
rect 2353 2693 2367 2707
rect 2333 2653 2347 2667
rect 2333 2573 2347 2587
rect 2333 2474 2347 2488
rect 2273 2432 2287 2446
rect 2313 2433 2327 2447
rect 2213 2352 2227 2366
rect 2193 2313 2207 2327
rect 2173 2253 2187 2267
rect 2273 2253 2287 2267
rect 2153 2212 2167 2226
rect 2193 2212 2207 2226
rect 2133 2173 2147 2187
rect 2233 2173 2247 2187
rect 2153 2033 2167 2047
rect 2193 1954 2207 1968
rect 2293 2173 2307 2187
rect 2273 2033 2287 2047
rect 2253 1953 2267 1967
rect 2093 1893 2107 1907
rect 2133 1893 2147 1907
rect 2173 1873 2187 1887
rect 2293 2013 2307 2027
rect 2273 1853 2287 1867
rect 2173 1833 2187 1847
rect 2133 1793 2147 1807
rect 2053 1773 2067 1787
rect 2053 1733 2067 1747
rect 2133 1734 2147 1748
rect 2212 1793 2226 1807
rect 2233 1793 2247 1807
rect 2033 1553 2047 1567
rect 2113 1553 2127 1567
rect 1933 1513 1947 1527
rect 1913 1493 1927 1507
rect 1973 1493 1987 1507
rect 2153 1453 2167 1467
rect 1973 1413 1987 1427
rect 2233 1734 2247 1748
rect 1873 1392 1887 1406
rect 1913 1392 1927 1406
rect 2093 1392 2107 1406
rect 2053 1353 2067 1367
rect 1993 1293 2007 1307
rect 1893 1253 1907 1267
rect 1853 1214 1867 1228
rect 1933 1214 1947 1228
rect 1973 1214 1987 1228
rect 1833 1172 1847 1186
rect 1893 1172 1907 1186
rect 2213 1392 2227 1406
rect 2133 1313 2147 1327
rect 2133 1292 2147 1306
rect 2093 1214 2107 1228
rect 2053 1153 2067 1167
rect 1953 1133 1967 1147
rect 1813 1073 1827 1087
rect 1893 1033 1907 1047
rect 1813 1013 1827 1027
rect 1853 1013 1867 1027
rect 1713 914 1727 928
rect 1793 914 1807 928
rect 1833 914 1847 928
rect 1573 872 1587 886
rect 1653 872 1667 886
rect 1693 872 1707 886
rect 1733 833 1747 847
rect 1613 694 1627 708
rect 1633 652 1647 666
rect 1533 613 1547 627
rect 1593 613 1607 627
rect 1593 573 1607 587
rect 1433 553 1447 567
rect 1573 453 1587 467
rect 1133 333 1147 347
rect 1233 333 1247 347
rect 1053 313 1067 327
rect 1213 253 1227 267
rect 973 213 987 227
rect 933 173 947 187
rect 1113 152 1127 166
rect 1213 152 1227 166
rect 1333 313 1347 327
rect 1313 293 1327 307
rect 1253 273 1267 287
rect 1893 993 1907 1007
rect 1893 914 1907 928
rect 1933 914 1947 928
rect 1832 873 1846 887
rect 1853 873 1867 887
rect 1913 872 1927 886
rect 1793 813 1807 827
rect 1953 813 1967 827
rect 1833 733 1847 747
rect 1773 693 1787 707
rect 1873 713 1887 727
rect 2013 733 2027 747
rect 2193 1214 2207 1228
rect 2233 1214 2247 1228
rect 2113 1133 2127 1147
rect 2213 1133 2227 1147
rect 2173 1113 2187 1127
rect 2213 1073 2227 1087
rect 2113 993 2127 1007
rect 2233 953 2247 967
rect 2133 914 2147 928
rect 2393 3013 2407 3027
rect 2493 3013 2507 3027
rect 2433 2952 2447 2966
rect 2473 2952 2487 2966
rect 2473 2813 2487 2827
rect 2433 2793 2447 2807
rect 2413 2732 2427 2746
rect 2373 2653 2387 2667
rect 2373 2333 2387 2347
rect 2533 3553 2547 3567
rect 2613 4273 2627 4287
rect 2633 3793 2647 3807
rect 2613 3733 2627 3747
rect 2753 4973 2767 4987
rect 2733 4913 2747 4927
rect 2733 4554 2747 4568
rect 2693 4512 2707 4526
rect 2673 4353 2687 4367
rect 2713 4393 2727 4407
rect 2833 5332 2847 5346
rect 2813 5293 2827 5307
rect 2853 5193 2867 5207
rect 2853 5033 2867 5047
rect 2833 4953 2847 4967
rect 2793 4933 2807 4947
rect 2853 4913 2867 4927
rect 2773 4873 2787 4887
rect 2833 4854 2847 4868
rect 2833 4793 2847 4807
rect 2813 4773 2827 4787
rect 2813 4533 2827 4547
rect 2753 4373 2767 4387
rect 2753 4334 2767 4348
rect 2793 4334 2807 4348
rect 2713 4293 2727 4307
rect 2773 4113 2787 4127
rect 2753 4053 2767 4067
rect 2673 4032 2687 4046
rect 2693 4033 2707 4047
rect 2713 4034 2727 4048
rect 2673 3973 2687 3987
rect 2793 3972 2807 3986
rect 2693 3814 2707 3828
rect 2733 3832 2747 3846
rect 2653 3753 2667 3767
rect 2733 3753 2747 3767
rect 2633 3713 2647 3727
rect 2593 3693 2607 3707
rect 2572 3653 2586 3667
rect 2593 3653 2607 3667
rect 2573 3573 2587 3587
rect 2573 3533 2587 3547
rect 2573 3473 2587 3487
rect 2653 3693 2667 3707
rect 2633 3613 2647 3627
rect 2613 3513 2627 3527
rect 2652 3514 2666 3528
rect 2673 3513 2687 3527
rect 2633 3472 2647 3486
rect 2713 3453 2727 3467
rect 2713 3413 2727 3427
rect 2673 3373 2687 3387
rect 2633 3294 2647 3308
rect 2713 3293 2727 3307
rect 2753 3433 2767 3447
rect 2653 3252 2667 3266
rect 2573 3233 2587 3247
rect 2613 3193 2627 3207
rect 2573 3153 2587 3167
rect 2553 3133 2567 3147
rect 2533 3073 2547 3087
rect 2552 3053 2566 3067
rect 2573 3053 2587 3067
rect 2573 2993 2587 3007
rect 2633 3073 2647 3087
rect 2633 2994 2647 3008
rect 2733 3252 2747 3266
rect 2693 3013 2707 3027
rect 2713 2994 2727 3008
rect 2633 2953 2647 2967
rect 2613 2932 2627 2946
rect 2673 2933 2687 2947
rect 2553 2793 2567 2807
rect 2593 2793 2607 2807
rect 2533 2713 2547 2727
rect 2533 2653 2547 2667
rect 2513 2593 2527 2607
rect 2453 2533 2467 2547
rect 2653 2793 2667 2807
rect 2653 2774 2667 2788
rect 2693 2774 2707 2788
rect 2613 2753 2627 2767
rect 2593 2693 2607 2707
rect 2613 2613 2627 2627
rect 2473 2474 2487 2488
rect 2433 2313 2447 2327
rect 2352 2273 2366 2287
rect 2373 2273 2387 2287
rect 2413 2273 2427 2287
rect 2573 2474 2587 2488
rect 2553 2313 2567 2327
rect 2493 2273 2507 2287
rect 2473 2254 2487 2268
rect 2373 2212 2387 2226
rect 2413 2212 2427 2226
rect 2473 2133 2487 2147
rect 2413 2013 2427 2027
rect 2333 1973 2347 1987
rect 2373 1973 2387 1987
rect 2453 1993 2467 2007
rect 2413 1954 2427 1968
rect 2393 1893 2407 1907
rect 2453 1853 2467 1867
rect 2313 1793 2327 1807
rect 2453 1793 2467 1807
rect 2313 1734 2327 1748
rect 2353 1734 2367 1748
rect 2393 1734 2407 1748
rect 2293 1653 2307 1667
rect 2373 1692 2387 1706
rect 2313 1493 2327 1507
rect 2353 1434 2367 1448
rect 2453 1692 2467 1706
rect 2413 1433 2427 1447
rect 2433 1434 2447 1448
rect 2433 1253 2447 1267
rect 2393 1214 2407 1228
rect 2493 1833 2507 1847
rect 2413 1172 2427 1186
rect 2473 1173 2487 1187
rect 2273 1033 2287 1047
rect 2353 953 2367 967
rect 2393 914 2407 928
rect 2433 913 2447 927
rect 2153 872 2167 886
rect 2253 872 2267 886
rect 2353 853 2367 867
rect 2113 813 2127 827
rect 2093 713 2107 727
rect 2073 694 2087 708
rect 2333 793 2347 807
rect 2293 713 2307 727
rect 2213 693 2227 707
rect 1813 652 1827 666
rect 1773 613 1787 627
rect 1953 652 1967 666
rect 2013 652 2027 666
rect 2053 652 2067 666
rect 2093 652 2107 666
rect 1853 573 1867 587
rect 1733 414 1747 428
rect 1933 453 1947 467
rect 1833 413 1847 427
rect 1693 372 1707 386
rect 1813 373 1827 387
rect 1693 213 1707 227
rect 1253 154 1267 168
rect 1333 154 1347 168
rect 1393 154 1407 168
rect 833 93 847 107
rect 913 93 927 107
rect 1273 73 1287 87
rect 2133 394 2147 408
rect 2313 652 2327 666
rect 2433 853 2447 867
rect 2453 793 2467 807
rect 2393 693 2407 707
rect 2373 613 2387 627
rect 2153 352 2167 366
rect 2213 352 2227 366
rect 1953 313 1967 327
rect 2193 293 2207 307
rect 2093 213 2107 227
rect 1793 112 1807 126
rect 2133 154 2147 168
rect 2333 433 2347 447
rect 2393 573 2407 587
rect 2513 1633 2527 1647
rect 2513 1533 2527 1547
rect 2653 2533 2667 2547
rect 2633 2493 2647 2507
rect 2633 2433 2647 2447
rect 2613 2313 2627 2327
rect 2773 3293 2787 3307
rect 2753 3073 2767 3087
rect 2753 3013 2767 3027
rect 2773 2952 2787 2966
rect 2753 2733 2767 2747
rect 2813 3793 2827 3807
rect 2893 6333 2907 6347
rect 2933 6173 2947 6187
rect 2893 6133 2907 6147
rect 2933 6113 2947 6127
rect 2893 6093 2907 6107
rect 2933 6072 2947 6086
rect 2893 6053 2907 6067
rect 2893 5993 2907 6007
rect 2913 5933 2927 5947
rect 2893 5873 2907 5887
rect 2933 5833 2947 5847
rect 2913 5733 2927 5747
rect 2893 5553 2907 5567
rect 2893 5473 2907 5487
rect 2993 6473 3007 6487
rect 3053 6833 3067 6847
rect 3033 6453 3047 6467
rect 3033 6413 3047 6427
rect 2993 6393 3007 6407
rect 3013 6233 3027 6247
rect 3013 6153 3027 6167
rect 2973 6113 2987 6127
rect 3233 6912 3247 6926
rect 3473 7493 3487 7507
rect 3473 7393 3487 7407
rect 3453 7193 3467 7207
rect 3453 7154 3467 7168
rect 3453 6933 3467 6947
rect 3393 6813 3407 6827
rect 3433 6813 3447 6827
rect 3433 6792 3447 6806
rect 3093 6753 3107 6767
rect 3233 6753 3247 6767
rect 3313 6753 3327 6767
rect 3333 6753 3347 6767
rect 3073 6693 3087 6707
rect 3152 6693 3166 6707
rect 3173 6693 3187 6707
rect 3093 6634 3107 6648
rect 3153 6633 3167 6647
rect 3133 6553 3147 6567
rect 3153 6513 3167 6527
rect 3273 6733 3287 6747
rect 3233 6634 3247 6648
rect 3173 6493 3187 6507
rect 3413 6673 3427 6687
rect 3353 6634 3367 6648
rect 3273 6593 3287 6607
rect 3373 6592 3387 6606
rect 3413 6592 3427 6606
rect 3312 6553 3326 6567
rect 3333 6553 3347 6567
rect 3293 6533 3307 6547
rect 3193 6473 3207 6487
rect 3233 6473 3247 6487
rect 3073 6414 3087 6428
rect 3113 6414 3127 6428
rect 3153 6414 3167 6428
rect 3193 6414 3207 6428
rect 3053 6393 3067 6407
rect 3053 6293 3067 6307
rect 3053 6213 3067 6227
rect 3033 6113 3047 6127
rect 2993 6053 3007 6067
rect 3093 6373 3107 6387
rect 3173 6333 3187 6347
rect 3153 6253 3167 6267
rect 3093 6153 3107 6167
rect 3133 6153 3147 6167
rect 3133 6072 3147 6086
rect 3313 6333 3327 6347
rect 3293 6293 3307 6307
rect 3233 6173 3247 6187
rect 3253 6153 3267 6167
rect 3213 6114 3227 6128
rect 2973 5973 2987 5987
rect 3073 5973 3087 5987
rect 3113 5933 3127 5947
rect 2993 5893 3007 5907
rect 3053 5894 3067 5908
rect 3153 5894 3167 5908
rect 2993 5852 3007 5866
rect 3073 5852 3087 5866
rect 3133 5853 3147 5867
rect 3013 5813 3027 5827
rect 2973 5793 2987 5807
rect 3053 5673 3067 5687
rect 3013 5594 3027 5608
rect 3033 5552 3047 5566
rect 2953 5413 2967 5427
rect 3153 5613 3167 5627
rect 3133 5553 3147 5567
rect 3013 5393 3027 5407
rect 3113 5393 3127 5407
rect 3053 5374 3067 5388
rect 2973 5353 2987 5367
rect 2933 5333 2947 5347
rect 2973 5293 2987 5307
rect 3013 5273 3027 5287
rect 3033 5213 3047 5227
rect 3013 5153 3027 5167
rect 3093 5333 3107 5347
rect 3073 5233 3087 5247
rect 3193 6072 3207 6086
rect 3273 6072 3287 6086
rect 3233 5933 3247 5947
rect 3233 5894 3247 5908
rect 3233 5853 3247 5867
rect 3253 5753 3267 5767
rect 3193 5594 3207 5608
rect 3313 6053 3327 6067
rect 3393 6414 3407 6428
rect 3393 6353 3407 6367
rect 3373 6153 3387 6167
rect 3373 6132 3387 6146
rect 3333 6013 3347 6027
rect 3333 5992 3347 6006
rect 3293 5953 3307 5967
rect 3373 5973 3387 5987
rect 3453 6293 3467 6307
rect 3693 7533 3707 7547
rect 3553 7454 3567 7468
rect 3533 7412 3547 7426
rect 3493 7353 3507 7367
rect 3493 7213 3507 7227
rect 3473 6253 3487 6267
rect 3453 6153 3467 6167
rect 3433 6133 3447 6147
rect 3513 7193 3527 7207
rect 3513 7113 3527 7127
rect 3593 7413 3607 7427
rect 3733 7593 3747 7607
rect 3793 7652 3807 7666
rect 3753 7573 3767 7587
rect 3793 7553 3807 7567
rect 3773 7513 3787 7527
rect 3853 7953 3867 7967
rect 3833 7853 3847 7867
rect 3853 7793 3867 7807
rect 3813 7493 3827 7507
rect 3793 7473 3807 7487
rect 3573 7373 3587 7387
rect 3633 7154 3647 7168
rect 3713 7133 3727 7147
rect 3533 7093 3547 7107
rect 3553 7073 3567 7087
rect 3533 7013 3547 7027
rect 3573 7013 3587 7027
rect 3553 6993 3567 7007
rect 3653 7093 3667 7107
rect 3653 7013 3667 7027
rect 3613 6973 3627 6987
rect 3553 6933 3567 6947
rect 3613 6934 3627 6948
rect 3693 6953 3707 6967
rect 3533 6813 3547 6827
rect 3513 6773 3527 6787
rect 3533 6753 3547 6767
rect 3513 6733 3527 6747
rect 3593 6873 3607 6887
rect 3633 6833 3647 6847
rect 3613 6813 3627 6827
rect 3593 6793 3607 6807
rect 3573 6693 3587 6707
rect 3573 6592 3587 6606
rect 3533 6553 3547 6567
rect 3533 6433 3547 6447
rect 3573 6433 3587 6447
rect 3433 6072 3447 6086
rect 3433 6051 3447 6065
rect 3413 5973 3427 5987
rect 3393 5833 3407 5847
rect 3393 5812 3407 5826
rect 3373 5773 3387 5787
rect 3353 5753 3367 5767
rect 3313 5673 3327 5687
rect 3173 5333 3187 5347
rect 3213 5513 3227 5527
rect 3273 5533 3287 5547
rect 3233 5393 3247 5407
rect 3313 5533 3327 5547
rect 3293 5513 3307 5527
rect 3313 5374 3327 5388
rect 3353 5374 3367 5388
rect 3213 5313 3227 5327
rect 3153 5273 3167 5287
rect 3193 5273 3207 5287
rect 3113 5233 3127 5247
rect 3033 5073 3047 5087
rect 2893 4993 2907 5007
rect 2913 4893 2927 4907
rect 2913 4854 2927 4868
rect 2953 4854 2967 4868
rect 2933 4773 2947 4787
rect 3033 4973 3047 4987
rect 3033 4854 3047 4868
rect 3113 5074 3127 5088
rect 3153 5074 3167 5088
rect 3253 5313 3267 5327
rect 3093 5032 3107 5046
rect 2953 4733 2967 4747
rect 2973 4713 2987 4727
rect 2953 4653 2967 4667
rect 3073 4793 3087 4807
rect 3053 4733 3067 4747
rect 3073 4673 3087 4687
rect 2973 4573 2987 4587
rect 3013 4573 3027 4587
rect 2893 4413 2907 4427
rect 2873 4233 2887 4247
rect 2953 4512 2967 4526
rect 2933 4373 2947 4387
rect 2913 4333 2927 4347
rect 2913 4273 2927 4287
rect 2853 4213 2867 4227
rect 2893 4213 2907 4227
rect 2873 4013 2887 4027
rect 3233 5073 3247 5087
rect 3173 5032 3187 5046
rect 3233 5033 3247 5047
rect 3213 5013 3227 5027
rect 3173 4993 3187 5007
rect 3153 4833 3167 4847
rect 3153 4793 3167 4807
rect 3193 4953 3207 4967
rect 3173 4773 3187 4787
rect 3153 4554 3167 4568
rect 3113 4473 3127 4487
rect 3073 4393 3087 4407
rect 2993 4334 3007 4348
rect 3033 4334 3047 4348
rect 3073 4334 3087 4348
rect 3013 4292 3027 4306
rect 3053 4292 3067 4306
rect 2973 4273 2987 4287
rect 2933 4253 2947 4267
rect 3033 4253 3047 4267
rect 3053 4213 3067 4227
rect 3013 4053 3027 4067
rect 2973 4034 2987 4048
rect 3033 4033 3047 4047
rect 2933 3992 2947 4006
rect 2913 3973 2927 3987
rect 2993 3992 3007 4006
rect 3033 3993 3047 4007
rect 2973 3973 2987 3987
rect 2953 3893 2967 3907
rect 2913 3814 2927 3828
rect 2833 3733 2847 3747
rect 2813 3713 2827 3727
rect 2893 3733 2907 3747
rect 2873 3693 2887 3707
rect 2833 3514 2847 3528
rect 2933 3633 2947 3647
rect 2913 3612 2927 3626
rect 2993 3893 3007 3907
rect 3033 3813 3047 3827
rect 3013 3733 3027 3747
rect 3092 4113 3106 4127
rect 3113 4113 3127 4127
rect 3313 5313 3327 5327
rect 3273 5233 3287 5247
rect 3293 5173 3307 5187
rect 3273 5113 3287 5127
rect 3333 5273 3347 5287
rect 3313 5013 3327 5027
rect 3293 4993 3307 5007
rect 3253 4953 3267 4967
rect 3313 4873 3327 4887
rect 3273 4854 3287 4868
rect 3293 4813 3307 4827
rect 3253 4773 3267 4787
rect 3273 4673 3287 4687
rect 3233 4573 3247 4587
rect 3213 4553 3227 4567
rect 3253 4554 3267 4568
rect 3153 4493 3167 4507
rect 3193 4493 3207 4507
rect 3173 4393 3187 4407
rect 3153 4273 3167 4287
rect 3213 4334 3227 4348
rect 3273 4533 3287 4547
rect 3353 5133 3367 5147
rect 3353 4873 3367 4887
rect 3333 4813 3347 4827
rect 3393 5553 3407 5567
rect 3393 5473 3407 5487
rect 3413 5313 3427 5327
rect 3453 6013 3467 6027
rect 3473 5933 3487 5947
rect 3473 5873 3487 5887
rect 3453 5813 3467 5827
rect 3673 6634 3687 6648
rect 3713 6873 3727 6887
rect 3793 7393 3807 7407
rect 3853 7253 3867 7267
rect 3833 7193 3847 7207
rect 3993 8193 4007 8207
rect 3913 8173 3927 8187
rect 3953 8153 3967 8167
rect 3933 8133 3947 8147
rect 4013 8152 4027 8166
rect 4093 8593 4107 8607
rect 4233 9073 4247 9087
rect 4213 9033 4227 9047
rect 4253 9014 4267 9028
rect 4213 8873 4227 8887
rect 4193 8793 4207 8807
rect 4173 8593 4187 8607
rect 4293 9313 4307 9327
rect 4293 9273 4307 9287
rect 4293 9213 4307 9227
rect 4473 9754 4487 9768
rect 4473 9713 4487 9727
rect 4373 9573 4387 9587
rect 4433 9573 4447 9587
rect 4413 9553 4427 9567
rect 4633 9873 4647 9887
rect 4613 9853 4627 9867
rect 4593 9793 4607 9807
rect 4553 9754 4567 9768
rect 4533 9673 4547 9687
rect 4573 9653 4587 9667
rect 4533 9633 4547 9647
rect 4493 9534 4507 9548
rect 4373 9492 4387 9506
rect 4433 9492 4447 9506
rect 4473 9453 4487 9467
rect 4333 9253 4347 9267
rect 4453 9253 4467 9267
rect 4333 9193 4347 9207
rect 4373 9192 4387 9206
rect 4313 8993 4327 9007
rect 4273 8913 4287 8927
rect 4233 8853 4247 8867
rect 4273 8773 4287 8787
rect 4253 8713 4267 8727
rect 4233 8672 4247 8686
rect 4213 8593 4227 8607
rect 4193 8573 4207 8587
rect 4353 9153 4367 9167
rect 4433 9153 4447 9167
rect 4513 9453 4527 9467
rect 4493 9273 4507 9287
rect 4613 9553 4627 9567
rect 4673 10413 4687 10427
rect 4813 10473 4827 10487
rect 4793 10333 4807 10347
rect 4693 10233 4707 10247
rect 4673 10113 4687 10127
rect 4773 10153 4787 10167
rect 4753 10133 4767 10147
rect 4713 10113 4727 10127
rect 4693 10073 4707 10087
rect 4773 10093 4787 10107
rect 4713 10034 4727 10048
rect 4753 10034 4767 10048
rect 4693 9833 4707 9847
rect 4653 9693 4667 9707
rect 4693 9673 4707 9687
rect 4693 9593 4707 9607
rect 4793 10033 4807 10047
rect 5073 11133 5087 11147
rect 4873 11094 4887 11108
rect 5013 11094 5027 11108
rect 4853 10533 4867 10547
rect 4993 11052 5007 11066
rect 4973 11013 4987 11027
rect 4933 10613 4947 10627
rect 4893 10532 4907 10546
rect 5213 11094 5227 11108
rect 5393 11094 5407 11108
rect 5353 10853 5367 10867
rect 5133 10574 5147 10588
rect 4953 10513 4967 10527
rect 5113 10513 5127 10527
rect 4833 10453 4847 10467
rect 4853 10373 4867 10387
rect 4853 10333 4867 10347
rect 4833 10233 4847 10247
rect 5173 10473 5187 10487
rect 5113 10293 5127 10307
rect 5613 11133 5627 11147
rect 5493 10873 5507 10887
rect 5353 10613 5367 10627
rect 5273 10574 5287 10588
rect 5333 10574 5347 10588
rect 5213 10473 5227 10487
rect 5193 10393 5207 10407
rect 5013 10254 5027 10268
rect 4833 10193 4847 10207
rect 4873 10193 4887 10207
rect 4813 9993 4827 10007
rect 5093 10153 5107 10167
rect 4873 10113 4887 10127
rect 4853 10013 4867 10027
rect 4853 9992 4867 10006
rect 4833 9973 4847 9987
rect 4793 9953 4807 9967
rect 4733 9873 4747 9887
rect 4773 9833 4787 9847
rect 4733 9753 4747 9767
rect 4813 9754 4827 9768
rect 4793 9712 4807 9726
rect 4773 9693 4787 9707
rect 4753 9673 4767 9687
rect 4713 9553 4727 9567
rect 4733 9534 4747 9548
rect 4673 9433 4687 9447
rect 4693 9413 4707 9427
rect 4753 9413 4767 9427
rect 4713 9393 4727 9407
rect 4693 9353 4707 9367
rect 4693 9273 4707 9287
rect 4493 9193 4507 9207
rect 4473 9093 4487 9107
rect 4433 9053 4447 9067
rect 4393 9014 4407 9028
rect 4473 9014 4487 9028
rect 4353 8973 4367 8987
rect 4413 8953 4427 8967
rect 4333 8933 4347 8947
rect 4393 8753 4407 8767
rect 4313 8713 4327 8727
rect 4353 8714 4367 8728
rect 4393 8713 4407 8727
rect 4273 8653 4287 8667
rect 4352 8633 4366 8647
rect 4373 8633 4387 8647
rect 4433 8933 4447 8947
rect 4413 8613 4427 8627
rect 4293 8593 4307 8607
rect 4353 8593 4367 8607
rect 4393 8593 4407 8607
rect 4473 8913 4487 8927
rect 4253 8533 4267 8547
rect 4132 8493 4146 8507
rect 4153 8493 4167 8507
rect 4113 8452 4127 8466
rect 4093 8213 4107 8227
rect 3973 8133 3987 8147
rect 3953 8113 3967 8127
rect 4033 8053 4047 8067
rect 3993 8033 4007 8047
rect 3933 8013 3947 8027
rect 3913 7993 3927 8007
rect 3953 7974 3967 7988
rect 4053 7993 4067 8007
rect 4033 7974 4047 7988
rect 4093 7974 4107 7988
rect 4073 7953 4087 7967
rect 3913 7932 3927 7946
rect 3973 7932 3987 7946
rect 4013 7932 4027 7946
rect 3893 7393 3907 7407
rect 4053 7932 4067 7946
rect 4033 7893 4047 7907
rect 3973 7873 3987 7887
rect 4013 7873 4027 7887
rect 3933 7733 3947 7747
rect 4033 7853 4047 7867
rect 4093 7932 4107 7946
rect 4073 7793 4087 7807
rect 4013 7753 4027 7767
rect 4053 7753 4067 7767
rect 4073 7673 4087 7687
rect 3933 7652 3947 7666
rect 3993 7613 4007 7627
rect 3973 7573 3987 7587
rect 3953 7513 3967 7527
rect 4013 7593 4027 7607
rect 4013 7533 4027 7547
rect 3993 7513 4007 7527
rect 4073 7553 4087 7567
rect 3973 7493 3987 7507
rect 4033 7493 4047 7507
rect 4073 7493 4087 7507
rect 4033 7472 4047 7486
rect 4093 7473 4107 7487
rect 3993 7454 4007 7468
rect 3973 7413 3987 7427
rect 3913 7273 3927 7287
rect 3893 7233 3907 7247
rect 3873 7173 3887 7187
rect 3773 7112 3787 7126
rect 3873 7112 3887 7126
rect 3753 6893 3767 6907
rect 3793 7053 3807 7067
rect 3853 6953 3867 6967
rect 3953 7313 3967 7327
rect 4013 7412 4027 7426
rect 4093 7412 4107 7426
rect 4053 7393 4067 7407
rect 3993 7373 4007 7387
rect 3973 7293 3987 7307
rect 3953 7173 3967 7187
rect 3733 6813 3747 6827
rect 3753 6753 3767 6767
rect 3753 6693 3767 6707
rect 3753 6634 3767 6648
rect 3833 6793 3847 6807
rect 3733 6592 3747 6606
rect 3673 6353 3687 6367
rect 3593 6233 3607 6247
rect 3553 6114 3567 6128
rect 3533 6053 3547 6067
rect 3593 6073 3607 6087
rect 3553 6033 3567 6047
rect 3573 5973 3587 5987
rect 3513 5953 3527 5967
rect 3533 5894 3547 5908
rect 3553 5852 3567 5866
rect 3813 6592 3827 6606
rect 3893 6753 3907 6767
rect 3733 6233 3747 6247
rect 3713 6153 3727 6167
rect 3633 6073 3647 6087
rect 3613 5833 3627 5847
rect 3453 5552 3467 5566
rect 3533 5493 3547 5507
rect 3573 5493 3587 5507
rect 3493 5453 3507 5467
rect 3513 5332 3527 5346
rect 3433 5093 3447 5107
rect 3533 5093 3547 5107
rect 3553 5074 3567 5088
rect 3533 5032 3547 5046
rect 3453 4993 3467 5007
rect 3393 4973 3407 4987
rect 3393 4952 3407 4966
rect 3473 4933 3487 4947
rect 3413 4854 3427 4868
rect 3513 4854 3527 4868
rect 3393 4813 3407 4827
rect 3373 4793 3387 4807
rect 3353 4713 3367 4727
rect 3393 4713 3407 4727
rect 3333 4653 3347 4667
rect 3373 4573 3387 4587
rect 3253 4273 3267 4287
rect 3172 4193 3186 4207
rect 3193 4193 3207 4207
rect 3173 4133 3187 4147
rect 3073 4073 3087 4087
rect 3073 4052 3087 4066
rect 3073 3933 3087 3947
rect 3213 4034 3227 4048
rect 3153 3973 3167 3987
rect 3213 3973 3227 3987
rect 3193 3953 3207 3967
rect 3213 3933 3227 3947
rect 3213 3912 3227 3926
rect 3153 3893 3167 3907
rect 3113 3853 3127 3867
rect 3053 3753 3067 3767
rect 3033 3713 3047 3727
rect 3053 3693 3067 3707
rect 3013 3673 3027 3687
rect 2993 3513 3007 3527
rect 3053 3514 3067 3528
rect 2833 3393 2847 3407
rect 2893 3393 2907 3407
rect 2893 3353 2907 3367
rect 2833 3333 2847 3347
rect 2813 3273 2827 3287
rect 2813 3213 2827 3227
rect 2813 3093 2827 3107
rect 2813 2893 2827 2907
rect 2933 3294 2947 3308
rect 2973 3273 2987 3287
rect 2913 3252 2927 3266
rect 2953 3252 2967 3266
rect 2893 3153 2907 3167
rect 2853 3113 2867 3127
rect 2893 3113 2907 3127
rect 2793 2693 2807 2707
rect 2793 2672 2807 2686
rect 2733 2553 2747 2567
rect 2693 2493 2707 2507
rect 2733 2474 2747 2488
rect 2713 2432 2727 2446
rect 2753 2413 2767 2427
rect 2653 2273 2667 2287
rect 2693 2273 2707 2287
rect 2673 2212 2687 2226
rect 2613 2173 2627 2187
rect 2693 2173 2707 2187
rect 2573 2073 2587 2087
rect 2593 1954 2607 1968
rect 2633 1954 2647 1968
rect 2553 1873 2567 1887
rect 2653 1873 2667 1887
rect 2613 1813 2627 1827
rect 2593 1734 2607 1748
rect 2673 1734 2687 1748
rect 2653 1713 2667 1727
rect 2613 1692 2627 1706
rect 2653 1652 2667 1666
rect 2653 1613 2667 1627
rect 2533 1473 2547 1487
rect 2553 1434 2567 1448
rect 2533 1333 2547 1347
rect 2673 1333 2687 1347
rect 2553 1214 2567 1228
rect 2593 1214 2607 1228
rect 2633 1214 2647 1228
rect 2553 1153 2567 1167
rect 2593 1033 2607 1047
rect 2613 953 2627 967
rect 2573 914 2587 928
rect 2593 872 2607 886
rect 2633 872 2647 886
rect 2533 773 2547 787
rect 2633 753 2647 767
rect 2673 753 2687 767
rect 2453 493 2467 507
rect 2413 394 2427 408
rect 2573 694 2587 708
rect 2553 652 2567 666
rect 2513 633 2527 647
rect 2713 1773 2727 1787
rect 2733 1733 2747 1747
rect 2773 2353 2787 2367
rect 3153 3633 3167 3647
rect 3133 3514 3147 3528
rect 3073 3472 3087 3486
rect 3113 3472 3127 3486
rect 3033 3453 3047 3467
rect 3153 3453 3167 3467
rect 3133 3433 3147 3447
rect 3013 3294 3027 3308
rect 3133 3373 3147 3387
rect 3113 3353 3127 3367
rect 3053 3333 3067 3347
rect 3033 3273 3047 3287
rect 3133 3294 3147 3308
rect 3193 3753 3207 3767
rect 3193 3413 3207 3427
rect 3113 3252 3127 3266
rect 3033 3233 3047 3247
rect 3013 3093 3027 3107
rect 2893 3032 2907 3046
rect 2993 3033 3007 3047
rect 2933 2994 2947 3008
rect 2993 2994 3007 3008
rect 2913 2952 2927 2966
rect 2993 2953 3007 2967
rect 2993 2913 3007 2927
rect 2853 2774 2867 2788
rect 2853 2693 2867 2707
rect 2833 2553 2847 2567
rect 2813 2413 2827 2427
rect 2813 2254 2827 2268
rect 2793 2193 2807 2207
rect 2813 2173 2827 2187
rect 2873 2673 2887 2687
rect 3093 3193 3107 3207
rect 3113 3173 3127 3187
rect 3093 3153 3107 3167
rect 3073 3053 3087 3067
rect 3073 2994 3087 3008
rect 3033 2893 3047 2907
rect 3013 2853 3027 2867
rect 3053 2813 3067 2827
rect 3133 3113 3147 3127
rect 3113 3053 3127 3067
rect 3233 3893 3247 3907
rect 3233 3793 3247 3807
rect 3293 4233 3307 4247
rect 3273 4133 3287 4147
rect 3273 4093 3287 4107
rect 3273 3814 3287 3828
rect 3233 3753 3247 3767
rect 3253 3733 3267 3747
rect 3253 3673 3267 3687
rect 3353 4473 3367 4487
rect 3433 4813 3447 4827
rect 3333 4453 3347 4467
rect 3413 4453 3427 4467
rect 3313 3973 3327 3987
rect 3553 4813 3567 4827
rect 3493 4793 3507 4807
rect 3453 4773 3467 4787
rect 3473 4693 3487 4707
rect 3473 4533 3487 4547
rect 3353 4413 3367 4427
rect 3373 4334 3387 4348
rect 3513 4753 3527 4767
rect 3532 4653 3546 4667
rect 3553 4653 3567 4667
rect 3553 4613 3567 4627
rect 3773 6493 3787 6507
rect 3832 6493 3846 6507
rect 3853 6493 3867 6507
rect 3813 6414 3827 6428
rect 3873 6372 3887 6386
rect 3773 6293 3787 6307
rect 3773 6173 3787 6187
rect 3773 6093 3787 6107
rect 3693 6033 3707 6047
rect 3653 5973 3667 5987
rect 3713 5973 3727 5987
rect 3653 5952 3667 5966
rect 3633 5333 3647 5347
rect 3833 6273 3847 6287
rect 3813 6072 3827 6086
rect 3833 5993 3847 6007
rect 3813 5973 3827 5987
rect 3753 5852 3767 5866
rect 3933 6853 3947 6867
rect 3933 6813 3947 6827
rect 3913 6333 3927 6347
rect 3973 7093 3987 7107
rect 3973 7053 3987 7067
rect 4153 8413 4167 8427
rect 4133 8152 4147 8166
rect 4233 8494 4247 8508
rect 4193 8433 4207 8447
rect 4193 8412 4207 8426
rect 4193 8293 4207 8307
rect 4233 8393 4247 8407
rect 4213 8253 4227 8267
rect 4173 8233 4187 8247
rect 4313 8313 4327 8327
rect 4253 8273 4267 8287
rect 4293 8273 4307 8287
rect 4173 8193 4187 8207
rect 4213 8193 4227 8207
rect 4173 8073 4187 8087
rect 4273 8152 4287 8166
rect 4233 8113 4247 8127
rect 4213 8093 4227 8107
rect 4193 8053 4207 8067
rect 4253 8033 4267 8047
rect 4293 7993 4307 8007
rect 4253 7974 4267 7988
rect 4193 7932 4207 7946
rect 4233 7913 4247 7927
rect 4173 7873 4187 7887
rect 4133 7833 4147 7847
rect 4173 7833 4187 7847
rect 4133 7733 4147 7747
rect 4173 7793 4187 7807
rect 4153 7493 4167 7507
rect 4153 7412 4167 7426
rect 4133 7393 4147 7407
rect 4093 7154 4107 7168
rect 4033 7093 4047 7107
rect 4113 7073 4127 7087
rect 4113 6993 4127 7007
rect 4073 6953 4087 6967
rect 4033 6893 4047 6907
rect 4173 7373 4187 7387
rect 4173 7154 4187 7168
rect 4293 7853 4307 7867
rect 4493 8813 4507 8827
rect 4672 9214 4686 9228
rect 4693 9213 4707 9227
rect 4533 9193 4547 9207
rect 4533 9133 4547 9147
rect 4753 9113 4767 9127
rect 4573 9093 4587 9107
rect 4553 9053 4567 9067
rect 4553 8972 4567 8986
rect 4533 8893 4547 8907
rect 4673 9073 4687 9087
rect 4613 9013 4627 9027
rect 4653 9014 4667 9028
rect 4693 9014 4707 9028
rect 4673 8972 4687 8986
rect 4713 8953 4727 8967
rect 4613 8933 4627 8947
rect 4573 8753 4587 8767
rect 4593 8733 4607 8747
rect 4553 8714 4567 8728
rect 4693 8714 4707 8728
rect 4653 8693 4667 8707
rect 4573 8672 4587 8686
rect 4793 9593 4807 9607
rect 4793 9492 4807 9506
rect 4833 9453 4847 9467
rect 4813 9393 4827 9407
rect 4793 9353 4807 9367
rect 4793 9273 4807 9287
rect 4833 9313 4847 9327
rect 4833 9273 4847 9287
rect 4953 10054 4967 10068
rect 5033 10053 5047 10067
rect 5073 10054 5087 10068
rect 4973 10012 4987 10026
rect 5093 10033 5107 10047
rect 5073 10013 5087 10027
rect 5133 10252 5147 10266
rect 5153 10233 5167 10247
rect 5233 10233 5247 10247
rect 5233 10212 5247 10226
rect 5213 10153 5227 10167
rect 5153 10054 5167 10068
rect 5193 10054 5207 10068
rect 5253 10053 5267 10067
rect 4893 9973 4907 9987
rect 5033 9973 5047 9987
rect 5013 9873 5027 9887
rect 4913 9754 4927 9768
rect 5093 9853 5107 9867
rect 5053 9754 5067 9768
rect 4893 9633 4907 9647
rect 4993 9712 5007 9726
rect 5033 9653 5047 9667
rect 4953 9553 4967 9567
rect 5013 9553 5027 9567
rect 4933 9492 4947 9506
rect 4973 9473 4987 9487
rect 4873 9453 4887 9467
rect 4953 9453 4967 9467
rect 4893 9393 4907 9407
rect 4873 9333 4887 9347
rect 4813 9253 4827 9267
rect 4793 9193 4807 9207
rect 4853 9153 4867 9167
rect 4793 9093 4807 9107
rect 4833 9053 4847 9067
rect 4813 8993 4827 9007
rect 4733 8893 4747 8907
rect 4713 8693 4727 8707
rect 4733 8673 4747 8687
rect 4693 8613 4707 8627
rect 4673 8593 4687 8607
rect 4653 8573 4667 8587
rect 4513 8533 4527 8547
rect 4493 8513 4507 8527
rect 4553 8513 4567 8527
rect 4453 8494 4467 8508
rect 4353 8373 4367 8387
rect 4473 8452 4487 8466
rect 4453 8433 4467 8447
rect 4453 8373 4467 8387
rect 4433 8353 4447 8367
rect 4373 8333 4387 8347
rect 4353 7893 4367 7907
rect 4333 7813 4347 7827
rect 4353 7773 4367 7787
rect 4393 8273 4407 8287
rect 4453 8194 4467 8208
rect 4493 8193 4507 8207
rect 4393 7993 4407 8007
rect 4393 7972 4407 7986
rect 4373 7753 4387 7767
rect 4353 7713 4367 7727
rect 4273 7693 4287 7707
rect 4313 7693 4327 7707
rect 4293 7632 4307 7646
rect 4253 7613 4267 7627
rect 4353 7613 4367 7627
rect 4493 8152 4507 8166
rect 4493 8093 4507 8107
rect 4473 7974 4487 7988
rect 4433 7893 4447 7907
rect 4533 8493 4547 8507
rect 4533 8452 4547 8466
rect 4513 7913 4527 7927
rect 4513 7873 4527 7887
rect 4493 7793 4507 7807
rect 4433 7733 4447 7747
rect 4433 7673 4447 7687
rect 4493 7674 4507 7688
rect 4793 8953 4807 8967
rect 4773 8873 4787 8887
rect 4973 9413 4987 9427
rect 4953 9333 4967 9347
rect 4953 9293 4967 9307
rect 4913 9193 4927 9207
rect 4953 9113 4967 9127
rect 4933 9093 4947 9107
rect 4913 9014 4927 9028
rect 5053 9633 5067 9647
rect 5113 9754 5127 9768
rect 5053 9473 5067 9487
rect 5053 9353 5067 9367
rect 5053 9313 5067 9327
rect 5033 9293 5047 9307
rect 5233 10013 5247 10027
rect 5213 9973 5227 9987
rect 5253 9933 5267 9947
rect 5233 9913 5247 9927
rect 5393 10613 5407 10627
rect 5313 10532 5327 10546
rect 5373 10533 5387 10547
rect 5293 10353 5307 10367
rect 5173 9893 5187 9907
rect 5273 9893 5287 9907
rect 5253 9754 5267 9768
rect 5133 9713 5147 9727
rect 5173 9712 5187 9726
rect 5233 9712 5247 9726
rect 5092 9573 5106 9587
rect 5113 9573 5127 9587
rect 5113 9534 5127 9548
rect 5213 9613 5227 9627
rect 5553 10853 5567 10867
rect 5733 11133 5747 11147
rect 5593 10752 5607 10766
rect 5713 10752 5727 10766
rect 5693 10693 5707 10707
rect 5593 10613 5607 10627
rect 5673 10574 5687 10588
rect 5573 10532 5587 10546
rect 5533 10413 5547 10427
rect 5393 10353 5407 10367
rect 5513 10353 5527 10367
rect 5493 10313 5507 10327
rect 5393 10293 5407 10307
rect 5433 10274 5447 10288
rect 5473 10274 5487 10288
rect 5313 10253 5327 10267
rect 5373 10232 5387 10246
rect 5493 10233 5507 10247
rect 5333 10193 5347 10207
rect 5313 10113 5327 10127
rect 5313 9853 5327 9867
rect 5313 9793 5327 9807
rect 5313 9633 5327 9647
rect 5153 9433 5167 9447
rect 5193 9433 5207 9447
rect 5093 9353 5107 9367
rect 5073 9293 5087 9307
rect 5153 9293 5167 9307
rect 5093 9253 5107 9267
rect 5073 9192 5087 9206
rect 5033 9153 5047 9167
rect 5073 9153 5087 9167
rect 5053 9133 5067 9147
rect 4993 9073 5007 9087
rect 4933 8972 4947 8986
rect 4993 8972 5007 8986
rect 4913 8951 4927 8965
rect 4893 8933 4907 8947
rect 4953 8933 4967 8947
rect 4853 8913 4867 8927
rect 4873 8853 4887 8867
rect 4813 8793 4827 8807
rect 4993 8913 5007 8927
rect 4953 8813 4967 8827
rect 4893 8793 4907 8807
rect 4973 8793 4987 8807
rect 4933 8773 4947 8787
rect 4793 8714 4807 8728
rect 4833 8714 4847 8728
rect 4893 8714 4907 8728
rect 4773 8673 4787 8687
rect 4813 8672 4827 8686
rect 4853 8672 4867 8686
rect 4833 8653 4847 8667
rect 4933 8733 4947 8747
rect 4933 8693 4947 8707
rect 4913 8673 4927 8687
rect 4893 8633 4907 8647
rect 4813 8613 4827 8627
rect 4873 8613 4887 8627
rect 4793 8573 4807 8587
rect 4773 8473 4787 8487
rect 4633 8453 4647 8467
rect 4553 8413 4567 8427
rect 4573 8233 4587 8247
rect 4553 8033 4567 8047
rect 4553 7933 4567 7947
rect 4653 8393 4667 8407
rect 4753 8453 4767 8467
rect 4733 8333 4747 8347
rect 4693 8233 4707 8247
rect 4573 7853 4587 7867
rect 4553 7813 4567 7827
rect 4513 7632 4527 7646
rect 4473 7593 4487 7607
rect 4453 7573 4467 7587
rect 4513 7573 4527 7587
rect 4413 7553 4427 7567
rect 4393 7513 4407 7527
rect 4453 7533 4467 7547
rect 4473 7493 4487 7507
rect 4413 7453 4427 7467
rect 4213 7353 4227 7367
rect 4373 7413 4387 7427
rect 4453 7412 4467 7426
rect 4353 7353 4367 7367
rect 4293 7193 4307 7207
rect 4333 7173 4347 7187
rect 4573 7674 4587 7688
rect 4613 8053 4627 8067
rect 4793 8373 4807 8387
rect 4973 8653 4987 8667
rect 4933 8573 4947 8587
rect 4953 8553 4967 8567
rect 4913 8533 4927 8547
rect 4973 8493 4987 8507
rect 4853 8473 4867 8487
rect 4873 8353 4887 8367
rect 4913 8413 4927 8427
rect 4893 8333 4907 8347
rect 4813 8313 4827 8327
rect 4873 8313 4887 8327
rect 4833 8233 4847 8247
rect 4873 8194 4887 8208
rect 4773 8033 4787 8047
rect 4853 8152 4867 8166
rect 5013 8873 5027 8887
rect 5073 9013 5087 9027
rect 5073 8972 5087 8986
rect 5173 9173 5187 9187
rect 5133 9113 5147 9127
rect 5113 9053 5127 9067
rect 5113 9014 5127 9028
rect 5433 10153 5447 10167
rect 5353 10054 5367 10068
rect 5393 10054 5407 10068
rect 5473 10113 5487 10127
rect 5353 10013 5367 10027
rect 5413 9993 5427 10007
rect 5673 10473 5687 10487
rect 5653 10413 5667 10427
rect 5533 10032 5547 10046
rect 5513 9993 5527 10007
rect 5433 9953 5447 9967
rect 5393 9893 5407 9907
rect 5353 9853 5367 9867
rect 5353 9793 5367 9807
rect 5293 9473 5307 9487
rect 5333 9473 5347 9487
rect 5273 9413 5287 9427
rect 5213 9373 5227 9387
rect 5213 9333 5227 9347
rect 5273 9293 5287 9307
rect 5253 9273 5267 9287
rect 5233 9234 5247 9248
rect 5233 9193 5247 9207
rect 5433 9793 5447 9807
rect 5433 9754 5447 9768
rect 5473 9754 5487 9768
rect 5493 9712 5507 9726
rect 5453 9673 5467 9687
rect 5433 9534 5447 9548
rect 5393 9473 5407 9487
rect 5353 9433 5367 9447
rect 5333 9234 5347 9248
rect 5313 9192 5327 9206
rect 5353 9192 5367 9206
rect 5293 9153 5307 9167
rect 5193 9093 5207 9107
rect 5253 9073 5267 9087
rect 5173 9014 5187 9028
rect 5233 9014 5247 9028
rect 5153 8972 5167 8986
rect 5193 8972 5207 8986
rect 5093 8913 5107 8927
rect 5033 8853 5047 8867
rect 5133 8913 5147 8927
rect 5113 8813 5127 8827
rect 5013 8713 5027 8727
rect 5073 8733 5087 8747
rect 5053 8672 5067 8686
rect 5113 8652 5127 8666
rect 5053 8633 5067 8647
rect 5073 8613 5087 8627
rect 5013 8553 5027 8567
rect 5033 8533 5047 8547
rect 5013 8513 5027 8527
rect 5053 8493 5067 8507
rect 5033 8473 5047 8487
rect 4933 8393 4947 8407
rect 4933 8194 4947 8208
rect 4913 8113 4927 8127
rect 4833 8073 4847 8087
rect 4933 8073 4947 8087
rect 4813 7993 4827 8007
rect 4713 7974 4727 7988
rect 4653 7893 4667 7907
rect 4813 7933 4827 7947
rect 4733 7893 4747 7907
rect 4633 7872 4647 7886
rect 4693 7873 4707 7887
rect 4813 7873 4827 7887
rect 4613 7813 4627 7827
rect 4573 7593 4587 7607
rect 4493 7313 4507 7327
rect 4553 7313 4567 7327
rect 4713 7833 4727 7847
rect 4813 7833 4827 7847
rect 4653 7773 4667 7787
rect 4793 7733 4807 7747
rect 4753 7674 4767 7688
rect 4733 7632 4747 7646
rect 4813 7632 4827 7646
rect 4693 7593 4707 7607
rect 4653 7573 4667 7587
rect 4753 7553 4767 7567
rect 4633 7513 4647 7527
rect 4713 7513 4727 7527
rect 4653 7493 4667 7507
rect 4633 7453 4647 7467
rect 4793 7493 4807 7507
rect 4673 7413 4687 7427
rect 4653 7373 4667 7387
rect 4633 7333 4647 7347
rect 4733 7412 4747 7426
rect 4692 7353 4706 7367
rect 4713 7353 4727 7367
rect 4673 7273 4687 7287
rect 4453 7233 4467 7247
rect 4613 7233 4627 7247
rect 4473 7213 4487 7227
rect 4413 7173 4427 7187
rect 4453 7173 4467 7187
rect 4153 7133 4167 7147
rect 4153 7013 4167 7027
rect 4073 6853 4087 6867
rect 4053 6733 4067 6747
rect 4053 6633 4067 6647
rect 4073 6612 4087 6626
rect 4133 6873 4147 6887
rect 4193 6953 4207 6967
rect 4133 6753 4147 6767
rect 4013 6533 4027 6547
rect 4073 6473 4087 6487
rect 3973 6433 3987 6447
rect 4133 6573 4147 6587
rect 4133 6513 4147 6527
rect 4133 6453 4147 6467
rect 3953 6414 3967 6428
rect 3993 6413 4007 6427
rect 4053 6414 4067 6428
rect 4093 6414 4107 6428
rect 4153 6414 4167 6428
rect 3933 6273 3947 6287
rect 3893 6072 3907 6086
rect 3793 5753 3807 5767
rect 3713 5733 3727 5747
rect 3833 5693 3847 5707
rect 3713 5613 3727 5627
rect 3673 5413 3687 5427
rect 3713 5374 3727 5388
rect 3753 5374 3767 5388
rect 3813 5373 3827 5387
rect 3773 5332 3787 5346
rect 3753 5313 3767 5327
rect 3733 5233 3747 5247
rect 3633 5074 3647 5088
rect 3613 5032 3627 5046
rect 3633 4993 3647 5007
rect 3613 4613 3627 4627
rect 3573 4593 3587 4607
rect 3593 4554 3607 4568
rect 3573 4512 3587 4526
rect 3613 4493 3627 4507
rect 3793 5293 3807 5307
rect 3773 5273 3787 5287
rect 3773 5173 3787 5187
rect 3753 4913 3767 4927
rect 3713 4854 3727 4868
rect 3753 4854 3767 4868
rect 3753 4834 3767 4848
rect 3693 4812 3707 4826
rect 3733 4813 3747 4827
rect 3653 4773 3667 4787
rect 3693 4713 3707 4727
rect 3653 4693 3667 4707
rect 3673 4673 3687 4687
rect 3653 4593 3667 4607
rect 3653 4554 3667 4568
rect 3513 4473 3527 4487
rect 3593 4473 3607 4487
rect 3633 4473 3647 4487
rect 3493 4413 3507 4427
rect 3553 4393 3567 4407
rect 3453 4334 3467 4348
rect 3493 4334 3507 4348
rect 3453 4273 3467 4287
rect 3433 4133 3447 4147
rect 3413 4093 3427 4107
rect 3473 4213 3487 4227
rect 3473 4133 3487 4147
rect 3453 4073 3467 4087
rect 3513 4073 3527 4087
rect 3473 4053 3487 4067
rect 3413 3992 3427 4006
rect 3393 3973 3407 3987
rect 3373 3873 3387 3887
rect 3433 3933 3447 3947
rect 3393 3853 3407 3867
rect 3353 3833 3367 3847
rect 3333 3814 3347 3828
rect 3373 3814 3387 3828
rect 3453 3893 3467 3907
rect 3453 3853 3467 3867
rect 3313 3773 3327 3787
rect 3353 3772 3367 3786
rect 3393 3772 3407 3786
rect 3453 3772 3467 3786
rect 3293 3693 3307 3707
rect 3273 3633 3287 3647
rect 3453 3733 3467 3747
rect 3373 3693 3387 3707
rect 3353 3673 3367 3687
rect 3353 3633 3367 3647
rect 3273 3573 3287 3587
rect 3233 3553 3247 3567
rect 3313 3514 3327 3528
rect 3253 3453 3267 3467
rect 3253 3413 3267 3427
rect 3233 3353 3247 3367
rect 3233 3252 3247 3266
rect 3213 3093 3227 3107
rect 3173 2994 3187 3008
rect 3213 2993 3227 3007
rect 3153 2952 3167 2966
rect 3193 2952 3207 2966
rect 3153 2893 3167 2907
rect 3193 2893 3207 2907
rect 3093 2773 3107 2787
rect 3133 2773 3147 2787
rect 3013 2733 3027 2747
rect 3073 2732 3087 2746
rect 3113 2733 3127 2747
rect 3093 2693 3107 2707
rect 3073 2653 3087 2667
rect 2993 2593 3007 2607
rect 3033 2593 3047 2607
rect 2893 2513 2907 2527
rect 2933 2474 2947 2488
rect 2893 2453 2907 2467
rect 2953 2432 2967 2446
rect 3013 2553 3027 2567
rect 2933 2413 2947 2427
rect 2893 2254 2907 2268
rect 2953 2353 2967 2367
rect 2953 2253 2967 2267
rect 2913 2212 2927 2226
rect 2933 2153 2947 2167
rect 2833 2053 2847 2067
rect 2873 2053 2887 2067
rect 2793 2033 2807 2047
rect 2833 1954 2847 1968
rect 2953 2033 2967 2047
rect 2853 1912 2867 1926
rect 2813 1893 2827 1907
rect 2773 1793 2787 1807
rect 2953 1913 2967 1927
rect 2893 1773 2907 1787
rect 2933 1773 2947 1787
rect 2853 1734 2867 1748
rect 2913 1734 2927 1748
rect 2793 1692 2807 1706
rect 2753 1553 2767 1567
rect 2753 1434 2767 1448
rect 2873 1673 2887 1687
rect 2833 1633 2847 1647
rect 2833 1553 2847 1567
rect 2713 1353 2727 1367
rect 2713 1273 2727 1287
rect 2773 1392 2787 1406
rect 2893 1493 2907 1507
rect 2893 1393 2907 1407
rect 2833 1353 2847 1367
rect 2833 1293 2847 1307
rect 2733 1253 2747 1267
rect 2713 1213 2727 1227
rect 2933 1673 2947 1687
rect 2993 2432 3007 2446
rect 2993 2373 3007 2387
rect 2993 2133 3007 2147
rect 3053 2474 3067 2488
rect 3053 2133 3067 2147
rect 3033 2053 3047 2067
rect 3033 1993 3047 2007
rect 3213 2753 3227 2767
rect 3193 2653 3207 2667
rect 3153 2613 3167 2627
rect 3173 2474 3187 2488
rect 3153 2413 3167 2427
rect 3193 2393 3207 2407
rect 3293 3453 3307 3467
rect 3313 3313 3327 3327
rect 3293 3213 3307 3227
rect 3293 3073 3307 3087
rect 3253 2893 3267 2907
rect 3293 2774 3307 2788
rect 3233 2373 3247 2387
rect 3113 2313 3127 2327
rect 3453 3693 3467 3707
rect 3393 3673 3407 3687
rect 3393 3633 3407 3647
rect 3493 3813 3507 3827
rect 3553 4093 3567 4107
rect 3673 4512 3687 4526
rect 3673 4393 3687 4407
rect 3913 5993 3927 6007
rect 3993 6372 4007 6386
rect 4033 6313 4047 6327
rect 4013 6053 4027 6067
rect 3973 6033 3987 6047
rect 4113 6372 4127 6386
rect 4133 6293 4147 6307
rect 4073 6233 4087 6247
rect 4133 6173 4147 6187
rect 4093 6113 4107 6127
rect 4053 6053 4067 6067
rect 4033 5993 4047 6007
rect 4013 5973 4027 5987
rect 3973 5894 3987 5908
rect 4013 5894 4027 5908
rect 4053 5894 4067 5908
rect 4053 5874 4067 5888
rect 4133 6033 4147 6047
rect 4113 6013 4127 6027
rect 4113 5953 4127 5967
rect 4133 5873 4147 5887
rect 3953 5853 3967 5867
rect 3933 5813 3947 5827
rect 3933 5713 3947 5727
rect 3913 5653 3927 5667
rect 3893 5594 3907 5608
rect 3873 5552 3887 5566
rect 4033 5853 4047 5867
rect 3993 5833 4007 5847
rect 3953 5693 3967 5707
rect 3993 5812 4007 5826
rect 3973 5673 3987 5687
rect 3933 5533 3947 5547
rect 4013 5613 4027 5627
rect 3993 5473 4007 5487
rect 3853 5373 3867 5387
rect 3973 5374 3987 5388
rect 3853 5332 3867 5346
rect 3833 5213 3847 5227
rect 4133 5833 4147 5847
rect 4093 5813 4107 5827
rect 4033 5553 4047 5567
rect 4353 7153 4367 7167
rect 4373 7132 4387 7146
rect 4413 7132 4427 7146
rect 4313 7112 4327 7126
rect 4273 7093 4287 7107
rect 4233 7013 4247 7027
rect 4213 6853 4227 6867
rect 4193 6813 4207 6827
rect 4373 7013 4387 7027
rect 4393 6973 4407 6987
rect 4273 6953 4287 6967
rect 4333 6953 4347 6967
rect 4373 6953 4387 6967
rect 4293 6934 4307 6948
rect 4253 6833 4267 6847
rect 4233 6793 4247 6807
rect 4313 6892 4327 6906
rect 4293 6793 4307 6807
rect 4273 6733 4287 6747
rect 4413 6892 4427 6906
rect 4313 6753 4327 6767
rect 4353 6753 4367 6767
rect 4293 6713 4307 6727
rect 4613 7134 4627 7148
rect 4793 7213 4807 7227
rect 4733 7132 4747 7146
rect 4793 7073 4807 7087
rect 4993 8333 5007 8347
rect 4973 8233 4987 8247
rect 5013 8293 5027 8307
rect 5113 8593 5127 8607
rect 5153 8733 5167 8747
rect 5133 8533 5147 8547
rect 5213 8873 5227 8887
rect 5173 8653 5187 8667
rect 5133 8494 5147 8508
rect 5213 8613 5227 8627
rect 5273 8972 5287 8986
rect 5253 8913 5267 8927
rect 5233 8533 5247 8547
rect 5213 8513 5227 8527
rect 5113 8353 5127 8367
rect 5093 8293 5107 8307
rect 5053 8273 5067 8287
rect 5053 8194 5067 8208
rect 5153 8413 5167 8427
rect 5153 8333 5167 8347
rect 5153 8213 5167 8227
rect 5193 8193 5207 8207
rect 4973 8113 4987 8127
rect 4953 8053 4967 8067
rect 4973 8013 4987 8027
rect 4933 7974 4947 7988
rect 4993 7993 5007 8007
rect 5073 8152 5087 8166
rect 5053 8133 5067 8147
rect 5153 8153 5167 8167
rect 5053 8073 5067 8087
rect 5033 8013 5047 8027
rect 5033 7973 5047 7987
rect 4893 7933 4907 7947
rect 4853 7913 4867 7927
rect 4833 7613 4847 7627
rect 4833 7573 4847 7587
rect 4873 7753 4887 7767
rect 4873 7633 4887 7647
rect 4853 7513 4867 7527
rect 4833 7412 4847 7426
rect 4833 7273 4847 7287
rect 4873 7353 4887 7367
rect 4853 7253 4867 7267
rect 4852 7232 4866 7246
rect 4873 7233 4887 7247
rect 4833 7213 4847 7227
rect 4853 7154 4867 7168
rect 4812 7053 4826 7067
rect 4833 7053 4847 7067
rect 4653 7013 4667 7027
rect 4713 7013 4727 7027
rect 4793 7013 4807 7027
rect 4513 6973 4527 6987
rect 4553 6934 4567 6948
rect 4493 6892 4507 6906
rect 4533 6892 4547 6906
rect 4593 6892 4607 6906
rect 4553 6813 4567 6827
rect 4453 6693 4467 6707
rect 4533 6653 4547 6667
rect 4433 6612 4447 6626
rect 4513 6613 4527 6627
rect 4413 6573 4427 6587
rect 4433 6553 4447 6567
rect 4253 6513 4267 6527
rect 4393 6513 4407 6527
rect 4233 6493 4247 6507
rect 4233 6453 4247 6467
rect 4193 6353 4207 6367
rect 4193 6093 4207 6107
rect 4293 6433 4307 6447
rect 4253 6114 4267 6128
rect 4213 6073 4227 6087
rect 4393 6372 4407 6386
rect 4573 6713 4587 6727
rect 4733 6973 4747 6987
rect 4833 6993 4847 7007
rect 4693 6953 4707 6967
rect 4813 6953 4827 6967
rect 4753 6934 4767 6948
rect 4693 6892 4707 6906
rect 4733 6892 4747 6906
rect 4773 6892 4787 6906
rect 4693 6853 4707 6867
rect 4653 6693 4667 6707
rect 4853 6933 4867 6947
rect 4873 6833 4887 6847
rect 4833 6813 4847 6827
rect 4833 6773 4847 6787
rect 4753 6693 4767 6707
rect 4693 6634 4707 6648
rect 4733 6634 4747 6648
rect 4673 6592 4687 6606
rect 4573 6433 4587 6447
rect 4593 6414 4607 6428
rect 4633 6414 4647 6428
rect 4493 6393 4507 6407
rect 4573 6372 4587 6386
rect 4433 6313 4447 6327
rect 4533 6313 4547 6327
rect 4573 6313 4587 6327
rect 4353 6273 4367 6287
rect 4393 6253 4407 6267
rect 4173 6033 4187 6047
rect 4313 6033 4327 6047
rect 4293 5813 4307 5827
rect 4293 5753 4307 5767
rect 4233 5733 4247 5747
rect 4193 5713 4207 5727
rect 4193 5633 4207 5647
rect 4173 5593 4187 5607
rect 4073 5533 4087 5547
rect 4113 5533 4127 5547
rect 4153 5533 4167 5547
rect 4033 5513 4047 5527
rect 4033 5393 4047 5407
rect 4093 5374 4107 5388
rect 4013 5293 4027 5307
rect 4073 5293 4087 5307
rect 3953 5193 3967 5207
rect 3853 5153 3867 5167
rect 3813 5073 3827 5087
rect 4093 5133 4107 5147
rect 3873 5032 3887 5046
rect 4153 5374 4167 5388
rect 4253 5594 4267 5608
rect 4293 5594 4307 5608
rect 4333 5594 4347 5608
rect 4233 5413 4247 5427
rect 4173 5332 4187 5346
rect 4213 5313 4227 5327
rect 4312 5533 4326 5547
rect 4333 5533 4347 5547
rect 4313 5413 4327 5427
rect 4113 4993 4127 5007
rect 4193 5074 4207 5088
rect 4053 4973 4067 4987
rect 3833 4953 3847 4967
rect 4093 4913 4107 4927
rect 3813 4873 3827 4887
rect 3853 4873 3867 4887
rect 3793 4753 3807 4767
rect 3833 4733 3847 4747
rect 3733 4693 3747 4707
rect 3753 4673 3767 4687
rect 3733 4653 3747 4667
rect 3813 4573 3827 4587
rect 3773 4512 3787 4526
rect 3793 4473 3807 4487
rect 3753 4393 3767 4407
rect 3693 4353 3707 4367
rect 3733 4353 3747 4367
rect 3673 4333 3687 4347
rect 3693 4292 3707 4306
rect 3733 4273 3747 4287
rect 3633 4253 3647 4267
rect 3593 4053 3607 4067
rect 3713 4173 3727 4187
rect 3673 4053 3687 4067
rect 3693 4033 3707 4047
rect 3553 3993 3567 4007
rect 3653 3992 3667 4006
rect 3633 3973 3647 3987
rect 3613 3933 3627 3947
rect 3533 3913 3547 3927
rect 3513 3753 3527 3767
rect 3493 3733 3507 3747
rect 3653 3814 3667 3828
rect 3553 3772 3567 3786
rect 3593 3772 3607 3786
rect 3633 3772 3647 3786
rect 3673 3772 3687 3786
rect 3533 3673 3547 3687
rect 3693 3693 3707 3707
rect 3473 3593 3487 3607
rect 3433 3573 3447 3587
rect 3493 3553 3507 3567
rect 3673 3653 3687 3667
rect 3673 3593 3687 3607
rect 3613 3573 3627 3587
rect 3533 3513 3547 3527
rect 3593 3513 3607 3527
rect 3393 3453 3407 3467
rect 3433 3453 3447 3467
rect 3513 3472 3527 3486
rect 3733 4133 3747 4147
rect 3733 3993 3747 4007
rect 3773 4313 3787 4327
rect 3773 4213 3787 4227
rect 3773 4033 3787 4047
rect 3753 3913 3767 3927
rect 3733 3814 3747 3828
rect 3733 3773 3747 3787
rect 3713 3653 3727 3667
rect 3653 3553 3667 3567
rect 3693 3553 3707 3567
rect 3613 3473 3627 3487
rect 3633 3453 3647 3467
rect 3353 3313 3367 3327
rect 3413 3294 3427 3308
rect 3333 3233 3347 3247
rect 3373 3233 3387 3247
rect 3393 3013 3407 3027
rect 3513 3333 3527 3347
rect 3473 3294 3487 3308
rect 3453 3273 3467 3287
rect 3453 3213 3467 3227
rect 3633 3333 3647 3347
rect 3673 3473 3687 3487
rect 3733 3393 3747 3407
rect 3733 3313 3747 3327
rect 3553 3294 3567 3308
rect 3613 3294 3627 3308
rect 3533 3253 3547 3267
rect 3472 3113 3486 3127
rect 3493 3113 3507 3127
rect 3433 2973 3447 2987
rect 3333 2773 3347 2787
rect 3313 2673 3327 2687
rect 3273 2613 3287 2627
rect 3333 2593 3347 2607
rect 3413 2833 3427 2847
rect 3273 2433 3287 2447
rect 3513 2774 3527 2788
rect 3473 2713 3487 2727
rect 3453 2673 3467 2687
rect 3433 2553 3447 2567
rect 3413 2513 3427 2527
rect 3373 2474 3387 2488
rect 3413 2474 3427 2488
rect 3333 2393 3347 2407
rect 3293 2313 3307 2327
rect 3273 2293 3287 2307
rect 3153 2254 3167 2268
rect 3253 2254 3267 2268
rect 3093 2213 3107 2227
rect 3133 2212 3147 2226
rect 3093 2153 3107 2167
rect 3213 2113 3227 2127
rect 3173 2093 3187 2107
rect 3113 2053 3127 2067
rect 3073 1993 3087 2007
rect 3153 1993 3167 2007
rect 3093 1954 3107 1968
rect 3073 1873 3087 1887
rect 3013 1833 3027 1847
rect 3113 1813 3127 1827
rect 3073 1793 3087 1807
rect 3033 1734 3047 1748
rect 3033 1673 3047 1687
rect 2973 1593 2987 1607
rect 2993 1473 3007 1487
rect 3093 1673 3107 1687
rect 3073 1653 3087 1667
rect 3053 1613 3067 1627
rect 3093 1573 3107 1587
rect 2913 1153 2927 1167
rect 2852 993 2866 1007
rect 2873 993 2887 1007
rect 2733 913 2747 927
rect 2813 913 2827 927
rect 2713 872 2727 886
rect 2793 873 2807 887
rect 2753 773 2767 787
rect 2693 713 2707 727
rect 2733 713 2747 727
rect 2833 872 2847 886
rect 2833 713 2847 727
rect 2672 652 2686 666
rect 2693 652 2707 666
rect 2733 652 2747 666
rect 2673 593 2687 607
rect 2673 533 2687 547
rect 2733 533 2747 547
rect 2333 352 2347 366
rect 2393 352 2407 366
rect 2473 352 2487 366
rect 2433 333 2447 347
rect 2653 352 2667 366
rect 2653 293 2667 307
rect 2613 273 2627 287
rect 2293 213 2307 227
rect 2393 213 2407 227
rect 2553 174 2567 188
rect 2613 174 2627 188
rect 2813 653 2827 667
rect 2773 493 2787 507
rect 2813 433 2827 447
rect 2793 413 2807 427
rect 2733 154 2747 168
rect 2413 132 2427 146
rect 2553 133 2567 147
rect 2633 132 2647 146
rect 2713 132 2727 146
rect 2093 113 2107 127
rect 2593 113 2607 127
rect 3033 1434 3047 1448
rect 3013 1392 3027 1406
rect 3013 1313 3027 1327
rect 2993 1273 3007 1287
rect 2973 1214 2987 1228
rect 2973 1113 2987 1127
rect 3233 2053 3247 2067
rect 3213 2033 3227 2047
rect 3193 1873 3207 1887
rect 3173 1734 3187 1748
rect 3153 1673 3167 1687
rect 3153 1573 3167 1587
rect 3133 1273 3147 1287
rect 3053 1214 3067 1228
rect 3093 1214 3107 1228
rect 3013 1193 3027 1207
rect 3033 1172 3047 1186
rect 3073 1172 3087 1186
rect 3113 1172 3127 1186
rect 2993 1053 3007 1067
rect 3033 1053 3047 1067
rect 3033 1013 3047 1027
rect 3073 933 3087 947
rect 3113 913 3127 927
rect 2973 713 2987 727
rect 2933 694 2947 708
rect 3013 694 3027 708
rect 2993 652 3007 666
rect 3113 773 3127 787
rect 3093 713 3107 727
rect 3113 652 3127 666
rect 3033 613 3047 627
rect 3073 613 3087 627
rect 3053 473 3067 487
rect 3093 473 3107 487
rect 2853 453 2867 467
rect 2913 394 2927 408
rect 2793 293 2807 307
rect 2833 352 2847 366
rect 2873 352 2887 366
rect 2813 213 2827 227
rect 2853 333 2867 347
rect 2853 293 2867 307
rect 2873 213 2887 227
rect 2833 174 2847 188
rect 2913 174 2927 188
rect 3433 2433 3447 2447
rect 3393 2293 3407 2307
rect 3413 2273 3427 2287
rect 3353 2254 3367 2268
rect 3293 2213 3307 2227
rect 3333 2212 3347 2226
rect 3273 2173 3287 2187
rect 3373 2173 3387 2187
rect 3273 2113 3287 2127
rect 3413 2093 3427 2107
rect 3253 1993 3267 2007
rect 3253 1954 3267 1968
rect 3313 1954 3327 1968
rect 3233 1913 3247 1927
rect 3333 1912 3347 1926
rect 3373 1913 3387 1927
rect 3293 1793 3307 1807
rect 3253 1734 3267 1748
rect 3493 2673 3507 2687
rect 3473 2553 3487 2567
rect 3473 2393 3487 2407
rect 3473 2253 3487 2267
rect 3473 2213 3487 2227
rect 3513 2453 3527 2467
rect 3513 2273 3527 2287
rect 3653 3293 3667 3307
rect 3713 3293 3727 3307
rect 3593 3252 3607 3266
rect 3573 3173 3587 3187
rect 3613 3233 3627 3247
rect 3553 3133 3567 3147
rect 3593 3133 3607 3147
rect 3613 3113 3627 3127
rect 3553 3013 3567 3027
rect 3673 3252 3687 3266
rect 3713 3073 3727 3087
rect 3573 2994 3587 3008
rect 3633 2994 3647 3008
rect 3693 3013 3707 3027
rect 3673 2992 3687 3006
rect 3593 2952 3607 2966
rect 3653 2953 3667 2967
rect 3613 2873 3627 2887
rect 3553 2753 3567 2767
rect 3613 2653 3627 2667
rect 3673 2913 3687 2927
rect 3693 2813 3707 2827
rect 3733 2893 3747 2907
rect 3813 4353 3827 4367
rect 4013 4833 4027 4847
rect 3993 4793 4007 4807
rect 4013 4773 4027 4787
rect 3913 4693 3927 4707
rect 4033 4693 4047 4707
rect 3853 4453 3867 4467
rect 3893 4413 3907 4427
rect 3933 4673 3947 4687
rect 3993 4653 4007 4667
rect 3953 4613 3967 4627
rect 4033 4573 4047 4587
rect 4053 4554 4067 4568
rect 3953 4512 3967 4526
rect 3993 4512 4007 4526
rect 3933 4473 3947 4487
rect 4013 4473 4027 4487
rect 3913 4393 3927 4407
rect 3893 4334 3907 4348
rect 3953 4334 3967 4348
rect 3993 4334 4007 4348
rect 3853 4273 3867 4287
rect 3933 4273 3947 4287
rect 3813 4233 3827 4247
rect 3833 4193 3847 4207
rect 3973 4253 3987 4267
rect 3953 4213 3967 4227
rect 3853 4173 3867 4187
rect 3853 4034 3867 4048
rect 3873 3992 3887 4006
rect 3913 3992 3927 4006
rect 3813 3973 3827 3987
rect 3853 3973 3867 3987
rect 3793 3893 3807 3907
rect 3893 3853 3907 3867
rect 3853 3833 3867 3847
rect 3833 3772 3847 3786
rect 3773 3453 3787 3467
rect 3833 3693 3847 3707
rect 3953 3953 3967 3967
rect 3933 3893 3947 3907
rect 3913 3693 3927 3707
rect 3873 3553 3887 3567
rect 3953 3873 3967 3887
rect 3993 4213 4007 4227
rect 3993 4073 4007 4087
rect 3993 4013 4007 4027
rect 3993 3992 4007 4006
rect 3973 3753 3987 3767
rect 3933 3533 3947 3547
rect 3873 3453 3887 3467
rect 3913 3453 3927 3467
rect 3933 3433 3947 3447
rect 3873 3393 3887 3407
rect 3853 3252 3867 3266
rect 3833 3193 3847 3207
rect 3793 3173 3807 3187
rect 3833 3093 3847 3107
rect 3913 3233 3927 3247
rect 3873 3173 3887 3187
rect 3893 3153 3907 3167
rect 3873 3133 3887 3147
rect 3853 3053 3867 3067
rect 3813 2933 3827 2947
rect 3753 2833 3767 2847
rect 3673 2633 3687 2647
rect 3653 2573 3667 2587
rect 3613 2474 3627 2488
rect 3633 2393 3647 2407
rect 3553 2333 3567 2347
rect 3593 2333 3607 2347
rect 3593 2273 3607 2287
rect 3593 2254 3607 2268
rect 3533 2173 3547 2187
rect 3492 2113 3506 2127
rect 3513 2113 3527 2127
rect 3473 1993 3487 2007
rect 3453 1953 3467 1967
rect 3433 1913 3447 1927
rect 3413 1873 3427 1887
rect 3393 1773 3407 1787
rect 3613 2213 3627 2227
rect 3573 1993 3587 2007
rect 3553 1912 3567 1926
rect 3553 1873 3567 1887
rect 3493 1853 3507 1867
rect 3593 1833 3607 1847
rect 3553 1813 3567 1827
rect 3413 1733 3427 1747
rect 3553 1773 3567 1787
rect 3553 1733 3567 1747
rect 3273 1692 3287 1706
rect 3373 1693 3387 1707
rect 3533 1692 3547 1706
rect 3573 1692 3587 1706
rect 3493 1673 3507 1687
rect 3533 1653 3547 1667
rect 3413 1553 3427 1567
rect 3473 1553 3487 1567
rect 3413 1473 3427 1487
rect 3213 1453 3227 1467
rect 3253 1453 3267 1467
rect 3393 1413 3407 1427
rect 3173 1393 3187 1407
rect 3173 1333 3187 1347
rect 3193 1293 3207 1307
rect 3193 1172 3207 1186
rect 3273 1392 3287 1406
rect 3353 1373 3367 1387
rect 3253 1213 3267 1227
rect 3313 1214 3327 1228
rect 3393 1213 3407 1227
rect 3253 1172 3267 1186
rect 3293 1172 3307 1186
rect 3333 1073 3347 1087
rect 3233 1053 3247 1067
rect 3233 933 3247 947
rect 3273 914 3287 928
rect 3573 1553 3587 1567
rect 3553 1513 3567 1527
rect 3553 1453 3567 1467
rect 3453 1392 3467 1406
rect 3593 1433 3607 1447
rect 3593 1393 3607 1407
rect 3593 1372 3607 1386
rect 3573 1293 3587 1307
rect 3653 2254 3667 2268
rect 3653 2173 3667 2187
rect 3693 2293 3707 2307
rect 3693 2212 3707 2226
rect 3693 2153 3707 2167
rect 3693 2113 3707 2127
rect 3673 2093 3687 2107
rect 3673 1953 3687 1967
rect 3793 2733 3807 2747
rect 3753 2693 3767 2707
rect 3853 2773 3867 2787
rect 3813 2693 3827 2707
rect 3873 2753 3887 2767
rect 3853 2613 3867 2627
rect 3793 2593 3807 2607
rect 3753 2573 3767 2587
rect 3873 2513 3887 2527
rect 3813 2474 3827 2488
rect 3873 2473 3887 2487
rect 3793 2432 3807 2446
rect 3753 2373 3767 2387
rect 3833 2373 3847 2387
rect 3773 2333 3787 2347
rect 3813 2254 3827 2268
rect 3733 2233 3747 2247
rect 3793 2212 3807 2226
rect 3833 2212 3847 2226
rect 3733 2133 3747 2147
rect 3713 2073 3727 2087
rect 3773 2053 3787 2067
rect 3952 3393 3966 3407
rect 3973 3393 3987 3407
rect 3973 3313 3987 3327
rect 4033 4133 4047 4147
rect 4313 5193 4327 5207
rect 4253 5153 4267 5167
rect 4293 5074 4307 5088
rect 4693 6513 4707 6527
rect 4693 6433 4707 6447
rect 4713 6413 4727 6427
rect 4673 6372 4687 6386
rect 4653 6333 4667 6347
rect 4633 6193 4647 6207
rect 4593 6173 4607 6187
rect 4453 6114 4467 6128
rect 4553 6113 4567 6127
rect 4433 6072 4447 6086
rect 4553 6072 4567 6086
rect 4573 5973 4587 5987
rect 4413 5874 4427 5888
rect 4513 5874 4527 5888
rect 4573 5853 4587 5867
rect 4573 5832 4587 5846
rect 4573 5673 4587 5687
rect 4713 6133 4727 6147
rect 4633 6072 4647 6086
rect 4693 6053 4707 6067
rect 4673 6033 4687 6047
rect 4613 5993 4627 6007
rect 4593 5633 4607 5647
rect 4553 5594 4567 5608
rect 4393 5533 4407 5547
rect 4433 5513 4447 5527
rect 4413 5473 4427 5487
rect 4373 5413 4387 5427
rect 4353 5373 4367 5387
rect 4433 5393 4447 5407
rect 4433 5293 4447 5307
rect 4533 5552 4547 5566
rect 4573 5533 4587 5547
rect 4573 5453 4587 5467
rect 4553 5413 4567 5427
rect 4533 5353 4547 5367
rect 4513 5332 4527 5346
rect 4553 5333 4567 5347
rect 4393 5233 4407 5247
rect 4473 5233 4487 5247
rect 4373 5213 4387 5227
rect 4373 5153 4387 5167
rect 4393 5113 4407 5127
rect 4473 5074 4487 5088
rect 4273 5032 4287 5046
rect 4333 5033 4347 5047
rect 4493 5032 4507 5046
rect 4553 5073 4567 5087
rect 4213 4873 4227 4887
rect 4193 4833 4207 4847
rect 4113 4773 4127 4787
rect 4153 4713 4167 4727
rect 4213 4713 4227 4727
rect 4373 4832 4387 4846
rect 4273 4593 4287 4607
rect 4433 4593 4447 4607
rect 4493 4593 4507 4607
rect 4133 4554 4147 4568
rect 4233 4554 4247 4568
rect 4193 4533 4207 4547
rect 4133 4513 4147 4527
rect 4253 4512 4267 4526
rect 4193 4473 4207 4487
rect 4333 4433 4347 4447
rect 4233 4393 4247 4407
rect 4113 4333 4127 4347
rect 4153 4334 4167 4348
rect 4193 4334 4207 4348
rect 4113 4133 4127 4147
rect 4093 4073 4107 4087
rect 4053 4034 4067 4048
rect 4073 3992 4087 4006
rect 4013 3933 4027 3947
rect 4033 3893 4047 3907
rect 4013 3873 4027 3887
rect 4053 3833 4067 3847
rect 4013 3813 4027 3827
rect 4173 4292 4187 4306
rect 4433 4393 4447 4407
rect 4373 4334 4387 4348
rect 4413 4334 4427 4348
rect 4453 4334 4467 4348
rect 4433 4293 4447 4307
rect 4433 4233 4447 4247
rect 4333 4193 4347 4207
rect 4413 4173 4427 4187
rect 4133 4093 4147 4107
rect 4193 4093 4207 4107
rect 4233 4093 4247 4107
rect 4133 3933 4147 3947
rect 4113 3813 4127 3827
rect 3993 3153 4007 3167
rect 3933 3113 3947 3127
rect 3993 3093 4007 3107
rect 3993 3053 4007 3067
rect 3973 2994 3987 3008
rect 3933 2952 3947 2966
rect 3913 2933 3927 2947
rect 3953 2913 3967 2927
rect 3973 2853 3987 2867
rect 4113 3773 4127 3787
rect 4033 3533 4047 3547
rect 4053 3493 4067 3507
rect 4033 3294 4047 3308
rect 4193 3773 4207 3787
rect 4253 4034 4267 4048
rect 4352 4033 4366 4047
rect 4373 4033 4387 4047
rect 4273 3992 4287 4006
rect 4373 3992 4387 4006
rect 4413 3993 4427 4007
rect 4413 3953 4427 3967
rect 4313 3913 4327 3927
rect 4353 3913 4367 3927
rect 4273 3814 4287 3828
rect 4413 3893 4427 3907
rect 4353 3814 4367 3828
rect 4253 3753 4267 3767
rect 4133 3733 4147 3747
rect 4233 3514 4247 3528
rect 4353 3773 4367 3787
rect 4293 3733 4307 3747
rect 4473 4293 4487 4307
rect 4793 6673 4807 6687
rect 4773 6634 4787 6648
rect 4813 6653 4827 6667
rect 4793 6593 4807 6607
rect 5013 7933 5027 7947
rect 5053 7953 5067 7967
rect 4953 7813 4967 7827
rect 4933 7613 4947 7627
rect 4973 7593 4987 7607
rect 4953 7573 4967 7587
rect 5033 7812 5047 7826
rect 5073 7932 5087 7946
rect 5073 7773 5087 7787
rect 5053 7753 5067 7767
rect 4993 7513 5007 7527
rect 5033 7453 5047 7467
rect 5193 8113 5207 8127
rect 5133 8053 5147 8067
rect 5173 8033 5187 8047
rect 5133 7974 5147 7988
rect 5173 7974 5187 7988
rect 5153 7932 5167 7946
rect 5173 7913 5187 7927
rect 5172 7873 5186 7887
rect 5193 7873 5207 7887
rect 5213 7853 5227 7867
rect 5133 7793 5147 7807
rect 5113 7773 5127 7787
rect 5133 7713 5147 7727
rect 5113 7674 5127 7688
rect 5093 7553 5107 7567
rect 5073 7513 5087 7527
rect 4993 7412 5007 7426
rect 5033 7412 5047 7426
rect 5033 7333 5047 7347
rect 4913 7193 4927 7207
rect 5053 7313 5067 7327
rect 5053 7273 5067 7287
rect 4993 7253 5007 7267
rect 5033 7253 5047 7267
rect 5033 7154 5047 7168
rect 4933 7133 4947 7147
rect 5013 7112 5027 7126
rect 4913 7093 4927 7107
rect 4973 7093 4987 7107
rect 4933 7073 4947 7087
rect 5033 7073 5047 7087
rect 4933 6993 4947 7007
rect 4953 6973 4967 6987
rect 5053 7053 5067 7067
rect 5033 6953 5047 6967
rect 5093 7313 5107 7327
rect 5093 7133 5107 7147
rect 5073 6993 5087 7007
rect 4993 6934 5007 6948
rect 5053 6933 5067 6947
rect 4913 6892 4927 6906
rect 4893 6753 4907 6767
rect 4933 6713 4947 6727
rect 4893 6693 4907 6707
rect 4893 6634 4907 6648
rect 5013 6873 5027 6887
rect 5013 6833 5027 6847
rect 5013 6793 5027 6807
rect 5013 6753 5027 6767
rect 4833 6592 4847 6606
rect 4873 6592 4887 6606
rect 4913 6592 4927 6606
rect 4973 6593 4987 6607
rect 5013 6593 5027 6607
rect 5013 6572 5027 6586
rect 4813 6553 4827 6567
rect 4993 6533 5007 6547
rect 4833 6513 4847 6527
rect 4773 6353 4787 6367
rect 4773 6293 4787 6307
rect 4753 6233 4767 6247
rect 4793 6093 4807 6107
rect 4773 5993 4787 6007
rect 4733 5933 4747 5947
rect 4733 5894 4747 5908
rect 4773 5894 4787 5908
rect 4633 5853 4647 5867
rect 4673 5852 4687 5866
rect 4653 5793 4667 5807
rect 4713 5753 4727 5767
rect 4673 5533 4687 5547
rect 4633 5453 4647 5467
rect 4613 5413 4627 5427
rect 4813 6013 4827 6027
rect 4813 5713 4827 5727
rect 4793 5653 4807 5667
rect 4773 5533 4787 5547
rect 4873 6393 4887 6407
rect 4913 6353 4927 6367
rect 4913 6273 4927 6287
rect 4953 6233 4967 6247
rect 4913 6133 4927 6147
rect 5013 6273 5027 6287
rect 4993 6173 5007 6187
rect 4993 6114 5007 6128
rect 4933 5973 4947 5987
rect 4893 5953 4907 5967
rect 4933 5952 4947 5966
rect 4993 5953 5007 5967
rect 4973 5894 4987 5908
rect 5013 5892 5027 5906
rect 4913 5852 4927 5866
rect 4953 5753 4967 5767
rect 4893 5593 4907 5607
rect 4933 5594 4947 5608
rect 5013 5753 5027 5767
rect 5053 6873 5067 6887
rect 5053 6753 5067 6767
rect 5053 6732 5067 6746
rect 5073 6713 5087 6727
rect 5153 7632 5167 7646
rect 5193 7633 5207 7647
rect 5293 8953 5307 8967
rect 5273 8833 5287 8847
rect 5453 9453 5467 9467
rect 5453 9393 5467 9407
rect 5433 9253 5447 9267
rect 5432 9193 5446 9207
rect 5493 9373 5507 9387
rect 5453 9192 5467 9206
rect 5653 10313 5667 10327
rect 5573 10274 5587 10288
rect 5613 10274 5627 10288
rect 5593 10233 5607 10247
rect 5573 10093 5587 10107
rect 5573 10054 5587 10068
rect 5553 9953 5567 9967
rect 5553 9833 5567 9847
rect 5533 9333 5547 9347
rect 5653 10054 5667 10068
rect 5713 10273 5727 10287
rect 5853 11094 5867 11108
rect 5873 10794 5887 10808
rect 5793 10713 5807 10727
rect 5853 10673 5867 10687
rect 5813 10613 5827 10627
rect 5853 10574 5867 10588
rect 5793 10532 5807 10546
rect 5933 11094 5947 11108
rect 5913 10953 5927 10967
rect 5793 10413 5807 10427
rect 5773 10393 5787 10407
rect 5733 10233 5747 10247
rect 5733 10054 5747 10068
rect 5593 9673 5607 9687
rect 5713 9993 5727 10007
rect 5673 9953 5687 9967
rect 5833 10353 5847 10367
rect 5793 10313 5807 10327
rect 5773 9973 5787 9987
rect 5753 9853 5767 9867
rect 5733 9793 5747 9807
rect 5693 9773 5707 9787
rect 5673 9754 5687 9768
rect 5713 9712 5727 9726
rect 5653 9653 5667 9667
rect 5653 9573 5667 9587
rect 5713 9553 5727 9567
rect 5573 9393 5587 9407
rect 5553 9293 5567 9307
rect 5493 9234 5507 9248
rect 5653 9534 5667 9548
rect 5693 9534 5707 9548
rect 5633 9492 5647 9506
rect 5653 9433 5667 9447
rect 5593 9273 5607 9287
rect 5633 9273 5647 9287
rect 5593 9252 5607 9266
rect 5473 9173 5487 9187
rect 5393 9153 5407 9167
rect 5453 9153 5467 9167
rect 5353 9093 5367 9107
rect 5393 9033 5407 9047
rect 5393 9014 5407 9028
rect 5373 8972 5387 8986
rect 5353 8953 5367 8967
rect 5413 8773 5427 8787
rect 5313 8613 5327 8627
rect 5353 8613 5367 8627
rect 5273 8553 5287 8567
rect 5253 8393 5267 8407
rect 5293 8473 5307 8487
rect 5273 8373 5287 8387
rect 5353 8573 5367 8587
rect 5433 8714 5447 8728
rect 5393 8653 5407 8667
rect 5413 8633 5427 8647
rect 5393 8593 5407 8607
rect 5433 8613 5447 8627
rect 5413 8553 5427 8567
rect 5393 8533 5407 8547
rect 5373 8513 5387 8527
rect 5473 8972 5487 8986
rect 5533 9192 5547 9206
rect 5573 9173 5587 9187
rect 5513 9093 5527 9107
rect 5693 9373 5707 9387
rect 5693 9333 5707 9347
rect 5753 9393 5767 9407
rect 5893 10473 5907 10487
rect 5953 10573 5967 10587
rect 5933 10313 5947 10327
rect 6033 11133 6047 11147
rect 6093 10873 6107 10887
rect 6053 10833 6067 10847
rect 6053 10794 6067 10808
rect 6153 10794 6167 10808
rect 6073 10752 6087 10766
rect 6153 10753 6167 10767
rect 6193 10752 6207 10766
rect 6113 10713 6127 10727
rect 6053 10574 6067 10588
rect 5993 10532 6007 10546
rect 6033 10532 6047 10546
rect 5973 10513 5987 10527
rect 5973 10333 5987 10347
rect 5973 10232 5987 10246
rect 5953 10012 5967 10026
rect 5953 9973 5967 9987
rect 5913 9793 5927 9807
rect 5833 9753 5847 9767
rect 5873 9754 5887 9768
rect 5833 9713 5847 9727
rect 5853 9693 5867 9707
rect 5833 9673 5847 9687
rect 5872 9673 5886 9687
rect 5893 9673 5907 9687
rect 5813 9613 5827 9627
rect 5833 9553 5847 9567
rect 5853 9492 5867 9506
rect 5793 9433 5807 9447
rect 5773 9333 5787 9347
rect 5893 9473 5907 9487
rect 5873 9353 5887 9367
rect 5853 9313 5867 9327
rect 5793 9234 5807 9248
rect 5833 9234 5847 9248
rect 5733 9193 5747 9207
rect 5593 9053 5607 9067
rect 5633 9053 5647 9067
rect 5633 9014 5647 9028
rect 5613 8972 5627 8986
rect 5513 8933 5527 8947
rect 5633 8933 5647 8947
rect 5493 8913 5507 8927
rect 5593 8753 5607 8767
rect 5553 8714 5567 8728
rect 5533 8672 5547 8686
rect 5533 8613 5547 8627
rect 5313 8433 5327 8447
rect 5353 8433 5367 8447
rect 5413 8452 5427 8466
rect 5453 8453 5467 8467
rect 5633 8673 5647 8687
rect 5633 8494 5647 8508
rect 5313 8393 5327 8407
rect 5293 8273 5307 8287
rect 5253 8153 5267 8167
rect 5253 8132 5267 8146
rect 5233 7593 5247 7607
rect 5213 7553 5227 7567
rect 5193 7473 5207 7487
rect 5173 7454 5187 7468
rect 5213 7454 5227 7468
rect 5333 8153 5347 8167
rect 5313 8093 5327 8107
rect 5293 8073 5307 8087
rect 5273 7974 5287 7988
rect 5273 7833 5287 7847
rect 5273 7673 5287 7687
rect 5253 7453 5267 7467
rect 5133 7373 5147 7387
rect 5173 7333 5187 7347
rect 5153 7213 5167 7227
rect 5173 7154 5187 7168
rect 5373 8313 5387 8327
rect 5373 8233 5387 8247
rect 5353 8093 5367 8107
rect 5353 8053 5367 8067
rect 5353 7973 5367 7987
rect 5453 8373 5467 8387
rect 5413 8293 5427 8307
rect 5413 8113 5427 8127
rect 5393 8053 5407 8067
rect 5513 8293 5527 8307
rect 5413 7993 5427 8007
rect 5353 7933 5367 7947
rect 5353 7893 5367 7907
rect 5413 7893 5427 7907
rect 5353 7713 5367 7727
rect 5313 7673 5327 7687
rect 5393 7674 5407 7688
rect 5533 8093 5547 8107
rect 5513 8073 5527 8087
rect 5473 7853 5487 7867
rect 5433 7674 5447 7688
rect 5373 7632 5387 7646
rect 5413 7633 5427 7647
rect 5353 7613 5367 7627
rect 5333 7533 5347 7547
rect 5413 7592 5427 7606
rect 5473 7713 5487 7727
rect 5393 7412 5407 7426
rect 5353 7373 5367 7387
rect 5273 7353 5287 7367
rect 5373 7353 5387 7367
rect 5333 7313 5347 7327
rect 5333 7193 5347 7207
rect 5253 7173 5267 7187
rect 5313 7173 5327 7187
rect 5213 7154 5227 7168
rect 5233 7112 5247 7126
rect 5273 7112 5287 7126
rect 5193 7093 5207 7107
rect 5253 7073 5267 7087
rect 5173 7013 5187 7027
rect 5193 6993 5207 7007
rect 5133 6892 5147 6906
rect 5193 6793 5207 6807
rect 5173 6713 5187 6727
rect 5113 6693 5127 6707
rect 5093 6673 5107 6687
rect 5073 6634 5087 6648
rect 5133 6634 5147 6648
rect 5193 6673 5207 6687
rect 5193 6634 5207 6648
rect 5113 6592 5127 6606
rect 5153 6573 5167 6587
rect 5233 6533 5247 6547
rect 5273 6993 5287 7007
rect 5333 7112 5347 7126
rect 5353 7073 5367 7087
rect 5433 7373 5447 7387
rect 5413 7353 5427 7367
rect 5453 7353 5467 7367
rect 5393 7113 5407 7127
rect 5373 7053 5387 7067
rect 5593 8413 5607 8427
rect 5573 8393 5587 8407
rect 5573 8372 5587 8386
rect 5573 8213 5587 8227
rect 5613 8293 5627 8307
rect 5633 8273 5647 8287
rect 5613 8253 5627 8267
rect 5593 8133 5607 8147
rect 5552 8073 5566 8087
rect 5573 8073 5587 8087
rect 5633 8013 5647 8027
rect 5613 7992 5627 8006
rect 5653 7973 5667 7987
rect 5633 7932 5647 7946
rect 5553 7833 5567 7847
rect 5633 7773 5647 7787
rect 5593 7674 5607 7688
rect 5653 7713 5667 7727
rect 5573 7632 5587 7646
rect 5633 7633 5647 7647
rect 5533 7613 5547 7627
rect 5633 7612 5647 7626
rect 5513 7593 5527 7607
rect 5533 7473 5547 7487
rect 5493 7413 5507 7427
rect 5553 7333 5567 7347
rect 5533 7213 5547 7227
rect 5473 7154 5487 7168
rect 5513 7154 5527 7168
rect 5533 7113 5547 7127
rect 5493 7073 5507 7087
rect 5473 7053 5487 7067
rect 5513 7053 5527 7067
rect 5453 7033 5467 7047
rect 5433 6993 5447 7007
rect 5273 6953 5287 6967
rect 5313 6953 5327 6967
rect 5393 6953 5407 6967
rect 5273 6813 5287 6827
rect 5293 6773 5307 6787
rect 5273 6653 5287 6667
rect 5293 6533 5307 6547
rect 5073 6473 5087 6487
rect 5113 6473 5127 6487
rect 5113 6433 5127 6447
rect 5213 6433 5227 6447
rect 5093 6413 5107 6427
rect 5153 6414 5167 6428
rect 5173 6372 5187 6386
rect 5473 6973 5487 6987
rect 5373 6892 5387 6906
rect 5393 6833 5407 6847
rect 5373 6693 5387 6707
rect 5413 6713 5427 6727
rect 5453 6713 5467 6727
rect 5393 6673 5407 6687
rect 5373 6634 5387 6648
rect 5413 6634 5427 6648
rect 5473 6634 5487 6648
rect 5393 6592 5407 6606
rect 5453 6593 5467 6607
rect 5513 6933 5527 6947
rect 5513 6892 5527 6906
rect 5773 9192 5787 9206
rect 5873 9193 5887 9207
rect 5833 9173 5847 9187
rect 5813 9153 5827 9167
rect 5853 9033 5867 9047
rect 5913 9433 5927 9447
rect 5893 9013 5907 9027
rect 5833 8933 5847 8947
rect 5733 8893 5747 8907
rect 5813 8893 5827 8907
rect 5733 8672 5747 8686
rect 5733 8651 5747 8665
rect 5773 8653 5787 8667
rect 5713 8633 5727 8647
rect 5713 8494 5727 8508
rect 5713 8433 5727 8447
rect 5693 8373 5707 8387
rect 5713 8333 5727 8347
rect 5753 8494 5767 8508
rect 5893 8973 5907 8987
rect 5873 8893 5887 8907
rect 5873 8813 5887 8827
rect 5873 8713 5887 8727
rect 5893 8673 5907 8687
rect 5873 8593 5887 8607
rect 5833 8573 5847 8587
rect 5853 8553 5867 8567
rect 5813 8494 5827 8508
rect 5853 8433 5867 8447
rect 5813 8353 5827 8367
rect 5773 8333 5787 8347
rect 5733 8253 5747 8267
rect 5713 8213 5727 8227
rect 5693 8194 5707 8208
rect 5733 8133 5747 8147
rect 5713 8113 5727 8127
rect 5713 8013 5727 8027
rect 5693 7973 5707 7987
rect 5693 7633 5707 7647
rect 5673 7613 5687 7627
rect 5653 7513 5667 7527
rect 5573 7154 5587 7168
rect 5553 7073 5567 7087
rect 5653 7412 5667 7426
rect 5753 8113 5767 8127
rect 5833 8194 5847 8208
rect 5833 8053 5847 8067
rect 5873 8413 5887 8427
rect 5873 8373 5887 8387
rect 5933 9393 5947 9407
rect 5933 9053 5947 9067
rect 5933 9013 5947 9027
rect 5953 8933 5967 8947
rect 6073 10513 6087 10527
rect 6193 10673 6207 10687
rect 6173 10613 6187 10627
rect 6173 10573 6187 10587
rect 6113 10473 6127 10487
rect 6073 10413 6087 10427
rect 6193 10413 6207 10427
rect 6013 10273 6027 10287
rect 6113 10373 6127 10387
rect 5993 10013 6007 10027
rect 6053 10232 6067 10246
rect 6093 10232 6107 10246
rect 6193 10233 6207 10247
rect 6133 10193 6147 10207
rect 6313 11033 6327 11047
rect 6273 10794 6287 10808
rect 6353 10794 6367 10808
rect 6333 10752 6347 10766
rect 6493 11173 6507 11187
rect 10253 11173 10267 11187
rect 10453 11173 10467 11187
rect 6413 11094 6427 11108
rect 6453 11094 6467 11108
rect 6593 11133 6607 11147
rect 6853 11133 6867 11147
rect 6933 11133 6947 11147
rect 7073 11133 7087 11147
rect 7373 11133 7387 11147
rect 7813 11133 7827 11147
rect 8953 11133 8967 11147
rect 9073 11133 9087 11147
rect 6553 11093 6567 11107
rect 6473 11033 6487 11047
rect 6453 10873 6467 10887
rect 6413 10733 6427 10747
rect 6293 10693 6307 10707
rect 6313 10532 6327 10546
rect 6253 10473 6267 10487
rect 6153 10113 6167 10127
rect 6213 10113 6227 10127
rect 6193 10054 6207 10068
rect 6053 10012 6067 10026
rect 6133 10012 6147 10026
rect 6193 9993 6207 10007
rect 6173 9973 6187 9987
rect 6133 9873 6147 9887
rect 6093 9754 6107 9768
rect 6053 9693 6067 9707
rect 6153 9713 6167 9727
rect 6113 9633 6127 9647
rect 6093 9534 6107 9548
rect 6133 9534 6147 9548
rect 6013 9473 6027 9487
rect 5993 9273 6007 9287
rect 6113 9493 6127 9507
rect 6073 9413 6087 9427
rect 5993 9193 6007 9207
rect 6013 9173 6027 9187
rect 6013 9152 6027 9166
rect 5993 8913 6007 8927
rect 5973 8873 5987 8887
rect 5933 8833 5947 8847
rect 5993 8813 6007 8827
rect 6093 9373 6107 9387
rect 6133 9453 6147 9467
rect 6113 9153 6127 9167
rect 6073 8972 6087 8986
rect 6133 8973 6147 8987
rect 6113 8933 6127 8947
rect 6053 8913 6067 8927
rect 6013 8753 6027 8767
rect 5973 8672 5987 8686
rect 6013 8633 6027 8647
rect 6013 8573 6027 8587
rect 5953 8533 5967 8547
rect 5993 8533 6007 8547
rect 5913 8353 5927 8367
rect 5993 8373 6007 8387
rect 5973 8293 5987 8307
rect 5953 8273 5967 8287
rect 5893 8213 5907 8227
rect 5973 8213 5987 8227
rect 5873 8133 5887 8147
rect 5953 8194 5967 8208
rect 6073 8733 6087 8747
rect 6093 8593 6107 8607
rect 6052 8533 6066 8547
rect 6073 8533 6087 8547
rect 6133 8673 6147 8687
rect 6113 8573 6127 8587
rect 6093 8493 6107 8507
rect 6173 9653 6187 9667
rect 6213 9753 6227 9767
rect 6493 10853 6507 10867
rect 6553 10833 6567 10847
rect 6713 11094 6727 11108
rect 6693 10933 6707 10947
rect 6813 10813 6827 10827
rect 6633 10794 6647 10808
rect 6733 10794 6747 10808
rect 6773 10794 6787 10808
rect 6493 10752 6507 10766
rect 6573 10733 6587 10747
rect 6633 10733 6647 10747
rect 6373 10673 6387 10687
rect 6453 10673 6467 10687
rect 6533 10673 6547 10687
rect 6733 10673 6747 10687
rect 6273 10073 6287 10087
rect 6473 10633 6487 10647
rect 6733 10613 6747 10627
rect 6473 10573 6487 10587
rect 6513 10574 6527 10588
rect 6633 10573 6647 10587
rect 6493 10532 6507 10546
rect 6573 10493 6587 10507
rect 6533 10433 6547 10447
rect 6473 10353 6487 10367
rect 6453 10274 6467 10288
rect 6393 10232 6407 10246
rect 6393 10073 6407 10087
rect 6413 10012 6427 10026
rect 6313 9993 6327 10007
rect 6353 9993 6367 10007
rect 6393 9993 6407 10007
rect 6353 9773 6367 9787
rect 6313 9754 6327 9768
rect 6273 9713 6287 9727
rect 6333 9712 6347 9726
rect 6373 9673 6387 9687
rect 6333 9573 6347 9587
rect 6373 9513 6387 9527
rect 6193 9493 6207 9507
rect 6233 9492 6247 9506
rect 6273 9492 6287 9506
rect 6173 9293 6187 9307
rect 6173 9234 6187 9248
rect 6273 9433 6287 9447
rect 6333 9473 6347 9487
rect 6313 9373 6327 9387
rect 6293 9353 6307 9367
rect 6233 9173 6247 9187
rect 6213 9053 6227 9067
rect 6193 8873 6207 8887
rect 6193 8833 6207 8847
rect 6413 9754 6427 9768
rect 6413 9713 6427 9727
rect 6433 9613 6447 9627
rect 6393 9433 6407 9447
rect 6333 9173 6347 9187
rect 6293 9053 6307 9067
rect 6313 9014 6327 9028
rect 6253 8973 6267 8987
rect 6233 8853 6247 8867
rect 6293 8813 6307 8827
rect 6173 8793 6187 8807
rect 6213 8793 6227 8807
rect 6293 8792 6307 8806
rect 6193 8713 6207 8727
rect 6213 8672 6227 8686
rect 6233 8613 6247 8627
rect 6313 8773 6327 8787
rect 6253 8593 6267 8607
rect 6293 8533 6307 8547
rect 6193 8494 6207 8508
rect 6233 8494 6247 8508
rect 6033 8393 6047 8407
rect 5893 8113 5907 8127
rect 5953 8113 5967 8127
rect 5933 8053 5947 8067
rect 5853 7974 5867 7988
rect 5793 7932 5807 7946
rect 5913 7974 5927 7988
rect 5873 7913 5887 7927
rect 5793 7893 5807 7907
rect 5833 7893 5847 7907
rect 5753 7733 5767 7747
rect 5893 7813 5907 7827
rect 5833 7713 5847 7727
rect 5793 7674 5807 7688
rect 5773 7632 5787 7646
rect 5813 7632 5827 7646
rect 5893 7633 5907 7647
rect 5913 7613 5927 7627
rect 5793 7553 5807 7567
rect 5773 7413 5787 7427
rect 5773 7373 5787 7387
rect 5633 7253 5647 7267
rect 5613 7113 5627 7127
rect 5353 6573 5367 6587
rect 5353 6533 5367 6547
rect 5253 6493 5267 6507
rect 5313 6493 5327 6507
rect 5293 6453 5307 6467
rect 5253 6414 5267 6428
rect 5073 6313 5087 6327
rect 5053 6073 5067 6087
rect 5033 5733 5047 5747
rect 5033 5653 5047 5667
rect 4753 5513 4767 5527
rect 4833 5513 4847 5527
rect 4693 5473 4707 5487
rect 4733 5473 4747 5487
rect 4673 5373 4687 5387
rect 4953 5552 4967 5566
rect 4993 5552 5007 5566
rect 4933 5533 4947 5547
rect 4993 5513 5007 5527
rect 4893 5473 4907 5487
rect 4753 5393 4767 5407
rect 4653 5332 4667 5346
rect 4753 5333 4767 5347
rect 4853 5333 4867 5347
rect 4633 5293 4647 5307
rect 4593 5273 4607 5287
rect 4593 5113 4607 5127
rect 4553 4933 4567 4947
rect 4533 4873 4547 4887
rect 4613 5032 4627 5046
rect 4613 4913 4627 4927
rect 4593 4833 4607 4847
rect 4533 4793 4547 4807
rect 4693 5273 4707 5287
rect 4693 5233 4707 5247
rect 5053 5592 5067 5606
rect 5053 5493 5067 5507
rect 5133 6273 5147 6287
rect 5213 6113 5227 6127
rect 5093 6072 5107 6086
rect 5153 6072 5167 6086
rect 5153 5953 5167 5967
rect 5113 5893 5127 5907
rect 5113 5793 5127 5807
rect 5213 5852 5227 5866
rect 5233 5833 5247 5847
rect 5173 5633 5187 5647
rect 5133 5594 5147 5608
rect 5213 5594 5227 5608
rect 5313 6413 5327 6427
rect 5393 6433 5407 6447
rect 5493 6592 5507 6606
rect 5473 6572 5487 6586
rect 5433 6413 5447 6427
rect 5293 6373 5307 6387
rect 5273 6233 5287 6247
rect 5293 6173 5307 6187
rect 5413 6353 5427 6367
rect 5333 6114 5347 6128
rect 5373 6114 5387 6128
rect 5413 6092 5427 6106
rect 5353 6072 5367 6086
rect 5313 6053 5327 6067
rect 5433 6013 5447 6027
rect 5413 5953 5427 5967
rect 5473 6213 5487 6227
rect 5473 6073 5487 6087
rect 5453 5993 5467 6007
rect 5453 5972 5467 5986
rect 5433 5913 5447 5927
rect 5353 5894 5367 5908
rect 5473 5953 5487 5967
rect 5453 5893 5467 5907
rect 5573 7033 5587 7047
rect 5613 7033 5627 7047
rect 5713 7154 5727 7168
rect 5753 7113 5767 7127
rect 5653 7053 5667 7067
rect 5693 7013 5707 7027
rect 5633 6973 5647 6987
rect 5573 6953 5587 6967
rect 5633 6952 5647 6966
rect 5613 6892 5627 6906
rect 5653 6853 5667 6867
rect 5613 6813 5627 6827
rect 5613 6713 5627 6727
rect 5653 6634 5667 6648
rect 5593 6592 5607 6606
rect 5533 6553 5547 6567
rect 5533 6493 5547 6507
rect 5593 6433 5607 6447
rect 5713 6634 5727 6648
rect 5693 6513 5707 6527
rect 5533 6253 5547 6267
rect 5733 6373 5747 6387
rect 5713 6253 5727 6267
rect 5593 6233 5607 6247
rect 5653 6094 5667 6108
rect 5573 5993 5587 6007
rect 5733 5993 5747 6007
rect 5713 5973 5727 5987
rect 5293 5833 5307 5847
rect 5293 5812 5307 5826
rect 5272 5773 5286 5787
rect 5293 5773 5307 5787
rect 5513 5853 5527 5867
rect 5373 5833 5387 5847
rect 5593 5852 5607 5866
rect 5553 5813 5567 5827
rect 5613 5813 5627 5827
rect 5513 5733 5527 5747
rect 5293 5673 5307 5687
rect 5333 5673 5347 5687
rect 5313 5633 5327 5647
rect 5293 5613 5307 5627
rect 5093 5513 5107 5527
rect 4993 5293 5007 5307
rect 4853 5273 4867 5287
rect 4833 5233 4847 5247
rect 4673 5113 4687 5127
rect 4713 5074 4727 5088
rect 4693 5013 4707 5027
rect 4653 4992 4667 5006
rect 4593 4773 4607 4787
rect 4633 4773 4647 4787
rect 4553 4334 4567 4348
rect 4813 5193 4827 5207
rect 4793 5153 4807 5167
rect 4793 5053 4807 5067
rect 4773 5013 4787 5027
rect 4673 4933 4687 4947
rect 4673 4773 4687 4787
rect 4653 4653 4667 4667
rect 4653 4554 4667 4568
rect 4733 4953 4747 4967
rect 4713 4933 4727 4947
rect 4813 4893 4827 4907
rect 5093 5453 5107 5467
rect 5253 5593 5267 5607
rect 5133 5453 5147 5467
rect 5233 5552 5247 5566
rect 5333 5572 5347 5586
rect 5533 5633 5547 5647
rect 5533 5573 5547 5587
rect 5213 5533 5227 5547
rect 5313 5552 5327 5566
rect 5313 5513 5327 5527
rect 5213 5493 5227 5507
rect 5213 5433 5227 5447
rect 5193 5393 5207 5407
rect 5533 5453 5547 5467
rect 5333 5413 5347 5427
rect 5053 5233 5067 5247
rect 4933 5213 4947 5227
rect 4873 5153 4887 5167
rect 4993 5113 5007 5127
rect 4913 5032 4927 5046
rect 4873 4973 4887 4987
rect 4853 4933 4867 4947
rect 4993 4993 5007 5007
rect 4953 4973 4967 4987
rect 4853 4853 4867 4867
rect 4753 4833 4767 4847
rect 4713 4713 4727 4727
rect 4633 4334 4647 4348
rect 4713 4512 4727 4526
rect 4573 4292 4587 4306
rect 4613 4292 4627 4306
rect 4653 4292 4667 4306
rect 4553 4273 4567 4287
rect 4533 4253 4547 4267
rect 4573 4193 4587 4207
rect 4673 4173 4687 4187
rect 4513 4153 4527 4167
rect 4773 4812 4787 4826
rect 4813 4812 4827 4826
rect 4833 4593 4847 4607
rect 5033 5133 5047 5147
rect 5133 5133 5147 5147
rect 5253 5374 5267 5388
rect 5293 5374 5307 5388
rect 5233 5253 5247 5267
rect 5093 5093 5107 5107
rect 5193 5094 5207 5108
rect 5313 5332 5327 5346
rect 5593 5313 5607 5327
rect 5553 5273 5567 5287
rect 5373 5253 5387 5267
rect 5373 5213 5387 5227
rect 5353 5193 5367 5207
rect 5253 5153 5267 5167
rect 5393 5133 5407 5147
rect 5293 5113 5307 5127
rect 5053 5012 5067 5026
rect 5073 4973 5087 4987
rect 5013 4933 5027 4947
rect 4953 4854 4967 4868
rect 5013 4873 5027 4887
rect 5193 5073 5207 5087
rect 5253 5053 5267 5067
rect 5133 5032 5147 5046
rect 5173 5013 5187 5027
rect 5253 4993 5267 5007
rect 5133 4973 5147 4987
rect 5113 4873 5127 4887
rect 5073 4812 5087 4826
rect 5033 4753 5047 4767
rect 5053 4653 5067 4667
rect 4953 4593 4967 4607
rect 4933 4554 4947 4568
rect 4853 4513 4867 4527
rect 4913 4512 4927 4526
rect 4893 4473 4907 4487
rect 4873 4393 4887 4407
rect 4833 4354 4847 4368
rect 4793 4333 4807 4347
rect 4833 4333 4847 4347
rect 4933 4453 4947 4467
rect 4913 4353 4927 4367
rect 4753 4273 4767 4287
rect 4713 4213 4727 4227
rect 4613 4133 4627 4147
rect 4693 4133 4707 4147
rect 4553 4093 4567 4107
rect 4593 4093 4607 4107
rect 4473 4053 4487 4067
rect 4493 4034 4507 4048
rect 4513 3992 4527 4006
rect 4573 3992 4587 4006
rect 4473 3913 4487 3927
rect 4493 3893 4507 3907
rect 4473 3873 4487 3887
rect 4533 3814 4547 3828
rect 4493 3772 4507 3786
rect 4273 3693 4287 3707
rect 4433 3693 4447 3707
rect 4473 3693 4487 3707
rect 4093 3333 4107 3347
rect 4093 3294 4107 3308
rect 4113 3252 4127 3266
rect 4213 3294 4227 3308
rect 4173 3233 4187 3247
rect 4053 3133 4067 3147
rect 4093 3133 4107 3147
rect 4033 3113 4047 3127
rect 4033 3073 4047 3087
rect 4033 3052 4047 3066
rect 4073 3053 4087 3067
rect 4033 3013 4047 3027
rect 4073 3013 4087 3027
rect 4053 2994 4067 3008
rect 4133 3052 4147 3066
rect 4113 2993 4127 3007
rect 4033 2952 4047 2966
rect 4013 2853 4027 2867
rect 3993 2793 4007 2807
rect 4053 2793 4067 2807
rect 3933 2774 3947 2788
rect 3973 2774 3987 2788
rect 4033 2753 4047 2767
rect 3913 2733 3927 2747
rect 3893 2393 3907 2407
rect 3893 2293 3907 2307
rect 3893 2013 3907 2027
rect 3813 1954 3827 1968
rect 3873 1954 3887 1968
rect 3933 2474 3947 2488
rect 3913 1953 3927 1967
rect 3693 1933 3707 1947
rect 3733 1813 3747 1827
rect 3673 1773 3687 1787
rect 3773 1753 3787 1767
rect 3753 1734 3767 1748
rect 3653 1653 3667 1667
rect 3653 1613 3667 1627
rect 3673 1593 3687 1607
rect 3653 1573 3667 1587
rect 3833 1912 3847 1926
rect 3913 1912 3927 1926
rect 3892 1873 3906 1887
rect 3913 1873 3927 1887
rect 3893 1793 3907 1807
rect 4013 2474 4027 2488
rect 4093 2933 4107 2947
rect 4073 2733 4087 2747
rect 4073 2513 4087 2527
rect 4113 2913 4127 2927
rect 4113 2774 4127 2788
rect 4093 2473 4107 2487
rect 3993 2432 4007 2446
rect 3973 2393 3987 2407
rect 4013 2393 4027 2407
rect 3993 2353 4007 2367
rect 3973 2333 3987 2347
rect 3953 2173 3967 2187
rect 4073 2432 4087 2446
rect 4072 2353 4086 2367
rect 4093 2353 4107 2367
rect 4033 2313 4047 2327
rect 4093 2212 4107 2226
rect 3993 2133 4007 2147
rect 4053 2133 4067 2147
rect 3973 2093 3987 2107
rect 4093 2113 4107 2127
rect 4033 2073 4047 2087
rect 3993 1954 4007 1968
rect 4013 1912 4027 1926
rect 3993 1873 4007 1887
rect 3933 1753 3947 1767
rect 3813 1734 3827 1748
rect 3773 1573 3787 1587
rect 3713 1553 3727 1567
rect 3673 1533 3687 1547
rect 3772 1533 3786 1547
rect 3793 1533 3807 1547
rect 3773 1453 3787 1467
rect 3733 1434 3747 1448
rect 3753 1393 3767 1407
rect 3693 1353 3707 1367
rect 3633 1333 3647 1347
rect 3673 1293 3687 1307
rect 3493 1213 3507 1227
rect 3553 1214 3567 1228
rect 3593 1214 3607 1228
rect 3473 1172 3487 1186
rect 3453 1113 3467 1127
rect 3533 1172 3547 1186
rect 3573 1172 3587 1186
rect 3613 1172 3627 1186
rect 3493 1033 3507 1047
rect 3613 1033 3627 1047
rect 3393 914 3407 928
rect 3453 913 3467 927
rect 3533 932 3547 946
rect 3573 914 3587 928
rect 3233 733 3247 747
rect 3173 673 3187 687
rect 3253 652 3267 666
rect 3213 573 3227 587
rect 3193 393 3207 407
rect 3373 873 3387 887
rect 3453 872 3467 886
rect 3513 872 3527 886
rect 3433 713 3447 727
rect 3473 694 3487 708
rect 3453 652 3467 666
rect 3513 652 3527 666
rect 3653 1214 3667 1228
rect 3653 1173 3667 1187
rect 3693 1253 3707 1267
rect 3893 1733 3907 1747
rect 3953 1734 3967 1748
rect 3873 1633 3887 1647
rect 3833 1553 3847 1567
rect 3813 1453 3827 1467
rect 3873 1513 3887 1527
rect 3853 1433 3867 1447
rect 3933 1692 3947 1706
rect 3913 1633 3927 1647
rect 3933 1613 3947 1627
rect 3972 1573 3986 1587
rect 3993 1573 4007 1587
rect 3953 1493 3967 1507
rect 4073 1533 4087 1547
rect 4173 2993 4187 3007
rect 4173 2933 4187 2947
rect 4153 2853 4167 2867
rect 4173 2833 4187 2847
rect 4253 3333 4267 3347
rect 4253 3213 4267 3227
rect 4533 3653 4547 3667
rect 4473 3613 4487 3627
rect 4473 3553 4487 3567
rect 4293 3514 4307 3528
rect 4373 3514 4387 3528
rect 4433 3514 4447 3528
rect 4333 3453 4347 3467
rect 4453 3472 4467 3486
rect 4413 3453 4427 3467
rect 4373 3433 4387 3447
rect 4433 3433 4447 3447
rect 4333 3393 4347 3407
rect 4293 3333 4307 3347
rect 4353 3373 4367 3387
rect 4333 3313 4347 3327
rect 4313 3294 4327 3308
rect 4413 3333 4427 3347
rect 4393 3313 4407 3327
rect 4453 3353 4467 3367
rect 4433 3313 4447 3327
rect 4413 3213 4427 3227
rect 4393 3133 4407 3147
rect 4313 2994 4327 3008
rect 4333 2973 4347 2987
rect 4233 2933 4247 2947
rect 4273 2933 4287 2947
rect 4313 2933 4327 2947
rect 4213 2893 4227 2907
rect 4193 2813 4207 2827
rect 4253 2793 4267 2807
rect 4213 2774 4227 2788
rect 4173 1954 4187 1968
rect 4213 2693 4227 2707
rect 4213 2633 4227 2647
rect 4293 2813 4307 2827
rect 4293 2732 4307 2746
rect 4273 2673 4287 2687
rect 4393 2952 4407 2966
rect 4353 2933 4367 2947
rect 4433 3013 4447 3027
rect 4433 2913 4447 2927
rect 4393 2853 4407 2867
rect 4333 2773 4347 2787
rect 4433 2813 4447 2827
rect 4432 2774 4446 2788
rect 4593 3933 4607 3947
rect 4552 3513 4566 3527
rect 4573 3513 4587 3527
rect 4533 3472 4547 3486
rect 4533 3393 4547 3407
rect 4573 3333 4587 3347
rect 4853 4292 4867 4306
rect 4693 4034 4707 4048
rect 4733 4034 4747 4048
rect 4793 4034 4807 4048
rect 4653 4013 4667 4027
rect 4693 3973 4707 3987
rect 4653 3773 4667 3787
rect 4613 3513 4627 3527
rect 4653 3514 4667 3528
rect 4633 3472 4647 3486
rect 4612 3333 4626 3347
rect 4633 3333 4647 3347
rect 4553 3294 4567 3308
rect 4513 3273 4527 3287
rect 4513 3193 4527 3207
rect 4513 3113 4527 3127
rect 4493 3013 4507 3027
rect 4573 3213 4587 3227
rect 4553 3053 4567 3067
rect 4553 3013 4567 3027
rect 4493 2952 4507 2966
rect 4453 2773 4467 2787
rect 4373 2732 4387 2746
rect 4313 2653 4327 2667
rect 4253 2593 4267 2607
rect 4213 2573 4227 2587
rect 4313 2613 4327 2627
rect 4353 2613 4367 2627
rect 4313 2573 4327 2587
rect 4213 2533 4227 2547
rect 4273 2533 4287 2547
rect 4453 2733 4467 2747
rect 4253 2513 4267 2527
rect 4293 2513 4307 2527
rect 4413 2513 4427 2527
rect 4213 2474 4227 2488
rect 4253 2474 4267 2488
rect 4353 2473 4367 2487
rect 4293 2413 4307 2427
rect 4273 2353 4287 2367
rect 4333 2353 4347 2367
rect 4253 2333 4267 2347
rect 4293 2333 4307 2347
rect 4213 2313 4227 2327
rect 4253 2293 4267 2307
rect 4253 2254 4267 2268
rect 4273 2212 4287 2226
rect 4233 2173 4247 2187
rect 4373 2393 4387 2407
rect 4353 2212 4367 2226
rect 4353 2173 4367 2187
rect 4233 2013 4247 2027
rect 4273 1954 4287 1968
rect 4173 1913 4187 1927
rect 4213 1873 4227 1887
rect 4173 1813 4187 1827
rect 4333 1813 4347 1827
rect 4213 1734 4227 1748
rect 4253 1734 4267 1748
rect 4193 1593 4207 1607
rect 4153 1573 4167 1587
rect 4153 1533 4167 1547
rect 4133 1473 4147 1487
rect 4253 1473 4267 1487
rect 4013 1453 4027 1467
rect 4213 1453 4227 1467
rect 3833 1293 3847 1307
rect 3993 1433 4007 1447
rect 3873 1392 3887 1406
rect 3933 1392 3947 1406
rect 3973 1392 3987 1406
rect 3873 1333 3887 1347
rect 3853 1253 3867 1267
rect 3753 1213 3767 1227
rect 3793 1213 3807 1227
rect 3893 1253 3907 1267
rect 3873 1213 3887 1227
rect 3773 1172 3787 1186
rect 3853 1172 3867 1186
rect 3873 1133 3887 1147
rect 3813 1113 3827 1127
rect 3693 1053 3707 1067
rect 3673 933 3687 947
rect 3773 1033 3787 1047
rect 3733 914 3747 928
rect 3873 1053 3887 1067
rect 3813 993 3827 1007
rect 3833 953 3847 967
rect 3693 872 3707 886
rect 3753 872 3767 886
rect 3793 872 3807 886
rect 3633 773 3647 787
rect 3673 694 3687 708
rect 3653 652 3667 666
rect 3613 593 3627 607
rect 3693 593 3707 607
rect 3913 1193 3927 1207
rect 3913 1153 3927 1167
rect 4093 1433 4107 1447
rect 4153 1434 4167 1448
rect 4013 1353 4027 1367
rect 4053 1214 4067 1228
rect 4173 1392 4187 1406
rect 4133 1313 4147 1327
rect 4133 1213 4147 1227
rect 3953 1153 3967 1167
rect 4073 1172 4087 1186
rect 4113 1172 4127 1186
rect 4053 1133 4067 1147
rect 4033 1113 4047 1127
rect 3933 1093 3947 1107
rect 3993 914 4007 928
rect 3953 873 3967 887
rect 4013 872 4027 886
rect 4053 872 4067 886
rect 3893 833 3907 847
rect 4233 1313 4247 1327
rect 4273 1293 4287 1307
rect 4253 1253 4267 1267
rect 4413 2313 4427 2327
rect 4493 2773 4507 2787
rect 4473 2473 4487 2487
rect 4553 2733 4567 2747
rect 4533 2673 4547 2687
rect 4633 3173 4647 3187
rect 4673 3353 4687 3367
rect 4753 3992 4767 4006
rect 4793 3973 4807 3987
rect 4713 3933 4727 3947
rect 4813 3933 4827 3947
rect 4853 4213 4867 4227
rect 4733 3913 4747 3927
rect 4833 3913 4847 3927
rect 4713 3814 4727 3828
rect 4773 3853 4787 3867
rect 4753 3733 4767 3747
rect 4873 4173 4887 4187
rect 4873 4034 4887 4048
rect 4973 4393 4987 4407
rect 5273 4933 5287 4947
rect 5573 5013 5587 5027
rect 5533 4953 5547 4967
rect 5533 4932 5547 4946
rect 5293 4913 5307 4927
rect 5413 4913 5427 4927
rect 5192 4893 5206 4907
rect 5213 4893 5227 4907
rect 5333 4893 5347 4907
rect 5173 4873 5187 4887
rect 5133 4633 5147 4647
rect 5113 4593 5127 4607
rect 5113 4554 5127 4568
rect 5093 4453 5107 4467
rect 5153 4334 5167 4348
rect 5013 4292 5027 4306
rect 5113 4292 5127 4306
rect 4973 4252 4987 4266
rect 5053 4253 5067 4267
rect 4933 4133 4947 4147
rect 4933 4034 4947 4048
rect 5093 4233 5107 4247
rect 5153 4233 5167 4247
rect 5053 4153 5067 4167
rect 5013 4034 5027 4048
rect 4893 3992 4907 4006
rect 4953 3992 4967 4006
rect 4933 3973 4947 3987
rect 4913 3953 4927 3967
rect 4913 3913 4927 3927
rect 4913 3813 4927 3827
rect 4853 3733 4867 3747
rect 4892 3693 4906 3707
rect 4913 3693 4927 3707
rect 4853 3633 4867 3647
rect 4793 3593 4807 3607
rect 4713 3573 4727 3587
rect 4833 3573 4847 3587
rect 4693 3293 4707 3307
rect 4673 3073 4687 3087
rect 4753 3553 4767 3567
rect 4733 3513 4747 3527
rect 4733 3472 4747 3486
rect 4893 3514 4907 3528
rect 4833 3472 4847 3486
rect 4873 3472 4887 3486
rect 4773 3453 4787 3467
rect 4893 3453 4907 3467
rect 4853 3393 4867 3407
rect 4833 3353 4847 3367
rect 4713 3252 4727 3266
rect 4793 3294 4807 3308
rect 4853 3294 4867 3308
rect 4773 3252 4787 3266
rect 4733 3213 4747 3227
rect 4813 3213 4827 3227
rect 4813 3173 4827 3187
rect 4713 3153 4727 3167
rect 4693 3013 4707 3027
rect 4773 3013 4787 3027
rect 4653 2893 4667 2907
rect 4753 2893 4767 2907
rect 4733 2853 4747 2867
rect 4693 2833 4707 2847
rect 4633 2774 4647 2788
rect 4553 2432 4567 2446
rect 4593 2432 4607 2446
rect 4513 2373 4527 2387
rect 4533 2353 4547 2367
rect 4453 2293 4467 2307
rect 4433 2253 4447 2267
rect 4493 2254 4507 2268
rect 4433 2212 4447 2226
rect 4473 2212 4487 2226
rect 4513 2212 4527 2226
rect 4473 2153 4487 2167
rect 4413 2093 4427 2107
rect 4373 2073 4387 2087
rect 4433 1993 4447 2007
rect 4533 2073 4547 2087
rect 4433 1853 4447 1867
rect 4393 1734 4407 1748
rect 4473 1893 4487 1907
rect 4493 1873 4507 1887
rect 4533 1873 4547 1887
rect 4473 1833 4487 1847
rect 4453 1813 4467 1827
rect 4513 1813 4527 1827
rect 4473 1773 4487 1787
rect 4393 1373 4407 1387
rect 4333 1193 4347 1207
rect 4393 1213 4407 1227
rect 4353 1033 4367 1047
rect 4213 953 4227 967
rect 4253 953 4267 967
rect 4153 913 4167 927
rect 4153 833 4167 847
rect 4133 773 4147 787
rect 3873 733 3887 747
rect 4113 733 4127 747
rect 3913 694 3927 708
rect 4153 694 4167 708
rect 3893 633 3907 647
rect 4093 613 4107 627
rect 4133 613 4147 627
rect 3833 533 3847 547
rect 3613 473 3627 487
rect 3953 473 3967 487
rect 3573 453 3587 467
rect 3353 433 3367 447
rect 3553 433 3567 447
rect 3553 412 3567 426
rect 3113 352 3127 366
rect 2913 133 2927 147
rect 3233 353 3247 367
rect 3253 333 3267 347
rect 3253 293 3267 307
rect 3253 272 3267 286
rect 3293 313 3307 327
rect 4233 833 4247 847
rect 4213 693 4227 707
rect 4093 433 4107 447
rect 4193 433 4207 447
rect 3693 413 3707 427
rect 3653 394 3667 408
rect 3953 413 3967 427
rect 3733 373 3747 387
rect 3573 352 3587 366
rect 3613 352 3627 366
rect 3933 352 3947 366
rect 3673 313 3687 327
rect 3733 313 3747 327
rect 3753 293 3767 307
rect 3373 273 3387 287
rect 3553 273 3567 287
rect 3293 233 3307 247
rect 3753 233 3767 247
rect 3953 233 3967 247
rect 3273 213 3287 227
rect 3313 174 3327 188
rect 3473 174 3487 188
rect 3513 174 3527 188
rect 3033 132 3047 146
rect 3193 132 3207 146
rect 3233 132 3247 146
rect 3553 173 3567 187
rect 3693 174 3707 188
rect 3733 174 3747 188
rect 3793 174 3807 188
rect 4153 394 4167 408
rect 4133 352 4147 366
rect 4373 913 4387 927
rect 4313 833 4327 847
rect 4453 1693 4467 1707
rect 4433 1393 4447 1407
rect 4433 1313 4447 1327
rect 4473 1513 4487 1527
rect 4453 1213 4467 1227
rect 4593 1833 4607 1847
rect 4673 2473 4687 2487
rect 4673 2353 4687 2367
rect 4813 2873 4827 2887
rect 4813 2852 4827 2866
rect 4773 2833 4787 2847
rect 4753 2732 4767 2746
rect 4713 2713 4727 2727
rect 4713 2593 4727 2607
rect 4913 3373 4927 3387
rect 4953 3953 4967 3967
rect 5033 3933 5047 3947
rect 4993 3893 5007 3907
rect 4993 3814 5007 3828
rect 5073 4133 5087 4147
rect 5053 3813 5067 3827
rect 4953 3773 4967 3787
rect 4953 3653 4967 3667
rect 4953 3514 4967 3528
rect 5013 3772 5027 3786
rect 4993 3733 5007 3747
rect 4973 3453 4987 3467
rect 4953 3393 4967 3407
rect 5073 3613 5087 3627
rect 5173 4213 5187 4227
rect 5353 4872 5367 4886
rect 5253 4854 5267 4868
rect 5293 4854 5307 4868
rect 5213 4812 5227 4826
rect 5313 4812 5327 4826
rect 5233 4713 5247 4727
rect 5233 4433 5247 4447
rect 5333 4753 5347 4767
rect 5293 4573 5307 4587
rect 5373 4853 5387 4867
rect 5373 4773 5387 4787
rect 5353 4653 5367 4667
rect 5373 4613 5387 4627
rect 5313 4512 5327 4526
rect 5293 4413 5307 4427
rect 5353 4413 5367 4427
rect 5313 4353 5327 4367
rect 5353 4353 5367 4367
rect 5373 4313 5387 4327
rect 5313 4292 5327 4306
rect 5353 4293 5367 4307
rect 5253 4253 5267 4267
rect 5313 4213 5327 4227
rect 5193 4153 5207 4167
rect 5293 4133 5307 4147
rect 5253 4073 5267 4087
rect 5113 4034 5127 4048
rect 5153 4034 5167 4048
rect 5213 4034 5227 4048
rect 5113 3993 5127 4007
rect 5153 3893 5167 3907
rect 5113 3813 5127 3827
rect 5093 3553 5107 3567
rect 5013 3514 5027 3528
rect 5013 3473 5027 3487
rect 5073 3514 5087 3528
rect 5153 3673 5167 3687
rect 5093 3472 5107 3486
rect 5033 3413 5047 3427
rect 5153 3413 5167 3427
rect 4993 3353 5007 3367
rect 5113 3353 5127 3367
rect 5093 3333 5107 3347
rect 5053 3313 5067 3327
rect 4953 3293 4967 3307
rect 5013 3294 5027 3308
rect 5053 3294 5067 3308
rect 4933 3273 4947 3287
rect 4913 3193 4927 3207
rect 4893 3173 4907 3187
rect 5093 3253 5107 3267
rect 5033 3233 5047 3247
rect 4953 3173 4967 3187
rect 5013 3173 5027 3187
rect 4893 3073 4907 3087
rect 4933 3073 4947 3087
rect 4893 2994 4907 3008
rect 4933 2994 4947 3008
rect 4913 2952 4927 2966
rect 4873 2933 4887 2947
rect 4853 2893 4867 2907
rect 4833 2813 4847 2827
rect 4793 2773 4807 2787
rect 4872 2853 4886 2867
rect 4893 2853 4907 2867
rect 4853 2793 4867 2807
rect 4913 2774 4927 2788
rect 5013 2952 5027 2966
rect 4973 2933 4987 2947
rect 4853 2732 4867 2746
rect 4793 2693 4807 2707
rect 4813 2673 4827 2687
rect 4793 2633 4807 2647
rect 4773 2493 4787 2507
rect 4753 2474 4767 2488
rect 4953 2732 4967 2746
rect 4913 2693 4927 2707
rect 4893 2673 4907 2687
rect 4833 2653 4847 2667
rect 4813 2432 4827 2446
rect 4733 2333 4747 2347
rect 4753 2313 4767 2327
rect 4713 2254 4727 2268
rect 4792 2254 4806 2268
rect 4813 2253 4827 2267
rect 4673 2212 4687 2226
rect 4653 2133 4667 2147
rect 4633 2033 4647 2047
rect 4673 1993 4687 2007
rect 4713 1993 4727 2007
rect 4793 2213 4807 2227
rect 4773 2193 4787 2207
rect 4813 2153 4827 2167
rect 4773 2033 4787 2047
rect 4793 1954 4807 1968
rect 4693 1912 4707 1926
rect 4793 1913 4807 1927
rect 4613 1813 4627 1827
rect 4533 1753 4547 1767
rect 4573 1753 4587 1767
rect 4553 1713 4567 1727
rect 4993 2653 5007 2667
rect 5013 2593 5027 2607
rect 4993 2533 5007 2547
rect 4893 2513 4907 2527
rect 4973 2513 4987 2527
rect 4853 2493 4867 2507
rect 4833 1913 4847 1927
rect 4813 1733 4827 1747
rect 5013 2493 5027 2507
rect 4953 2474 4967 2488
rect 4933 2432 4947 2446
rect 4973 2432 4987 2446
rect 5013 2432 5027 2446
rect 4912 2373 4926 2387
rect 4933 2372 4947 2386
rect 4873 2333 4887 2347
rect 4913 2333 4927 2347
rect 5133 3333 5147 3347
rect 5153 3233 5167 3247
rect 5133 3133 5147 3147
rect 5153 3113 5167 3127
rect 5233 3992 5247 4006
rect 5293 3993 5307 4007
rect 5193 3933 5207 3947
rect 5213 3913 5227 3927
rect 5213 3873 5227 3887
rect 5253 3873 5267 3887
rect 5573 4913 5587 4927
rect 5673 5614 5687 5628
rect 5633 5572 5647 5586
rect 5653 5553 5667 5567
rect 5633 5453 5647 5467
rect 5833 7513 5847 7527
rect 5913 7513 5927 7527
rect 5873 7454 5887 7468
rect 5813 7413 5827 7427
rect 5793 7092 5807 7106
rect 5813 7073 5827 7087
rect 5913 7393 5927 7407
rect 5853 7373 5867 7387
rect 5973 8073 5987 8087
rect 5973 7913 5987 7927
rect 5953 7893 5967 7907
rect 5933 7333 5947 7347
rect 5973 7673 5987 7687
rect 5973 7533 5987 7547
rect 5973 7493 5987 7507
rect 5973 7454 5987 7468
rect 5973 7293 5987 7307
rect 5953 7173 5967 7187
rect 5873 7154 5887 7168
rect 5913 7154 5927 7168
rect 5933 7112 5947 7126
rect 5872 7073 5886 7087
rect 5893 7073 5907 7087
rect 5793 6933 5807 6947
rect 5833 6933 5847 6947
rect 5813 6892 5827 6906
rect 5893 6953 5907 6967
rect 5873 6833 5887 6847
rect 5893 6753 5907 6767
rect 5913 6733 5927 6747
rect 5893 6713 5907 6727
rect 5793 6673 5807 6687
rect 5833 6673 5847 6687
rect 6053 8194 6067 8208
rect 6053 8113 6067 8127
rect 6033 8093 6047 8107
rect 6073 8073 6087 8087
rect 6033 7993 6047 8007
rect 6193 8393 6207 8407
rect 6113 8313 6127 8327
rect 6093 8013 6107 8027
rect 6273 8273 6287 8287
rect 6173 8233 6187 8247
rect 6253 8233 6267 8247
rect 6253 8212 6267 8226
rect 6153 8113 6167 8127
rect 6053 7913 6067 7927
rect 6113 7913 6127 7927
rect 6093 7893 6107 7907
rect 6073 7833 6087 7847
rect 6093 7773 6107 7787
rect 6073 7693 6087 7707
rect 6013 7674 6027 7688
rect 6013 7613 6027 7627
rect 6093 7593 6107 7607
rect 6133 7693 6147 7707
rect 6052 7393 6066 7407
rect 6073 7393 6087 7407
rect 6113 7393 6127 7407
rect 6053 7353 6067 7367
rect 6053 7233 6067 7247
rect 6033 7213 6047 7227
rect 6013 7113 6027 7127
rect 5993 7073 6007 7087
rect 6173 8093 6187 8107
rect 6173 8033 6187 8047
rect 6173 8012 6187 8026
rect 6273 8113 6287 8127
rect 6233 8053 6247 8067
rect 6193 7933 6207 7947
rect 6173 7813 6187 7827
rect 6213 7753 6227 7767
rect 6173 7733 6187 7747
rect 6333 8733 6347 8747
rect 6333 8672 6347 8686
rect 6373 9333 6387 9347
rect 6533 10313 6547 10327
rect 6533 10274 6547 10288
rect 6633 10473 6647 10487
rect 6633 10433 6647 10447
rect 6793 10553 6807 10567
rect 6713 10532 6727 10546
rect 7133 11094 7147 11108
rect 7193 11093 7207 11107
rect 7293 11094 7307 11108
rect 7333 11094 7347 11108
rect 7473 11094 7487 11108
rect 7593 11094 7607 11108
rect 7993 11113 8007 11127
rect 8273 11113 8287 11127
rect 7853 11094 7867 11108
rect 7073 11033 7087 11047
rect 7153 11052 7167 11066
rect 7113 11013 7127 11027
rect 7153 11013 7167 11027
rect 7033 10973 7047 10987
rect 6913 10813 6927 10827
rect 6933 10793 6947 10807
rect 6993 10794 7007 10808
rect 7113 10933 7127 10947
rect 7113 10794 7127 10808
rect 7013 10752 7027 10766
rect 6933 10733 6947 10747
rect 7053 10733 7067 10747
rect 6993 10693 7007 10707
rect 6893 10574 6907 10588
rect 6953 10574 6967 10588
rect 6733 10473 6747 10487
rect 6553 10232 6567 10246
rect 6593 10232 6607 10246
rect 6693 10274 6707 10288
rect 6693 10233 6707 10247
rect 6813 10393 6827 10407
rect 6773 10274 6787 10288
rect 7053 10573 7067 10587
rect 7133 10673 7147 10687
rect 6893 10473 6907 10487
rect 7013 10532 7027 10546
rect 7113 10533 7127 10547
rect 6973 10513 6987 10527
rect 6933 10453 6947 10467
rect 6853 10373 6867 10387
rect 6973 10373 6987 10387
rect 6933 10333 6947 10347
rect 6853 10313 6867 10327
rect 6893 10274 6907 10288
rect 6733 10213 6747 10227
rect 6793 10213 6807 10227
rect 6753 10193 6767 10207
rect 6633 10173 6647 10187
rect 6713 10133 6727 10147
rect 6493 10113 6507 10127
rect 6633 10113 6647 10127
rect 6473 10054 6487 10068
rect 6473 9793 6487 9807
rect 6553 10054 6567 10068
rect 6593 10054 6607 10068
rect 6673 10054 6687 10068
rect 6553 9973 6567 9987
rect 6653 9993 6667 10007
rect 6613 9933 6627 9947
rect 6533 9873 6547 9887
rect 6493 9753 6507 9767
rect 6613 9853 6627 9867
rect 6573 9793 6587 9807
rect 6693 9793 6707 9807
rect 6613 9754 6627 9768
rect 6473 9534 6487 9548
rect 6513 9534 6527 9548
rect 6533 9492 6547 9506
rect 6473 9473 6487 9487
rect 6553 9433 6567 9447
rect 6453 9413 6467 9427
rect 6513 9293 6527 9307
rect 6473 9234 6487 9248
rect 6453 9192 6467 9206
rect 6413 9153 6427 9167
rect 6373 9093 6387 9107
rect 6393 9053 6407 9067
rect 6373 8893 6387 8907
rect 6393 8873 6407 8887
rect 6613 9693 6627 9707
rect 6593 9633 6607 9647
rect 6593 9593 6607 9607
rect 6593 9534 6607 9548
rect 6593 9493 6607 9507
rect 6593 9413 6607 9427
rect 6573 9293 6587 9307
rect 6553 9273 6567 9287
rect 6473 9073 6487 9087
rect 6513 9073 6527 9087
rect 6473 8972 6487 8986
rect 6513 8913 6527 8927
rect 6373 8633 6387 8647
rect 6353 8553 6367 8567
rect 6333 8313 6347 8327
rect 6493 8833 6507 8847
rect 6453 8714 6467 8728
rect 6573 8733 6587 8747
rect 6433 8672 6447 8686
rect 6453 8653 6467 8667
rect 6413 8593 6427 8607
rect 6393 8573 6407 8587
rect 6373 8353 6387 8367
rect 6353 8273 6367 8287
rect 6333 8213 6347 8227
rect 6293 7974 6307 7988
rect 6513 8672 6527 8686
rect 6513 8633 6527 8647
rect 6473 8533 6487 8547
rect 6433 8493 6447 8507
rect 6473 8494 6487 8508
rect 6733 10053 6747 10067
rect 6733 9773 6747 9787
rect 6713 9693 6727 9707
rect 6693 9573 6707 9587
rect 6693 9534 6707 9548
rect 6833 10193 6847 10207
rect 6813 10173 6827 10187
rect 6933 10193 6947 10207
rect 7133 10413 7147 10427
rect 7053 10373 7067 10387
rect 7113 10373 7127 10387
rect 7013 10333 7027 10347
rect 7013 10274 7027 10288
rect 7113 10313 7127 10327
rect 7033 10213 7047 10227
rect 6913 10054 6927 10068
rect 6973 10052 6987 10066
rect 6853 10012 6867 10026
rect 6973 10013 6987 10027
rect 7053 9993 7067 10007
rect 6813 9953 6827 9967
rect 6853 9953 6867 9967
rect 6793 9853 6807 9867
rect 6813 9754 6827 9768
rect 6753 9713 6767 9727
rect 6793 9712 6807 9726
rect 6793 9633 6807 9647
rect 6713 9492 6727 9506
rect 6673 9373 6687 9387
rect 6713 9333 6727 9347
rect 6613 9193 6627 9207
rect 6693 9192 6707 9206
rect 6653 9153 6667 9167
rect 6753 9153 6767 9167
rect 6613 9014 6627 9028
rect 6833 9493 6847 9507
rect 6833 9234 6847 9248
rect 6873 9933 6887 9947
rect 6913 9754 6927 9768
rect 6953 9754 6967 9768
rect 7013 9754 7027 9768
rect 6873 9733 6887 9747
rect 6873 9712 6887 9726
rect 6993 9712 7007 9726
rect 7033 9712 7047 9726
rect 6913 9673 6927 9687
rect 6993 9673 7007 9687
rect 6933 9534 6947 9548
rect 6873 9513 6887 9527
rect 6913 9492 6927 9506
rect 6953 9393 6967 9407
rect 7053 9533 7067 9547
rect 7053 9492 7067 9506
rect 6993 9353 7007 9367
rect 6913 9313 6927 9327
rect 6953 9234 6967 9248
rect 7133 9653 7147 9667
rect 7173 10933 7187 10947
rect 7353 11052 7367 11066
rect 7393 11033 7407 11047
rect 7293 11013 7307 11027
rect 7433 10993 7447 11007
rect 7293 10833 7307 10847
rect 7333 10833 7347 10847
rect 7253 10794 7267 10808
rect 7373 10813 7387 10827
rect 7173 10753 7187 10767
rect 7353 10752 7367 10766
rect 7313 10733 7327 10747
rect 7273 10633 7287 10647
rect 7193 10613 7207 10627
rect 7233 10613 7247 10627
rect 7253 10532 7267 10546
rect 7353 10533 7367 10547
rect 7213 10513 7227 10527
rect 7333 10493 7347 10507
rect 7253 10393 7267 10407
rect 7313 10313 7327 10327
rect 7292 10274 7306 10288
rect 7313 10273 7327 10287
rect 7913 11093 7927 11107
rect 7933 11073 7947 11087
rect 7573 11052 7587 11066
rect 7513 11033 7527 11047
rect 7473 10933 7487 10947
rect 7473 10873 7487 10887
rect 7493 10833 7507 10847
rect 7553 10833 7567 10847
rect 7513 10813 7527 10827
rect 7433 10753 7447 10767
rect 7573 10813 7587 10827
rect 7593 10794 7607 10808
rect 7513 10752 7527 10766
rect 7553 10752 7567 10766
rect 7453 10653 7467 10667
rect 7493 10653 7507 10667
rect 7593 10573 7607 10587
rect 7393 10533 7407 10547
rect 7373 10313 7387 10327
rect 7233 10213 7247 10227
rect 7273 10213 7287 10227
rect 7173 10054 7187 10068
rect 7453 10532 7467 10546
rect 7493 10533 7507 10547
rect 7533 10433 7547 10447
rect 7433 10413 7447 10427
rect 7413 10293 7427 10307
rect 7393 10133 7407 10147
rect 7293 10012 7307 10026
rect 7193 9993 7207 10007
rect 7153 9633 7167 9647
rect 7173 9573 7187 9587
rect 7533 10353 7547 10367
rect 7553 10333 7567 10347
rect 7513 10313 7527 10327
rect 7473 10293 7487 10307
rect 7493 10232 7507 10246
rect 7433 10213 7447 10227
rect 7513 10193 7527 10207
rect 7553 10054 7567 10068
rect 7533 10012 7547 10026
rect 7493 9993 7507 10007
rect 7413 9953 7427 9967
rect 7273 9873 7287 9887
rect 7313 9873 7327 9887
rect 7233 9813 7247 9827
rect 7873 11052 7887 11066
rect 7913 11052 7927 11066
rect 7833 10973 7847 10987
rect 7913 10953 7927 10967
rect 7773 10794 7787 10808
rect 7813 10794 7827 10808
rect 7893 10794 7907 10808
rect 7753 10752 7767 10766
rect 7793 10752 7807 10766
rect 7793 10713 7807 10727
rect 7653 10633 7667 10647
rect 7633 10532 7647 10546
rect 7613 10493 7627 10507
rect 7693 10493 7707 10507
rect 7653 10453 7667 10467
rect 7673 10393 7687 10407
rect 7653 10273 7667 10287
rect 7713 10274 7727 10288
rect 7753 10274 7767 10288
rect 7653 10233 7667 10247
rect 7613 10173 7627 10187
rect 7953 11052 7967 11066
rect 7933 10893 7947 10907
rect 7933 10793 7947 10807
rect 7913 10773 7927 10787
rect 7933 10573 7947 10587
rect 8073 11094 8087 11108
rect 8313 11094 8327 11108
rect 8513 11094 8527 11108
rect 8733 11094 8747 11108
rect 8873 11093 8887 11107
rect 9093 11113 9107 11127
rect 9173 11113 9187 11127
rect 8993 11094 9007 11108
rect 9033 11094 9047 11108
rect 8053 11052 8067 11066
rect 8093 10993 8107 11007
rect 8033 10913 8047 10927
rect 8293 10913 8307 10927
rect 7993 10794 8007 10808
rect 8213 10833 8227 10847
rect 8253 10833 8267 10847
rect 8153 10794 8167 10808
rect 8213 10794 8227 10808
rect 8253 10793 8267 10807
rect 8013 10752 8027 10766
rect 8153 10753 8167 10767
rect 8133 10713 8147 10727
rect 8093 10653 8107 10667
rect 8033 10633 8047 10647
rect 7873 10532 7887 10546
rect 7873 10373 7887 10387
rect 7853 10333 7867 10347
rect 7813 10274 7827 10288
rect 7853 10274 7867 10288
rect 7813 10233 7827 10247
rect 7733 10192 7747 10206
rect 7693 10153 7707 10167
rect 7673 10133 7687 10147
rect 7613 10012 7627 10026
rect 7653 10012 7667 10026
rect 7613 9913 7627 9927
rect 7593 9813 7607 9827
rect 7433 9773 7447 9787
rect 7473 9773 7487 9787
rect 7273 9754 7287 9768
rect 7333 9754 7347 9768
rect 7413 9754 7427 9768
rect 7293 9693 7307 9707
rect 7413 9693 7427 9707
rect 7253 9633 7267 9647
rect 7233 9533 7247 9547
rect 7113 9492 7127 9506
rect 7213 9492 7227 9506
rect 7213 9453 7227 9467
rect 7313 9613 7327 9627
rect 7173 9433 7187 9447
rect 7093 9234 7107 9248
rect 7133 9234 7147 9248
rect 7173 9234 7187 9248
rect 6853 9193 6867 9207
rect 6933 9192 6947 9206
rect 7093 9193 7107 9207
rect 7153 9192 7167 9206
rect 6893 9153 6907 9167
rect 6833 9113 6847 9127
rect 6813 8972 6827 8986
rect 6853 8913 6867 8927
rect 7013 8992 7027 9006
rect 7153 8994 7167 9008
rect 7193 8994 7207 9008
rect 7013 8913 7027 8927
rect 6773 8813 6787 8827
rect 7013 8813 7027 8827
rect 7053 8813 7067 8827
rect 6913 8773 6927 8787
rect 7033 8773 7047 8787
rect 6873 8733 6887 8747
rect 6693 8714 6707 8728
rect 6753 8713 6767 8727
rect 6953 8733 6967 8747
rect 6673 8672 6687 8686
rect 6753 8672 6767 8686
rect 6853 8672 6867 8686
rect 6613 8633 6627 8647
rect 6453 8452 6467 8466
rect 6493 8453 6507 8467
rect 6473 8373 6487 8387
rect 6393 8293 6407 8307
rect 6433 8113 6447 8127
rect 6313 7932 6327 7946
rect 6353 7793 6367 7807
rect 6313 7753 6327 7767
rect 6233 7693 6247 7707
rect 6253 7674 6267 7688
rect 6193 7573 6207 7587
rect 6173 7513 6187 7527
rect 6273 7633 6287 7647
rect 6213 7453 6227 7467
rect 6473 8053 6487 8067
rect 6513 8393 6527 8407
rect 6513 8073 6527 8087
rect 6493 8013 6507 8027
rect 6473 7993 6487 8007
rect 6453 7973 6467 7987
rect 6393 7853 6407 7867
rect 6393 7793 6407 7807
rect 6393 7772 6407 7786
rect 6373 7753 6387 7767
rect 6353 7713 6367 7727
rect 6352 7674 6366 7688
rect 6373 7674 6387 7688
rect 6313 7454 6327 7468
rect 6193 7313 6207 7327
rect 6153 7253 6167 7267
rect 6133 7233 6147 7247
rect 6193 7193 6207 7207
rect 6133 7173 6147 7187
rect 6073 7154 6087 7168
rect 6173 7154 6187 7168
rect 6373 7633 6387 7647
rect 6353 7433 6367 7447
rect 6293 7412 6307 7426
rect 6253 7373 6267 7387
rect 6573 8493 6587 8507
rect 6933 8653 6947 8667
rect 6753 8472 6767 8486
rect 6613 8393 6627 8407
rect 6893 8472 6907 8486
rect 6933 8473 6947 8487
rect 6913 8432 6927 8446
rect 6813 8293 6827 8307
rect 6933 8293 6947 8307
rect 6793 8253 6807 8267
rect 6633 8233 6647 8247
rect 6653 8194 6667 8208
rect 6713 8194 6727 8208
rect 6633 8152 6647 8166
rect 6673 8152 6687 8166
rect 6613 8133 6627 8147
rect 6593 8093 6607 8107
rect 6573 8013 6587 8027
rect 6553 7973 6567 7987
rect 6533 7913 6547 7927
rect 6473 7833 6487 7847
rect 6473 7812 6487 7826
rect 6453 7753 6467 7767
rect 6433 7733 6447 7747
rect 6533 7733 6547 7747
rect 6433 7674 6447 7688
rect 6473 7674 6487 7688
rect 6413 7633 6427 7647
rect 6253 7352 6267 7366
rect 6333 7353 6347 7367
rect 6393 7353 6407 7367
rect 6273 7333 6287 7347
rect 6253 7193 6267 7207
rect 6053 7133 6067 7147
rect 6093 7093 6107 7107
rect 6073 7033 6087 7047
rect 6053 7013 6067 7027
rect 6033 6993 6047 7007
rect 5973 6973 5987 6987
rect 6153 7093 6167 7107
rect 6073 6934 6087 6948
rect 6113 6934 6127 6948
rect 5973 6892 5987 6906
rect 6013 6892 6027 6906
rect 6053 6892 6067 6906
rect 6033 6833 6047 6847
rect 5953 6753 5967 6767
rect 5953 6713 5967 6727
rect 5933 6673 5947 6687
rect 5913 6653 5927 6667
rect 5873 6634 5887 6648
rect 5853 6592 5867 6606
rect 5893 6592 5907 6606
rect 5793 6513 5807 6527
rect 5853 6353 5867 6367
rect 5813 6333 5827 6347
rect 5773 6253 5787 6267
rect 5813 6213 5827 6227
rect 5813 6134 5827 6148
rect 5973 6673 5987 6687
rect 5953 6593 5967 6607
rect 5933 6473 5947 6487
rect 6013 6653 6027 6667
rect 5973 6453 5987 6467
rect 5893 6293 5907 6307
rect 5973 6333 5987 6347
rect 5873 6253 5887 6267
rect 5933 6253 5947 6267
rect 5793 6093 5807 6107
rect 5853 6093 5867 6107
rect 5773 6053 5787 6067
rect 5753 5973 5767 5987
rect 5853 6072 5867 6086
rect 5833 6013 5847 6027
rect 5833 5893 5847 5907
rect 5733 5813 5747 5827
rect 5733 5673 5747 5687
rect 5733 5553 5747 5567
rect 5713 5453 5727 5467
rect 5673 5374 5687 5388
rect 5713 5374 5727 5388
rect 5773 5852 5787 5866
rect 5833 5853 5847 5867
rect 5773 5653 5787 5667
rect 5813 5653 5827 5667
rect 5793 5614 5807 5628
rect 5813 5513 5827 5527
rect 5813 5473 5827 5487
rect 5813 5373 5827 5387
rect 5673 5332 5687 5346
rect 5653 5273 5667 5287
rect 5613 5113 5627 5127
rect 5613 5053 5627 5067
rect 5693 5253 5707 5267
rect 6153 6993 6167 7007
rect 6153 6813 6167 6827
rect 6133 6773 6147 6787
rect 6113 6713 6127 6727
rect 6133 6673 6147 6687
rect 6053 6633 6067 6647
rect 6093 6634 6107 6648
rect 6073 6592 6087 6606
rect 6113 6592 6127 6606
rect 6073 6553 6087 6567
rect 6033 6313 6047 6327
rect 6193 7073 6207 7087
rect 6253 7154 6267 7168
rect 6313 7253 6327 7267
rect 6293 7233 6307 7247
rect 6273 7073 6287 7087
rect 6293 7053 6307 7067
rect 6273 7013 6287 7027
rect 6293 6993 6307 7007
rect 6193 6673 6207 6687
rect 6173 6533 6187 6547
rect 6133 6433 6147 6447
rect 6173 6414 6187 6428
rect 6293 6953 6307 6967
rect 6273 6892 6287 6906
rect 6493 7632 6507 7646
rect 6533 7632 6547 7646
rect 6493 7573 6507 7587
rect 6513 7454 6527 7468
rect 6573 7853 6587 7867
rect 6593 7713 6607 7727
rect 6573 7533 6587 7547
rect 6593 7513 6607 7527
rect 6553 7453 6567 7467
rect 6673 8093 6687 8107
rect 6793 8173 6807 8187
rect 6853 8194 6867 8208
rect 6913 8173 6927 8187
rect 6833 8153 6847 8167
rect 6833 8093 6847 8107
rect 6873 8093 6887 8107
rect 6813 8073 6827 8087
rect 6973 8693 6987 8707
rect 6993 8672 7007 8686
rect 6973 8613 6987 8627
rect 6973 8533 6987 8547
rect 6953 8133 6967 8147
rect 6933 8113 6947 8127
rect 6713 8053 6727 8067
rect 6913 8053 6927 8067
rect 6673 7993 6687 8007
rect 6633 7973 6647 7987
rect 7033 8493 7047 8507
rect 7033 8472 7047 8486
rect 7293 9233 7307 9247
rect 7273 9173 7287 9187
rect 7513 9754 7527 9768
rect 7433 9573 7447 9587
rect 7373 9534 7387 9548
rect 7433 9533 7447 9547
rect 7533 9693 7547 9707
rect 7493 9673 7507 9687
rect 7593 9693 7607 9707
rect 7573 9653 7587 9667
rect 7633 9873 7647 9887
rect 7613 9613 7627 9627
rect 7813 10073 7827 10087
rect 7773 10054 7787 10068
rect 7853 10053 7867 10067
rect 7753 10012 7767 10026
rect 7793 10012 7807 10026
rect 7853 10012 7867 10026
rect 7753 9813 7767 9827
rect 7673 9753 7687 9767
rect 7833 9773 7847 9787
rect 7793 9754 7807 9768
rect 7733 9673 7747 9687
rect 7773 9593 7787 9607
rect 7693 9573 7707 9587
rect 7593 9534 7607 9548
rect 7633 9534 7647 9548
rect 7672 9534 7686 9548
rect 7353 9492 7367 9506
rect 7393 9492 7407 9506
rect 7433 9492 7447 9506
rect 7533 9492 7547 9506
rect 7513 9453 7527 9467
rect 7453 9333 7467 9347
rect 7353 9234 7367 9248
rect 7393 9234 7407 9248
rect 7313 9173 7327 9187
rect 7293 9133 7307 9147
rect 7273 9073 7287 9087
rect 7253 8994 7267 9008
rect 7293 8994 7307 9008
rect 7293 8933 7307 8947
rect 7273 8833 7287 8847
rect 7253 8813 7267 8827
rect 7213 8793 7227 8807
rect 7153 8773 7167 8787
rect 7193 8714 7207 8728
rect 7093 8672 7107 8686
rect 7073 8613 7087 8627
rect 7133 8613 7147 8627
rect 7233 8613 7247 8627
rect 7053 8453 7067 8467
rect 7093 8593 7107 8607
rect 7033 8333 7047 8347
rect 7073 8333 7087 8347
rect 7013 8253 7027 8267
rect 7033 8233 7047 8247
rect 7013 8213 7027 8227
rect 7053 8152 7067 8166
rect 7053 8131 7067 8145
rect 6993 8113 7007 8127
rect 7013 8073 7027 8087
rect 6973 7973 6987 7987
rect 6813 7952 6827 7966
rect 6813 7913 6827 7927
rect 6813 7892 6827 7906
rect 6633 7753 6647 7767
rect 6673 7753 6687 7767
rect 6793 7713 6807 7727
rect 6773 7613 6787 7627
rect 6793 7593 6807 7607
rect 6713 7533 6727 7547
rect 6653 7453 6667 7467
rect 6693 7454 6707 7468
rect 6753 7454 6767 7468
rect 6493 7373 6507 7387
rect 6453 7353 6467 7367
rect 6413 7253 6427 7267
rect 6493 7253 6507 7267
rect 6473 7233 6487 7247
rect 6393 7154 6407 7168
rect 6433 7154 6447 7168
rect 6333 7093 6347 7107
rect 6353 7053 6367 7067
rect 6333 7013 6347 7027
rect 6333 6973 6347 6987
rect 6333 6853 6347 6867
rect 6313 6813 6327 6827
rect 6413 7112 6427 7126
rect 6393 7053 6407 7067
rect 6553 7413 6567 7427
rect 6613 7413 6627 7427
rect 6533 7213 6547 7227
rect 6773 7412 6787 7426
rect 6973 7853 6987 7867
rect 6873 7733 6887 7747
rect 6933 7733 6947 7747
rect 6833 7674 6847 7688
rect 6893 7693 6907 7707
rect 6833 7453 6847 7467
rect 6873 7454 6887 7468
rect 6753 7313 6767 7327
rect 6733 7293 6747 7307
rect 6713 7253 6727 7267
rect 6653 7233 6667 7247
rect 6573 7213 6587 7227
rect 6553 7113 6567 7127
rect 6413 6953 6427 6967
rect 6473 6954 6487 6968
rect 6393 6893 6407 6907
rect 6373 6833 6387 6847
rect 6333 6773 6347 6787
rect 6253 6753 6267 6767
rect 6313 6753 6327 6767
rect 6233 6634 6247 6648
rect 6233 6593 6247 6607
rect 6092 6373 6106 6387
rect 6113 6373 6127 6387
rect 6073 6293 6087 6307
rect 6013 6233 6027 6247
rect 5953 6213 5967 6227
rect 5933 6134 5947 6148
rect 5873 5853 5887 5867
rect 5933 6073 5947 6087
rect 5913 5953 5927 5967
rect 5893 5813 5907 5827
rect 6093 6193 6107 6207
rect 6053 6173 6067 6187
rect 5993 6133 6007 6147
rect 6213 6333 6227 6347
rect 6153 6313 6167 6327
rect 6113 6153 6127 6167
rect 6173 6133 6187 6147
rect 6113 6114 6127 6128
rect 5973 6053 5987 6067
rect 6013 5953 6027 5967
rect 6353 6733 6367 6747
rect 6353 6653 6367 6667
rect 6313 6634 6327 6648
rect 6313 6573 6327 6587
rect 6313 6533 6327 6547
rect 6273 6413 6287 6427
rect 6373 6573 6387 6587
rect 6473 6933 6487 6947
rect 6493 6892 6507 6906
rect 6613 7173 6627 7187
rect 6653 7154 6667 7168
rect 6573 6892 6587 6906
rect 6633 7013 6647 7027
rect 6633 6953 6647 6967
rect 6613 6933 6627 6947
rect 6613 6892 6627 6906
rect 6413 6513 6427 6527
rect 6433 6453 6447 6467
rect 6393 6414 6407 6428
rect 6473 6833 6487 6847
rect 6473 6693 6487 6707
rect 6593 6873 6607 6887
rect 6613 6773 6627 6787
rect 6592 6733 6606 6747
rect 6613 6733 6627 6747
rect 6513 6653 6527 6667
rect 6573 6653 6587 6667
rect 6493 6634 6507 6648
rect 6473 6593 6487 6607
rect 6453 6433 6467 6447
rect 6373 6372 6387 6386
rect 6333 6353 6347 6367
rect 6253 6313 6267 6327
rect 6333 6313 6347 6327
rect 6233 6033 6247 6047
rect 6313 6033 6327 6047
rect 6293 5993 6307 6007
rect 6253 5953 6267 5967
rect 6073 5933 6087 5947
rect 6113 5933 6127 5947
rect 6213 5933 6227 5947
rect 6033 5913 6047 5927
rect 6053 5894 6067 5908
rect 5953 5733 5967 5747
rect 5893 5693 5907 5707
rect 5973 5653 5987 5667
rect 5853 5613 5867 5627
rect 5933 5594 5947 5608
rect 5853 5413 5867 5427
rect 5733 5233 5747 5247
rect 5693 5213 5707 5227
rect 5753 5213 5767 5227
rect 5593 4873 5607 4887
rect 5573 4853 5587 4867
rect 5673 4913 5687 4927
rect 5593 4834 5607 4848
rect 5453 4812 5467 4826
rect 5433 4573 5447 4587
rect 5413 4253 5427 4267
rect 5553 4812 5567 4826
rect 5513 4673 5527 4687
rect 5453 4513 5467 4527
rect 5493 4513 5507 4527
rect 5573 4653 5587 4667
rect 5553 4613 5567 4627
rect 5573 4573 5587 4587
rect 5593 4554 5607 4568
rect 5633 4554 5647 4568
rect 5573 4512 5587 4526
rect 5793 5113 5807 5127
rect 5913 5552 5927 5566
rect 6053 5793 6067 5807
rect 6093 5673 6107 5687
rect 6133 5913 6147 5927
rect 6113 5653 6127 5667
rect 6033 5633 6047 5647
rect 6073 5633 6087 5647
rect 6213 5912 6227 5926
rect 6173 5894 6187 5908
rect 6273 5933 6287 5947
rect 6253 5893 6267 5907
rect 6233 5852 6247 5866
rect 6273 5852 6287 5866
rect 6193 5813 6207 5827
rect 6213 5653 6227 5667
rect 5993 5594 6007 5608
rect 6013 5553 6027 5567
rect 5973 5473 5987 5487
rect 5873 5293 5887 5307
rect 5973 5374 5987 5388
rect 6093 5513 6107 5527
rect 6053 5473 6067 5487
rect 5953 5332 5967 5346
rect 5993 5332 6007 5346
rect 6033 5332 6047 5346
rect 6113 5433 6127 5447
rect 6113 5373 6127 5387
rect 6093 5332 6107 5346
rect 5973 5293 5987 5307
rect 5913 5253 5927 5267
rect 5853 5233 5867 5247
rect 5853 5113 5867 5127
rect 5813 5073 5827 5087
rect 5853 5074 5867 5088
rect 5793 5013 5807 5027
rect 5933 5073 5947 5087
rect 5933 5032 5947 5046
rect 5753 4933 5767 4947
rect 5913 4933 5927 4947
rect 5933 4873 5947 4887
rect 5833 4832 5847 4846
rect 5933 4832 5947 4846
rect 6113 5273 6127 5287
rect 5993 5133 6007 5147
rect 6053 5093 6067 5107
rect 6093 5074 6107 5088
rect 5993 5053 6007 5067
rect 6033 5032 6047 5046
rect 6073 5032 6087 5046
rect 6033 4933 6047 4947
rect 5973 4893 5987 4907
rect 5933 4793 5947 4807
rect 5853 4713 5867 4727
rect 5813 4693 5827 4707
rect 5713 4573 5727 4587
rect 5733 4554 5747 4568
rect 5773 4554 5787 4568
rect 5913 4693 5927 4707
rect 5713 4513 5727 4527
rect 5633 4413 5647 4427
rect 5513 4393 5527 4407
rect 5593 4393 5607 4407
rect 5453 4373 5467 4387
rect 5513 4334 5527 4348
rect 5553 4334 5567 4348
rect 5453 4313 5467 4327
rect 5733 4373 5747 4387
rect 5653 4333 5667 4347
rect 5713 4334 5727 4348
rect 5793 4512 5807 4526
rect 5833 4393 5847 4407
rect 5813 4334 5827 4348
rect 5853 4313 5867 4327
rect 5493 4292 5507 4306
rect 5533 4292 5547 4306
rect 5593 4292 5607 4306
rect 5653 4292 5667 4306
rect 5733 4292 5747 4306
rect 5453 4273 5467 4287
rect 5433 4193 5447 4207
rect 5333 4033 5347 4047
rect 5313 3813 5327 3827
rect 5193 3773 5207 3787
rect 5233 3772 5247 3786
rect 5333 3772 5347 3786
rect 5753 4253 5767 4267
rect 5573 4193 5587 4207
rect 5553 4173 5567 4187
rect 5493 4093 5507 4107
rect 5553 4093 5567 4107
rect 5453 4034 5467 4048
rect 5473 3973 5487 3987
rect 5433 3953 5447 3967
rect 5513 3853 5527 3867
rect 5393 3814 5407 3828
rect 5473 3814 5487 3828
rect 5473 3753 5487 3767
rect 5553 3733 5567 3747
rect 5493 3713 5507 3727
rect 5473 3693 5487 3707
rect 5553 3693 5567 3707
rect 5453 3653 5467 3667
rect 5392 3633 5406 3647
rect 5413 3633 5427 3647
rect 5293 3472 5307 3486
rect 5273 3433 5287 3447
rect 5313 3433 5327 3447
rect 5233 3393 5247 3407
rect 5193 3294 5207 3308
rect 5273 3333 5287 3347
rect 5173 3093 5187 3107
rect 5053 2994 5067 3008
rect 5133 2994 5147 3008
rect 5173 2994 5187 3008
rect 5052 2913 5066 2927
rect 5073 2913 5087 2927
rect 5053 2673 5067 2687
rect 5033 2393 5047 2407
rect 4973 2373 4987 2387
rect 4953 2313 4967 2327
rect 5033 2272 5047 2286
rect 4933 2254 4947 2268
rect 4973 2254 4987 2268
rect 5013 2254 5027 2268
rect 4933 2053 4947 2067
rect 4893 1954 4907 1968
rect 4993 2193 5007 2207
rect 4992 2113 5006 2127
rect 5013 2113 5027 2127
rect 5013 2073 5027 2087
rect 4953 1993 4967 2007
rect 4993 1953 5007 1967
rect 4873 1913 4887 1927
rect 4913 1873 4927 1887
rect 4933 1853 4947 1867
rect 4913 1833 4927 1847
rect 4873 1733 4887 1747
rect 4733 1713 4747 1727
rect 4713 1673 4727 1687
rect 4693 1613 4707 1627
rect 4653 1573 4667 1587
rect 4613 1533 4627 1547
rect 4593 1493 4607 1507
rect 4573 1453 4587 1467
rect 4613 1453 4627 1467
rect 4533 1293 4547 1307
rect 4513 1234 4527 1248
rect 4513 1213 4527 1227
rect 4553 1213 4567 1227
rect 4553 1153 4567 1167
rect 4553 1113 4567 1127
rect 4553 1053 4567 1067
rect 4593 1333 4607 1347
rect 4613 1273 4627 1287
rect 4593 1073 4607 1087
rect 4573 1013 4587 1027
rect 4493 933 4507 947
rect 4433 914 4447 928
rect 4393 872 4407 886
rect 4453 872 4467 886
rect 4493 773 4507 787
rect 4373 733 4387 747
rect 4333 694 4347 708
rect 4393 652 4407 666
rect 4333 633 4347 647
rect 4433 633 4447 647
rect 4293 613 4307 627
rect 4333 593 4347 607
rect 4353 473 4367 487
rect 4233 433 4247 447
rect 4173 233 4187 247
rect 4093 174 4107 188
rect 4133 174 4147 188
rect 4173 174 4187 188
rect 3493 132 3507 146
rect 2753 113 2767 127
rect 1733 73 1747 87
rect 1853 73 1867 87
rect 1953 73 1967 87
rect 3713 132 3727 146
rect 3753 132 3767 146
rect 4313 393 4327 407
rect 4453 413 4467 427
rect 4393 394 4407 408
rect 4693 1513 4707 1527
rect 4853 1713 4867 1727
rect 4833 1653 4847 1667
rect 4893 1673 4907 1687
rect 4873 1613 4887 1627
rect 4832 1573 4846 1587
rect 4853 1573 4867 1587
rect 4793 1553 4807 1567
rect 4773 1533 4787 1547
rect 4733 1453 4747 1467
rect 4713 1434 4727 1448
rect 4813 1493 4827 1507
rect 4793 1453 4807 1467
rect 4813 1434 4827 1448
rect 4873 1473 4887 1487
rect 4813 1313 4827 1327
rect 4853 1313 4867 1327
rect 4793 1273 4807 1287
rect 4733 1253 4747 1267
rect 4773 1253 4787 1267
rect 4793 1213 4807 1227
rect 4693 1172 4707 1186
rect 4733 1172 4747 1186
rect 4773 1172 4787 1186
rect 4653 1073 4667 1087
rect 4793 1153 4807 1167
rect 4753 1133 4767 1147
rect 4713 1073 4727 1087
rect 4693 1013 4707 1027
rect 4613 913 4627 927
rect 4633 872 4647 886
rect 4673 872 4687 886
rect 4733 893 4747 907
rect 4613 813 4627 827
rect 4713 813 4727 827
rect 4593 713 4607 727
rect 4513 694 4527 708
rect 4573 694 4587 708
rect 4653 713 4667 727
rect 4513 613 4527 627
rect 4593 652 4607 666
rect 4653 652 4667 666
rect 4613 613 4627 627
rect 4553 533 4567 547
rect 4933 1753 4947 1767
rect 4933 1732 4947 1746
rect 4933 1573 4947 1587
rect 4933 1493 4947 1507
rect 4913 1473 4927 1487
rect 4993 1793 5007 1807
rect 5013 1713 5027 1727
rect 4993 1573 5007 1587
rect 4973 1553 4987 1567
rect 5013 1493 5027 1507
rect 5193 2952 5207 2966
rect 5193 2873 5207 2887
rect 5113 2793 5127 2807
rect 5153 2793 5167 2807
rect 5173 2773 5187 2787
rect 5093 2732 5107 2746
rect 5113 2713 5127 2727
rect 5093 2473 5107 2487
rect 5093 2413 5107 2427
rect 5153 2593 5167 2607
rect 5213 2774 5227 2788
rect 5273 3233 5287 3247
rect 5253 2932 5267 2946
rect 5253 2713 5267 2727
rect 5293 3173 5307 3187
rect 5293 3073 5307 3087
rect 5333 3313 5347 3327
rect 5313 2873 5327 2887
rect 5293 2853 5307 2867
rect 5313 2833 5327 2847
rect 5293 2793 5307 2807
rect 5273 2693 5287 2707
rect 5233 2633 5247 2647
rect 5273 2633 5287 2647
rect 5233 2593 5247 2607
rect 5193 2553 5207 2567
rect 5213 2533 5227 2547
rect 5173 2493 5187 2507
rect 5193 2473 5207 2487
rect 5153 2432 5167 2446
rect 5113 2313 5127 2327
rect 5073 2213 5087 2227
rect 5053 1833 5067 1847
rect 5073 1773 5087 1787
rect 5173 2273 5187 2287
rect 5253 2513 5267 2527
rect 5233 2253 5247 2267
rect 5193 2212 5207 2226
rect 5153 2173 5167 2187
rect 5173 2153 5187 2167
rect 5153 2093 5167 2107
rect 5152 1954 5166 1968
rect 5193 2053 5207 2067
rect 5173 1953 5187 1967
rect 5193 1932 5207 1946
rect 5273 2252 5287 2266
rect 5273 2173 5287 2187
rect 5373 3373 5387 3387
rect 5373 3173 5387 3187
rect 5373 3152 5387 3166
rect 5433 3553 5447 3567
rect 5413 3333 5427 3347
rect 5513 3533 5527 3547
rect 5593 4153 5607 4167
rect 5533 3472 5547 3486
rect 5453 3313 5467 3327
rect 5613 3893 5627 3907
rect 5493 3294 5507 3308
rect 5553 3293 5567 3307
rect 5593 3294 5607 3308
rect 5513 3252 5527 3266
rect 5473 3233 5487 3247
rect 5553 3173 5567 3187
rect 5753 3993 5767 4007
rect 5713 3973 5727 3987
rect 5813 4293 5827 4307
rect 5793 4233 5807 4247
rect 5793 3893 5807 3907
rect 5673 3853 5687 3867
rect 5693 3833 5707 3847
rect 5733 3814 5747 3828
rect 5793 3814 5807 3828
rect 5713 3772 5727 3786
rect 5753 3733 5767 3747
rect 5693 3693 5707 3707
rect 5673 3573 5687 3587
rect 5633 3533 5647 3547
rect 5653 3353 5667 3367
rect 5633 3253 5647 3267
rect 5613 3113 5627 3127
rect 5473 3073 5487 3087
rect 5593 3073 5607 3087
rect 5433 3033 5447 3047
rect 5393 3013 5407 3027
rect 5393 2913 5407 2927
rect 5373 2893 5387 2907
rect 5332 2793 5346 2807
rect 5353 2793 5367 2807
rect 5653 3213 5667 3227
rect 5573 2952 5587 2966
rect 5553 2933 5567 2947
rect 5513 2893 5527 2907
rect 5353 2732 5367 2746
rect 5393 2693 5407 2707
rect 5313 2473 5327 2487
rect 5373 2474 5387 2488
rect 5353 2432 5367 2446
rect 5393 2432 5407 2446
rect 5453 2773 5467 2787
rect 5453 2732 5467 2746
rect 5373 2373 5387 2387
rect 5433 2373 5447 2387
rect 5333 2293 5347 2307
rect 5253 2093 5267 2107
rect 5533 2873 5547 2887
rect 5613 2873 5627 2887
rect 5513 2293 5527 2307
rect 5393 2254 5407 2268
rect 5433 2254 5447 2268
rect 5493 2253 5507 2267
rect 5413 2173 5427 2187
rect 5353 2153 5367 2167
rect 5613 2793 5627 2807
rect 5573 2774 5587 2788
rect 5633 2732 5647 2746
rect 5593 2673 5607 2687
rect 5573 2653 5587 2667
rect 5773 3653 5787 3667
rect 5733 3514 5747 3528
rect 5833 4173 5847 4187
rect 5993 4753 6007 4767
rect 6033 4753 6047 4767
rect 6113 4973 6127 4987
rect 6173 5513 6187 5527
rect 6173 5374 6187 5388
rect 6193 5332 6207 5346
rect 6253 5733 6267 5747
rect 6353 6193 6367 6207
rect 6333 5733 6347 5747
rect 6333 5673 6347 5687
rect 6413 6233 6427 6247
rect 6393 6153 6407 6167
rect 6373 6073 6387 6087
rect 6393 5993 6407 6007
rect 6493 6333 6507 6347
rect 6473 6193 6487 6207
rect 6473 6114 6487 6128
rect 6553 6592 6567 6606
rect 6573 6553 6587 6567
rect 6553 6513 6567 6527
rect 6533 6372 6547 6386
rect 6532 6153 6546 6167
rect 6553 6153 6567 6167
rect 6493 6072 6507 6086
rect 6413 5953 6427 5967
rect 6373 5893 6387 5907
rect 6433 5894 6447 5908
rect 6453 5852 6467 5866
rect 6413 5813 6427 5827
rect 6373 5673 6387 5687
rect 6353 5653 6367 5667
rect 6493 5773 6507 5787
rect 6453 5753 6467 5767
rect 6493 5752 6507 5766
rect 6433 5673 6447 5687
rect 6373 5613 6387 5627
rect 6413 5613 6427 5627
rect 6473 5653 6487 5667
rect 6453 5593 6467 5607
rect 6353 5552 6367 5566
rect 6313 5533 6327 5547
rect 6333 5513 6347 5527
rect 6253 5413 6267 5427
rect 6193 5273 6207 5287
rect 6173 5253 6187 5267
rect 6153 4973 6167 4987
rect 6153 4952 6167 4966
rect 6133 4913 6147 4927
rect 6113 4893 6127 4907
rect 6053 4693 6067 4707
rect 6013 4613 6027 4627
rect 5953 4593 5967 4607
rect 5953 4553 5967 4567
rect 6113 4673 6127 4687
rect 6113 4613 6127 4627
rect 6073 4553 6087 4567
rect 5993 4533 6007 4547
rect 5933 4493 5947 4507
rect 5973 4393 5987 4407
rect 6073 4493 6087 4507
rect 6033 4353 6047 4367
rect 6013 4334 6027 4348
rect 5913 4193 5927 4207
rect 6293 5093 6307 5107
rect 6353 5433 6367 5447
rect 6473 5552 6487 5566
rect 6453 5433 6467 5447
rect 6353 5373 6367 5387
rect 6393 5373 6407 5387
rect 6433 5374 6447 5388
rect 6473 5373 6487 5387
rect 6353 5293 6367 5307
rect 6333 5253 6347 5267
rect 6333 5193 6347 5207
rect 6313 5073 6327 5087
rect 6273 5032 6287 5046
rect 6212 4953 6226 4967
rect 6233 4953 6247 4967
rect 6233 4913 6247 4927
rect 6193 4873 6207 4887
rect 6153 4833 6167 4847
rect 6253 4812 6267 4826
rect 6313 4793 6327 4807
rect 6173 4673 6187 4687
rect 6173 4413 6187 4427
rect 6313 4653 6327 4667
rect 6333 4593 6347 4607
rect 6293 4512 6307 4526
rect 6253 4493 6267 4507
rect 6333 4433 6347 4447
rect 6313 4393 6327 4407
rect 6153 4293 6167 4307
rect 6213 4253 6227 4267
rect 6133 4233 6147 4247
rect 5993 4213 6007 4227
rect 6093 4193 6107 4207
rect 5953 4113 5967 4127
rect 6013 4113 6027 4127
rect 5853 4093 5867 4107
rect 5893 4093 5907 4107
rect 5873 4073 5887 4087
rect 5853 4033 5867 4047
rect 5853 3893 5867 3907
rect 5833 3773 5847 3787
rect 5813 3573 5827 3587
rect 5793 3533 5807 3547
rect 5893 4033 5907 4047
rect 5933 3992 5947 4006
rect 5893 3893 5907 3907
rect 5973 3853 5987 3867
rect 5933 3814 5947 3828
rect 5892 3693 5906 3707
rect 5913 3693 5927 3707
rect 6033 4073 6047 4087
rect 6073 3893 6087 3907
rect 6033 3814 6047 3828
rect 6113 4033 6127 4047
rect 6152 4034 6166 4048
rect 6213 4073 6227 4087
rect 6173 4033 6187 4047
rect 6193 3992 6207 4006
rect 6133 3953 6147 3967
rect 6113 3913 6127 3927
rect 6093 3814 6107 3828
rect 6133 3814 6147 3828
rect 6173 3814 6187 3828
rect 6273 3913 6287 3927
rect 6233 3813 6247 3827
rect 6073 3793 6087 3807
rect 6153 3753 6167 3767
rect 6273 3733 6287 3747
rect 6013 3653 6027 3667
rect 5913 3633 5927 3647
rect 5973 3633 5987 3647
rect 6233 3633 6247 3647
rect 5933 3613 5947 3627
rect 5873 3553 5887 3567
rect 5693 3433 5707 3447
rect 5753 3393 5767 3407
rect 5733 3294 5747 3308
rect 5693 3252 5707 3266
rect 5713 3113 5727 3127
rect 5693 2813 5707 2827
rect 5693 2732 5707 2746
rect 5573 2533 5587 2547
rect 5673 2533 5687 2547
rect 5593 2474 5607 2488
rect 5693 2474 5707 2488
rect 5693 2313 5707 2327
rect 5653 2293 5667 2307
rect 5833 3433 5847 3447
rect 5853 3373 5867 3387
rect 5793 3253 5807 3267
rect 6233 3573 6247 3587
rect 6273 3573 6287 3587
rect 6073 3494 6087 3508
rect 6193 3492 6207 3506
rect 5893 3473 5907 3487
rect 6173 3433 6187 3447
rect 5893 3393 5907 3407
rect 5913 3373 5927 3387
rect 5953 3294 5967 3308
rect 6073 3293 6087 3307
rect 6193 3294 6207 3308
rect 5933 3213 5947 3227
rect 5873 3133 5887 3147
rect 5913 3033 5927 3047
rect 5833 2994 5847 3008
rect 5933 3013 5947 3027
rect 5813 2952 5827 2966
rect 5853 2952 5867 2966
rect 5773 2933 5787 2947
rect 5853 2913 5867 2927
rect 5753 2774 5767 2788
rect 5793 2774 5807 2788
rect 5813 2713 5827 2727
rect 5793 2693 5807 2707
rect 5833 2693 5847 2707
rect 5753 2593 5767 2607
rect 5753 2474 5767 2488
rect 5793 2474 5807 2488
rect 5833 2353 5847 2367
rect 5753 2293 5767 2307
rect 5793 2293 5807 2307
rect 5713 2273 5727 2287
rect 5773 2272 5787 2286
rect 5573 2213 5587 2227
rect 5753 2213 5767 2227
rect 5533 2173 5547 2187
rect 5673 2173 5687 2187
rect 5533 2133 5547 2147
rect 5493 2113 5507 2127
rect 5273 2073 5287 2087
rect 5333 2073 5347 2087
rect 5493 2073 5507 2087
rect 5293 2033 5307 2047
rect 5433 2033 5447 2047
rect 5273 1973 5287 1987
rect 5133 1873 5147 1887
rect 5213 1873 5227 1887
rect 5193 1833 5207 1847
rect 5093 1753 5107 1767
rect 5153 1753 5167 1767
rect 5113 1734 5127 1748
rect 5093 1692 5107 1706
rect 5053 1653 5067 1667
rect 5053 1613 5067 1627
rect 5133 1593 5147 1607
rect 5033 1433 5047 1447
rect 5073 1433 5087 1447
rect 4853 1273 4867 1287
rect 4893 1273 4907 1287
rect 4813 1113 4827 1127
rect 4833 1033 4847 1047
rect 4913 1233 4927 1247
rect 4873 1172 4887 1186
rect 4933 1053 4947 1067
rect 4853 993 4867 1007
rect 4893 993 4907 1007
rect 4893 953 4907 967
rect 4833 933 4847 947
rect 4813 914 4827 928
rect 4853 914 4867 928
rect 4753 872 4767 886
rect 4813 833 4827 847
rect 4813 773 4827 787
rect 4813 713 4827 727
rect 4793 633 4807 647
rect 4833 433 4847 447
rect 4733 413 4747 427
rect 4993 1293 5007 1307
rect 5013 1253 5027 1267
rect 4993 1233 5007 1247
rect 4493 373 4507 387
rect 4373 352 4387 366
rect 4313 293 4327 307
rect 4253 173 4267 187
rect 4293 173 4307 187
rect 3933 132 3947 146
rect 4193 132 4207 146
rect 4233 132 4247 146
rect 4153 113 4167 127
rect 3793 93 3807 107
rect 4453 352 4467 366
rect 4413 253 4427 267
rect 4373 174 4387 188
rect 4413 174 4427 188
rect 4473 174 4487 188
rect 4313 132 4327 146
rect 4393 132 4407 146
rect 4433 132 4447 146
rect 4293 113 4307 127
rect 4253 73 4267 87
rect 5113 1393 5127 1407
rect 5133 1373 5147 1387
rect 5073 1353 5087 1367
rect 5113 1353 5127 1367
rect 5073 1313 5087 1327
rect 5173 1734 5187 1748
rect 5273 1933 5287 1947
rect 5253 1853 5267 1867
rect 5293 1893 5307 1907
rect 5373 1833 5387 1847
rect 5293 1773 5307 1787
rect 5233 1753 5247 1767
rect 5273 1753 5287 1767
rect 5213 1713 5227 1727
rect 5193 1693 5207 1707
rect 5173 1513 5187 1527
rect 5333 1753 5347 1767
rect 5593 2013 5607 2027
rect 5653 2013 5667 2027
rect 5633 1953 5647 1967
rect 5553 1932 5567 1946
rect 5613 1933 5627 1947
rect 5593 1773 5607 1787
rect 5533 1753 5547 1767
rect 5573 1753 5587 1767
rect 5513 1734 5527 1748
rect 5493 1713 5507 1727
rect 5313 1692 5327 1706
rect 5373 1692 5387 1706
rect 5393 1673 5407 1687
rect 5273 1633 5287 1647
rect 5493 1613 5507 1627
rect 5393 1553 5407 1567
rect 5233 1493 5247 1507
rect 5293 1493 5307 1507
rect 5553 1493 5567 1507
rect 5233 1453 5247 1467
rect 5173 1273 5187 1287
rect 5073 1193 5087 1207
rect 5253 1233 5267 1247
rect 5073 1113 5087 1127
rect 5113 1013 5127 1027
rect 5193 1113 5207 1127
rect 5173 993 5187 1007
rect 5113 933 5127 947
rect 5153 933 5167 947
rect 5073 914 5087 928
rect 5093 872 5107 886
rect 5153 793 5167 807
rect 4973 713 4987 727
rect 5053 713 5067 727
rect 4993 693 5007 707
rect 5033 694 5047 708
rect 4973 652 4987 666
rect 5053 652 5067 666
rect 5133 413 5147 427
rect 5053 394 5067 408
rect 4513 352 4527 366
rect 4593 352 4607 366
rect 4633 352 4647 366
rect 4813 352 4827 366
rect 4633 313 4647 327
rect 4813 313 4827 327
rect 4893 352 4907 366
rect 4933 352 4947 366
rect 5073 352 5087 366
rect 5093 333 5107 347
rect 5033 313 5047 327
rect 4813 273 4827 287
rect 4853 273 4867 287
rect 4893 253 4907 267
rect 4653 193 4667 207
rect 4613 174 4627 188
rect 4953 193 4967 207
rect 4893 174 4907 188
rect 4953 174 4967 188
rect 5093 174 5107 188
rect 4493 133 4507 147
rect 5372 1473 5386 1487
rect 5393 1473 5407 1487
rect 5373 1392 5387 1406
rect 5333 1293 5347 1307
rect 5453 1434 5467 1448
rect 5533 1433 5547 1447
rect 5433 1392 5447 1406
rect 5473 1293 5487 1307
rect 5473 1233 5487 1247
rect 5433 1214 5447 1228
rect 5333 1193 5347 1207
rect 5553 1333 5567 1347
rect 5493 1213 5507 1227
rect 5533 1214 5547 1228
rect 5373 1172 5387 1186
rect 5413 1172 5427 1186
rect 5473 1172 5487 1186
rect 5333 1033 5347 1047
rect 5373 933 5387 947
rect 5353 872 5367 886
rect 5313 793 5327 807
rect 5273 713 5287 727
rect 5333 713 5347 727
rect 5253 694 5267 708
rect 5273 652 5287 666
rect 5233 593 5247 607
rect 5253 433 5267 447
rect 5193 393 5207 407
rect 5293 394 5307 408
rect 5193 352 5207 366
rect 5273 352 5287 366
rect 5233 273 5247 287
rect 5173 253 5187 267
rect 5153 174 5167 188
rect 5213 174 5227 188
rect 4853 132 4867 146
rect 4913 132 4927 146
rect 5133 132 5147 146
rect 4633 93 4647 107
rect 5313 133 5327 147
rect 5233 113 5247 127
rect 1573 53 1587 67
rect 3553 53 3567 67
rect 4473 53 4487 67
rect 5173 53 5187 67
rect 5513 1193 5527 1207
rect 5513 1153 5527 1167
rect 5513 973 5527 987
rect 5633 1833 5647 1847
rect 5653 1653 5667 1667
rect 5713 2193 5727 2207
rect 5713 2053 5727 2067
rect 5732 2033 5746 2047
rect 5753 2033 5767 2047
rect 5733 1933 5747 1947
rect 5813 2254 5827 2268
rect 5793 2193 5807 2207
rect 5773 1993 5787 2007
rect 5813 2133 5827 2147
rect 5793 1954 5807 1968
rect 5893 2474 5907 2488
rect 5993 2994 6007 3008
rect 6293 3493 6307 3507
rect 6273 3273 6287 3287
rect 6473 5332 6487 5346
rect 6493 5293 6507 5307
rect 6473 5253 6487 5267
rect 6453 5233 6467 5247
rect 6373 5153 6387 5167
rect 6393 5133 6407 5147
rect 6473 5133 6487 5147
rect 6473 5112 6487 5126
rect 6553 5973 6567 5987
rect 6533 5953 6547 5967
rect 6553 5852 6567 5866
rect 6653 6773 6667 6787
rect 6653 6752 6667 6766
rect 6653 6593 6667 6607
rect 6633 6493 6647 6507
rect 6613 6453 6627 6467
rect 6613 6414 6627 6428
rect 6773 7193 6787 7207
rect 6813 7373 6827 7387
rect 6813 7333 6827 7347
rect 6973 7674 6987 7688
rect 6953 7632 6967 7646
rect 7033 8033 7047 8047
rect 7033 7933 7047 7947
rect 7033 7674 7047 7688
rect 7033 7633 7047 7647
rect 6913 7533 6927 7547
rect 6953 7454 6967 7468
rect 6993 7454 7007 7468
rect 6913 7412 6927 7426
rect 7013 7412 7027 7426
rect 7173 8573 7187 8587
rect 7213 8494 7227 8508
rect 7113 8452 7127 8466
rect 7233 8452 7247 8466
rect 7193 8393 7207 8407
rect 7133 8373 7147 8387
rect 7133 8313 7147 8327
rect 7112 8233 7126 8247
rect 7133 8233 7147 8247
rect 7113 8152 7127 8166
rect 7173 8213 7187 8227
rect 7133 8093 7147 8107
rect 7113 8013 7127 8027
rect 7293 8713 7307 8727
rect 7273 8553 7287 8567
rect 7293 8513 7307 8527
rect 7273 8494 7287 8508
rect 7313 8393 7327 8407
rect 7293 8293 7307 8307
rect 7253 8213 7267 8227
rect 7273 8194 7287 8208
rect 7273 8093 7287 8107
rect 7253 8073 7267 8087
rect 7253 8033 7267 8047
rect 7173 7993 7187 8007
rect 7092 7773 7106 7787
rect 7113 7773 7127 7787
rect 7113 7713 7127 7727
rect 7253 7853 7267 7867
rect 7073 7693 7087 7707
rect 7133 7674 7147 7688
rect 7173 7674 7187 7688
rect 7233 7674 7247 7688
rect 7213 7633 7227 7647
rect 7313 8153 7327 8167
rect 7353 9093 7367 9107
rect 7413 9133 7427 9147
rect 7393 9073 7407 9087
rect 7373 9053 7387 9067
rect 7373 9014 7387 9028
rect 7353 8753 7367 8767
rect 7373 8733 7387 8747
rect 7493 9293 7507 9307
rect 7453 9014 7467 9028
rect 7493 9013 7507 9027
rect 7473 8972 7487 8986
rect 7613 9492 7627 9506
rect 7613 9234 7627 9248
rect 7553 9192 7567 9206
rect 7533 9073 7547 9087
rect 7573 9173 7587 9187
rect 7553 8973 7567 8987
rect 7433 8873 7447 8887
rect 7393 8714 7407 8728
rect 7453 8853 7467 8867
rect 7453 8673 7467 8687
rect 7433 8653 7447 8667
rect 7513 8913 7527 8927
rect 7513 8753 7527 8767
rect 7533 8713 7547 8727
rect 7693 9533 7707 9547
rect 7833 9534 7847 9548
rect 7893 10313 7907 10327
rect 7953 10533 7967 10547
rect 8073 10613 8087 10627
rect 8093 10593 8107 10607
rect 8173 10653 8187 10667
rect 8233 10752 8247 10766
rect 8333 11033 8347 11047
rect 8713 11033 8727 11047
rect 8533 11013 8547 11027
rect 8873 11052 8887 11066
rect 8933 11052 8947 11066
rect 8973 11013 8987 11027
rect 9073 10993 9087 11007
rect 8753 10953 8767 10967
rect 9033 10953 9047 10967
rect 8393 10873 8407 10887
rect 8353 10813 8367 10827
rect 8333 10793 8347 10807
rect 8193 10633 8207 10647
rect 8173 10573 8187 10587
rect 8033 10532 8047 10546
rect 8113 10532 8127 10546
rect 8213 10493 8227 10507
rect 8153 10373 8167 10387
rect 8113 10313 8127 10327
rect 7913 10273 7927 10287
rect 7933 10274 7947 10288
rect 7953 10232 7967 10246
rect 8313 10753 8327 10767
rect 8333 10713 8347 10727
rect 8313 10593 8327 10607
rect 8453 10853 8467 10867
rect 8513 10853 8527 10867
rect 8493 10813 8507 10827
rect 8593 10833 8607 10847
rect 8733 10833 8747 10847
rect 8513 10794 8527 10808
rect 8393 10752 8407 10766
rect 8433 10752 8447 10766
rect 8473 10633 8487 10647
rect 8553 10593 8567 10607
rect 8553 10574 8567 10588
rect 8693 10794 8707 10808
rect 8933 10794 8947 10808
rect 8653 10752 8667 10766
rect 8673 10693 8687 10707
rect 8653 10673 8667 10687
rect 8333 10532 8347 10546
rect 8433 10532 8447 10546
rect 8573 10513 8587 10527
rect 8913 10752 8927 10766
rect 8953 10752 8967 10766
rect 9033 10793 9047 10807
rect 8833 10713 8847 10727
rect 9013 10713 9027 10727
rect 8713 10653 8727 10667
rect 8753 10574 8767 10588
rect 8793 10574 8807 10588
rect 9073 10753 9087 10767
rect 8733 10553 8747 10567
rect 8673 10513 8687 10527
rect 8733 10493 8747 10507
rect 8653 10473 8667 10487
rect 8893 10573 8907 10587
rect 8773 10533 8787 10547
rect 8853 10532 8867 10546
rect 8893 10532 8907 10546
rect 8813 10473 8827 10487
rect 8732 10453 8746 10467
rect 8753 10453 8767 10467
rect 8373 10373 8387 10387
rect 8613 10373 8627 10387
rect 8273 10313 8287 10327
rect 8453 10313 8467 10327
rect 8593 10313 8607 10327
rect 8493 10274 8507 10288
rect 8193 10213 8207 10227
rect 8173 10193 8187 10207
rect 8133 10173 8147 10187
rect 8173 10153 8187 10167
rect 8113 10133 8127 10147
rect 7993 10054 8007 10068
rect 8313 10153 8327 10167
rect 8293 10133 8307 10147
rect 8233 10054 8247 10068
rect 8313 10113 8327 10127
rect 8313 10053 8327 10067
rect 8353 10054 8367 10068
rect 7933 9973 7947 9987
rect 7913 9853 7927 9867
rect 7853 9492 7867 9506
rect 7813 9413 7827 9427
rect 7993 9933 8007 9947
rect 7973 9853 7987 9867
rect 8213 10012 8227 10026
rect 8293 10012 8307 10026
rect 8253 9973 8267 9987
rect 8013 9913 8027 9927
rect 8013 9873 8027 9887
rect 8053 9754 8067 9768
rect 8153 9754 8167 9768
rect 8193 9754 8207 9768
rect 8233 9754 8247 9768
rect 7973 9712 7987 9726
rect 7913 9393 7927 9407
rect 7833 9273 7847 9287
rect 7913 9273 7927 9287
rect 7893 9253 7907 9267
rect 7813 9192 7827 9206
rect 7853 9192 7867 9206
rect 7953 9234 7967 9248
rect 8393 10213 8407 10227
rect 8693 10293 8707 10307
rect 8653 10274 8667 10288
rect 8433 10193 8447 10207
rect 8493 10193 8507 10207
rect 8533 10193 8547 10207
rect 8473 10113 8487 10127
rect 8433 10054 8447 10068
rect 8373 10012 8387 10026
rect 8453 10012 8467 10026
rect 8353 9973 8367 9987
rect 8433 9953 8447 9967
rect 8493 9953 8507 9967
rect 8373 9933 8387 9947
rect 8453 9793 8467 9807
rect 8513 9754 8527 9768
rect 8153 9653 8167 9667
rect 8113 9633 8127 9647
rect 8053 9593 8067 9607
rect 8113 9553 8127 9567
rect 8093 9534 8107 9548
rect 8253 9712 8267 9726
rect 8293 9712 8307 9726
rect 8433 9712 8447 9726
rect 8493 9712 8507 9726
rect 8473 9653 8487 9667
rect 8493 9633 8507 9647
rect 8253 9573 8267 9587
rect 8213 9513 8227 9527
rect 8113 9492 8127 9506
rect 8313 9553 8327 9567
rect 8453 9553 8467 9567
rect 8433 9513 8447 9527
rect 8253 9453 8267 9467
rect 8533 9573 8547 9587
rect 8593 10232 8607 10246
rect 8633 10232 8647 10246
rect 8713 10232 8727 10246
rect 8673 10193 8687 10207
rect 8753 10273 8767 10287
rect 8733 10193 8747 10207
rect 8713 10113 8727 10127
rect 8613 10053 8627 10067
rect 8673 10054 8687 10068
rect 8453 9492 8467 9506
rect 8513 9492 8527 9506
rect 8553 9492 8567 9506
rect 8593 9492 8607 9506
rect 8433 9453 8447 9467
rect 8293 9413 8307 9427
rect 8193 9353 8207 9367
rect 8073 9313 8087 9327
rect 8113 9313 8127 9327
rect 8073 9253 8087 9267
rect 7673 9173 7687 9187
rect 7653 9033 7667 9047
rect 7813 9033 7827 9047
rect 7713 9013 7727 9027
rect 7953 9193 7967 9207
rect 7973 9053 7987 9067
rect 7813 8972 7827 8986
rect 7593 8933 7607 8947
rect 7893 8972 7907 8986
rect 7633 8913 7647 8927
rect 7853 8913 7867 8927
rect 7673 8893 7687 8907
rect 7533 8672 7547 8686
rect 7373 8593 7387 8607
rect 7493 8593 7507 8607
rect 7353 8573 7367 8587
rect 7453 8553 7467 8567
rect 7533 8533 7547 8547
rect 7513 8453 7527 8467
rect 7393 8393 7407 8407
rect 7373 8353 7387 8367
rect 7353 8133 7367 8147
rect 7413 8253 7427 8267
rect 7493 8293 7507 8307
rect 7593 8672 7607 8686
rect 7773 8833 7787 8847
rect 7713 8773 7727 8787
rect 7693 8714 7707 8728
rect 7573 8653 7587 8667
rect 7553 8393 7567 8407
rect 7613 8613 7627 8627
rect 7593 8573 7607 8587
rect 7573 8353 7587 8367
rect 7533 8313 7547 8327
rect 7713 8673 7727 8687
rect 7733 8593 7747 8607
rect 7873 8773 7887 8787
rect 7833 8714 7847 8728
rect 8033 9234 8047 9248
rect 8273 9333 8287 9347
rect 8453 9333 8467 9347
rect 8193 9234 8207 9248
rect 8233 9234 8247 9248
rect 8413 9273 8427 9287
rect 8413 9234 8427 9248
rect 8533 9273 8547 9287
rect 8493 9234 8507 9248
rect 8053 9173 8067 9187
rect 8113 9173 8127 9187
rect 8013 9133 8027 9147
rect 8093 9093 8107 9107
rect 8153 9033 8167 9047
rect 8013 8972 8027 8986
rect 8073 8972 8087 8986
rect 8113 8972 8127 8986
rect 8153 8972 8167 8986
rect 8313 9053 8327 9067
rect 8253 9013 8267 9027
rect 8293 8972 8307 8986
rect 8513 9173 8527 9187
rect 8433 9153 8447 9167
rect 8273 8933 8287 8947
rect 8413 8933 8427 8947
rect 8193 8893 8207 8907
rect 8033 8833 8047 8847
rect 7993 8773 8007 8787
rect 7933 8692 7947 8706
rect 7973 8693 7987 8707
rect 7813 8673 7827 8687
rect 7733 8493 7747 8507
rect 7773 8493 7787 8507
rect 7753 8474 7767 8488
rect 7893 8593 7907 8607
rect 7993 8673 8007 8687
rect 8173 8733 8187 8747
rect 8033 8613 8047 8627
rect 7933 8573 7947 8587
rect 8232 8493 8246 8507
rect 8253 8493 8267 8507
rect 7673 8452 7687 8466
rect 7713 8452 7727 8466
rect 7673 8413 7687 8427
rect 7633 8373 7647 8387
rect 7853 8472 7867 8486
rect 7993 8472 8007 8486
rect 7833 8373 7847 8387
rect 7793 8313 7807 8327
rect 7593 8253 7607 8267
rect 7513 8233 7527 8247
rect 7533 8214 7547 8228
rect 7593 8214 7607 8228
rect 7433 8173 7447 8187
rect 7573 8172 7587 8186
rect 7693 8174 7707 8188
rect 7413 8113 7427 8127
rect 7513 8113 7527 8127
rect 7393 8093 7407 8107
rect 7353 8073 7367 8087
rect 7393 8072 7407 8086
rect 7373 8053 7387 8067
rect 7413 7974 7427 7988
rect 7453 7973 7467 7987
rect 7333 7893 7347 7907
rect 7313 7813 7327 7827
rect 7253 7633 7267 7647
rect 7193 7613 7207 7627
rect 7233 7613 7247 7627
rect 6893 7253 6907 7267
rect 7013 7213 7027 7227
rect 6893 7173 6907 7187
rect 6933 7173 6947 7187
rect 6853 7154 6867 7168
rect 6773 7112 6787 7126
rect 6833 7112 6847 7126
rect 6913 7112 6927 7126
rect 6893 7013 6907 7027
rect 6753 6993 6767 7007
rect 6833 6993 6847 7007
rect 6873 6993 6887 7007
rect 6693 6953 6707 6967
rect 6793 6934 6807 6948
rect 6893 6934 6907 6948
rect 6693 6892 6707 6906
rect 6833 6892 6847 6906
rect 6953 7154 6967 7168
rect 7013 7153 7027 7167
rect 6932 7073 6946 7087
rect 6953 7073 6967 7087
rect 7113 7513 7127 7527
rect 7093 7373 7107 7387
rect 7153 7553 7167 7567
rect 7133 7313 7147 7327
rect 7233 7533 7247 7547
rect 7273 7493 7287 7507
rect 7213 7293 7227 7307
rect 7153 7273 7167 7287
rect 7113 7233 7127 7247
rect 7053 7154 7067 7168
rect 7153 7112 7167 7126
rect 7113 7073 7127 7087
rect 7033 7053 7047 7067
rect 7153 7053 7167 7067
rect 7073 6953 7087 6967
rect 6933 6933 6947 6947
rect 6993 6934 7007 6948
rect 7033 6934 7047 6948
rect 6973 6892 6987 6906
rect 7013 6892 7027 6906
rect 6912 6833 6926 6847
rect 6933 6833 6947 6847
rect 6713 6773 6727 6787
rect 6693 6613 6707 6627
rect 7053 6753 7067 6767
rect 7013 6733 7027 6747
rect 7053 6713 7067 6727
rect 7033 6693 7047 6707
rect 6933 6653 6947 6667
rect 7033 6653 7047 6667
rect 6773 6634 6787 6648
rect 6813 6634 6827 6648
rect 6913 6613 6927 6627
rect 6673 6553 6687 6567
rect 6713 6553 6727 6567
rect 6753 6553 6767 6567
rect 6833 6593 6847 6607
rect 6813 6553 6827 6567
rect 6793 6513 6807 6527
rect 6753 6473 6767 6487
rect 6733 6433 6747 6447
rect 6633 6372 6647 6386
rect 6712 6293 6726 6307
rect 6733 6293 6747 6307
rect 6773 6453 6787 6467
rect 6773 6414 6787 6428
rect 6853 6553 6867 6567
rect 6913 6513 6927 6527
rect 6833 6493 6847 6507
rect 6973 6634 6987 6648
rect 7053 6573 7067 6587
rect 6933 6473 6947 6487
rect 7013 6433 7027 6447
rect 6893 6414 6907 6428
rect 7033 6413 7047 6427
rect 6753 6253 6767 6267
rect 6713 6233 6727 6247
rect 6633 6213 6647 6227
rect 6733 6213 6747 6227
rect 6613 6114 6627 6128
rect 6713 6193 6727 6207
rect 6733 6173 6747 6187
rect 6693 6114 6707 6128
rect 6633 6033 6647 6047
rect 6593 6013 6607 6027
rect 6573 5753 6587 5767
rect 6573 5732 6587 5746
rect 6533 5513 6547 5527
rect 6533 5473 6547 5487
rect 6533 5193 6547 5207
rect 6533 5113 6547 5127
rect 6513 5093 6527 5107
rect 6413 4933 6427 4947
rect 6453 5033 6467 5047
rect 6433 4913 6447 4927
rect 6493 5032 6507 5046
rect 6473 5013 6487 5027
rect 6513 4953 6527 4967
rect 6473 4853 6487 4867
rect 6413 4812 6427 4826
rect 6453 4812 6467 4826
rect 6393 4753 6407 4767
rect 6373 4633 6387 4647
rect 6393 4613 6407 4627
rect 6373 4593 6387 4607
rect 6373 4512 6387 4526
rect 6353 4393 6367 4407
rect 6533 4793 6547 4807
rect 6513 4713 6527 4727
rect 6473 4693 6487 4707
rect 6413 4593 6427 4607
rect 6513 4593 6527 4607
rect 6473 4554 6487 4568
rect 6573 5633 6587 5647
rect 6653 5933 6667 5947
rect 6693 5894 6707 5908
rect 6753 6113 6767 6127
rect 6753 6072 6767 6086
rect 6933 6372 6947 6386
rect 6873 6333 6887 6347
rect 6913 6333 6927 6347
rect 6913 6233 6927 6247
rect 7013 6372 7027 6386
rect 6972 6293 6986 6307
rect 6993 6293 7007 6307
rect 6953 6253 6967 6267
rect 6913 6173 6927 6187
rect 6793 6153 6807 6167
rect 6873 6153 6887 6167
rect 6773 6013 6787 6027
rect 6753 5953 6767 5967
rect 6673 5852 6687 5866
rect 6773 5894 6787 5908
rect 6753 5852 6767 5866
rect 6633 5813 6647 5827
rect 6713 5813 6727 5827
rect 6693 5733 6707 5747
rect 6613 5653 6627 5667
rect 6613 5594 6627 5608
rect 6673 5594 6687 5608
rect 6593 5533 6607 5547
rect 6653 5513 6667 5527
rect 6633 5374 6647 5388
rect 6573 5193 6587 5207
rect 6573 5153 6587 5167
rect 6573 5033 6587 5047
rect 6573 4854 6587 4868
rect 6573 4813 6587 4827
rect 6553 4733 6567 4747
rect 6553 4673 6567 4687
rect 6553 4613 6567 4627
rect 6533 4413 6547 4427
rect 6513 4393 6527 4407
rect 6493 4353 6507 4367
rect 6333 4292 6347 4306
rect 6353 4213 6367 4227
rect 6413 4213 6427 4227
rect 6413 4153 6427 4167
rect 6493 4153 6507 4167
rect 6353 3992 6367 4006
rect 6393 3992 6407 4006
rect 6433 3933 6447 3947
rect 6353 3853 6367 3867
rect 6393 3814 6407 3828
rect 6473 3814 6487 3828
rect 6373 3772 6387 3786
rect 6413 3772 6427 3786
rect 6473 3773 6487 3787
rect 6453 3653 6467 3667
rect 6373 3613 6387 3627
rect 6353 3493 6367 3507
rect 6313 3433 6327 3447
rect 6313 3412 6327 3426
rect 6433 3533 6447 3547
rect 6453 3513 6467 3527
rect 6473 3492 6487 3506
rect 6373 3393 6387 3407
rect 6613 5332 6627 5346
rect 6733 5594 6747 5608
rect 6713 5313 6727 5327
rect 6773 5793 6787 5807
rect 6913 6134 6927 6148
rect 6953 6133 6967 6147
rect 6813 6113 6827 6127
rect 6893 6113 6907 6127
rect 6873 6072 6887 6086
rect 6913 6072 6927 6086
rect 7053 6273 7067 6287
rect 7033 6253 7047 6267
rect 7013 6114 7027 6128
rect 6973 6093 6987 6107
rect 6873 6013 6887 6027
rect 6953 6013 6967 6027
rect 6813 5993 6827 6007
rect 6933 5993 6947 6007
rect 6793 5733 6807 5747
rect 6793 5613 6807 5627
rect 6793 5552 6807 5566
rect 6873 5633 6887 5647
rect 6933 5633 6947 5647
rect 6853 5613 6867 5627
rect 6973 5893 6987 5907
rect 7013 6073 7027 6087
rect 7053 6233 7067 6247
rect 7033 5953 7047 5967
rect 7093 6934 7107 6948
rect 7093 6853 7107 6867
rect 7093 6573 7107 6587
rect 7133 6934 7147 6948
rect 7113 6513 7127 6527
rect 7133 6493 7147 6507
rect 7133 6472 7147 6486
rect 7273 7373 7287 7387
rect 7193 7233 7207 7247
rect 7253 7233 7267 7247
rect 7213 7073 7227 7087
rect 7233 7053 7247 7067
rect 7213 7013 7227 7027
rect 7273 7033 7287 7047
rect 7453 7933 7467 7947
rect 7493 7913 7507 7927
rect 7433 7833 7447 7847
rect 7393 7733 7407 7747
rect 7493 7833 7507 7847
rect 7473 7813 7487 7827
rect 7393 7674 7407 7688
rect 7433 7673 7447 7687
rect 7313 7553 7327 7567
rect 7313 7493 7327 7507
rect 7293 6953 7307 6967
rect 7153 6453 7167 6467
rect 7133 6173 7147 6187
rect 7093 6114 7107 6128
rect 7273 6934 7287 6948
rect 7253 6892 7267 6906
rect 7213 6833 7227 6847
rect 7253 6833 7267 6847
rect 7213 6633 7227 6647
rect 7373 7573 7387 7587
rect 7413 7513 7427 7527
rect 7393 7473 7407 7487
rect 7373 7453 7387 7467
rect 7353 7373 7367 7387
rect 7373 7273 7387 7287
rect 7473 7673 7487 7687
rect 7453 7613 7467 7627
rect 7493 7573 7507 7587
rect 7473 7513 7487 7527
rect 7433 7473 7447 7487
rect 7413 7453 7427 7467
rect 7453 7454 7467 7468
rect 7433 7412 7447 7426
rect 7453 7393 7467 7407
rect 7453 7333 7467 7347
rect 7493 7373 7507 7387
rect 7473 7233 7487 7247
rect 7393 7193 7407 7207
rect 7453 7193 7467 7207
rect 7433 7154 7447 7168
rect 7473 7154 7487 7168
rect 7333 7112 7347 7126
rect 7453 7112 7467 7126
rect 7373 7073 7387 7087
rect 7433 7073 7447 7087
rect 7433 7033 7447 7047
rect 7753 8073 7767 8087
rect 7793 8073 7807 8087
rect 7593 8053 7607 8067
rect 7733 8053 7747 8067
rect 7573 8033 7587 8047
rect 7633 8013 7647 8027
rect 7713 8013 7727 8027
rect 7613 7932 7627 7946
rect 7653 7913 7667 7927
rect 7553 7873 7567 7887
rect 7693 7713 7707 7727
rect 7593 7674 7607 7688
rect 7673 7674 7687 7688
rect 7553 7573 7567 7587
rect 7533 7493 7547 7507
rect 7513 7333 7527 7347
rect 7513 7293 7527 7307
rect 7513 7272 7527 7286
rect 7493 7093 7507 7107
rect 7473 7033 7487 7047
rect 7373 7013 7387 7027
rect 7453 7013 7467 7027
rect 7353 6993 7367 7007
rect 7333 6934 7347 6948
rect 7593 7613 7607 7627
rect 7573 7533 7587 7547
rect 7573 7493 7587 7507
rect 7573 7373 7587 7387
rect 7573 7313 7587 7327
rect 7673 7593 7687 7607
rect 7713 7573 7727 7587
rect 7693 7533 7707 7547
rect 7613 7453 7627 7467
rect 7653 7454 7667 7468
rect 7773 7974 7787 7988
rect 7773 7893 7787 7907
rect 7933 8333 7947 8347
rect 7893 8313 7907 8327
rect 7873 8073 7887 8087
rect 7833 8053 7847 8067
rect 8153 8432 8167 8446
rect 8133 8393 8147 8407
rect 7933 8172 7947 8186
rect 7933 8133 7947 8147
rect 7893 8013 7907 8027
rect 7853 7974 7867 7988
rect 8193 8293 8207 8307
rect 8133 8273 8147 8287
rect 8153 8194 8167 8208
rect 8093 8172 8107 8186
rect 7973 8133 7987 8147
rect 8313 8873 8327 8887
rect 8333 8753 8347 8767
rect 8373 8753 8387 8767
rect 8312 8733 8326 8747
rect 8333 8734 8347 8748
rect 8293 8692 8307 8706
rect 8293 8633 8307 8647
rect 8253 8433 8267 8447
rect 8273 8353 8287 8367
rect 8133 8152 8147 8166
rect 8173 8093 8187 8107
rect 8093 8073 8107 8087
rect 7953 8033 7967 8047
rect 8193 8033 8207 8047
rect 8253 8033 8267 8047
rect 7833 7932 7847 7946
rect 7873 7893 7887 7907
rect 7793 7733 7807 7747
rect 7793 7674 7807 7688
rect 7833 7674 7847 7688
rect 7893 7873 7907 7887
rect 8073 7813 8087 7827
rect 8053 7753 8067 7767
rect 7913 7674 7927 7688
rect 8013 7674 8027 7688
rect 8133 7753 8147 7767
rect 8113 7733 8127 7747
rect 8093 7674 8107 7688
rect 7813 7632 7827 7646
rect 7873 7633 7887 7647
rect 7893 7613 7907 7627
rect 8053 7613 8067 7627
rect 7913 7553 7927 7567
rect 8073 7553 8087 7567
rect 7893 7533 7907 7547
rect 8053 7533 8067 7547
rect 7753 7473 7767 7487
rect 7813 7473 7827 7487
rect 7733 7453 7747 7467
rect 7593 7253 7607 7267
rect 7793 7434 7807 7448
rect 7673 7412 7687 7426
rect 7733 7393 7747 7407
rect 7753 7373 7767 7387
rect 7773 7253 7787 7267
rect 7713 7233 7727 7247
rect 7593 7173 7607 7187
rect 7533 7113 7547 7127
rect 7573 7113 7587 7127
rect 7513 7013 7527 7027
rect 7473 6973 7487 6987
rect 7453 6934 7467 6948
rect 7493 6934 7507 6948
rect 7553 6933 7567 6947
rect 7433 6893 7447 6907
rect 7333 6853 7347 6867
rect 7433 6853 7447 6867
rect 7413 6773 7427 6787
rect 7353 6713 7367 6727
rect 7333 6612 7347 6626
rect 7192 6513 7206 6527
rect 7213 6513 7227 6527
rect 7173 6113 7187 6127
rect 7273 6573 7287 6587
rect 7553 6892 7567 6906
rect 7573 6793 7587 6807
rect 7473 6733 7487 6747
rect 7713 7112 7727 7126
rect 7633 7073 7647 7087
rect 7593 6693 7607 6707
rect 7453 6633 7467 6647
rect 7433 6613 7447 6627
rect 7653 6953 7667 6967
rect 7633 6673 7647 6687
rect 7713 6993 7727 7007
rect 7753 7073 7767 7087
rect 7733 6953 7747 6967
rect 7913 7432 7927 7446
rect 7793 7112 7807 7126
rect 8013 7113 8027 7127
rect 7793 7073 7807 7087
rect 7793 6993 7807 7007
rect 7773 6953 7787 6967
rect 7693 6892 7707 6906
rect 7733 6853 7747 6867
rect 7733 6793 7747 6807
rect 7713 6673 7727 6687
rect 7653 6612 7667 6626
rect 7693 6612 7707 6626
rect 7593 6593 7607 6607
rect 7633 6593 7647 6607
rect 7353 6513 7367 6527
rect 7473 6513 7487 6527
rect 7513 6513 7527 6527
rect 7593 6513 7607 6527
rect 7233 6353 7247 6367
rect 7213 6233 7227 6247
rect 7233 6193 7247 6207
rect 7213 6113 7227 6127
rect 7093 5973 7107 5987
rect 7013 5933 7027 5947
rect 7053 5933 7067 5947
rect 6993 5852 7007 5866
rect 6973 5833 6987 5847
rect 6813 5513 6827 5527
rect 6893 5552 6907 5566
rect 6953 5513 6967 5527
rect 6853 5493 6867 5507
rect 6773 5473 6787 5487
rect 6813 5473 6827 5487
rect 6793 5433 6807 5447
rect 6773 5373 6787 5387
rect 6773 5332 6787 5346
rect 6733 5293 6747 5307
rect 6753 5273 6767 5287
rect 6773 5253 6787 5267
rect 6973 5413 6987 5427
rect 6853 5374 6867 5388
rect 6893 5374 6907 5388
rect 6933 5374 6947 5388
rect 6953 5353 6967 5367
rect 6833 5332 6847 5346
rect 6813 5253 6827 5267
rect 6653 5193 6667 5207
rect 6753 5232 6767 5246
rect 6753 5173 6767 5187
rect 6633 5113 6647 5127
rect 6793 5193 6807 5207
rect 6853 5273 6867 5287
rect 6833 5113 6847 5127
rect 6733 5074 6747 5088
rect 6813 5053 6827 5067
rect 6653 5033 6667 5047
rect 6693 4993 6707 5007
rect 6633 4953 6647 4967
rect 6653 4854 6667 4868
rect 6753 5032 6767 5046
rect 6713 4953 6727 4967
rect 6693 4733 6707 4747
rect 6673 4673 6687 4687
rect 6633 4533 6647 4547
rect 6593 4393 6607 4407
rect 6553 4373 6567 4387
rect 6593 4372 6607 4386
rect 6532 4334 6546 4348
rect 6553 4334 6567 4348
rect 6633 4334 6647 4348
rect 6613 4292 6627 4306
rect 6653 4292 6667 4306
rect 6633 4253 6647 4267
rect 6613 4233 6627 4247
rect 6633 4213 6647 4227
rect 6613 4173 6627 4187
rect 6653 4173 6667 4187
rect 6613 4133 6627 4147
rect 6713 4633 6727 4647
rect 6793 5013 6807 5027
rect 6793 4913 6807 4927
rect 6813 4893 6827 4907
rect 6793 4633 6807 4647
rect 6733 4613 6747 4627
rect 6733 4493 6747 4507
rect 6753 4333 6767 4347
rect 6733 4293 6747 4307
rect 6713 4153 6727 4167
rect 6693 4093 6707 4107
rect 6653 4033 6667 4047
rect 6633 3992 6647 4006
rect 6653 3933 6667 3947
rect 6693 3933 6707 3947
rect 6613 3853 6627 3867
rect 6653 3814 6667 3828
rect 6593 3772 6607 3786
rect 6633 3733 6647 3747
rect 6753 4193 6767 4207
rect 6773 4093 6787 4107
rect 6753 3953 6767 3967
rect 6933 5333 6947 5347
rect 6873 5253 6887 5267
rect 6993 5393 7007 5407
rect 6973 5233 6987 5247
rect 6953 5213 6967 5227
rect 6913 5193 6927 5207
rect 7053 5894 7067 5908
rect 7193 6072 7207 6086
rect 7153 6013 7167 6027
rect 7173 5953 7187 5967
rect 7113 5913 7127 5927
rect 7153 5913 7167 5927
rect 7073 5852 7087 5866
rect 7113 5852 7127 5866
rect 7133 5733 7147 5747
rect 7033 5613 7047 5627
rect 7013 5253 7027 5267
rect 7053 5594 7067 5608
rect 7093 5594 7107 5608
rect 7193 5894 7207 5908
rect 7173 5852 7187 5866
rect 7193 5833 7207 5847
rect 7193 5713 7207 5727
rect 7153 5613 7167 5627
rect 7053 5493 7067 5507
rect 7073 5473 7087 5487
rect 7153 5513 7167 5527
rect 7093 5332 7107 5346
rect 7093 5293 7107 5307
rect 7033 5193 7047 5207
rect 6993 5173 7007 5187
rect 6953 5133 6967 5147
rect 6933 5113 6947 5127
rect 6933 5053 6947 5067
rect 6893 4933 6907 4947
rect 7013 4893 7027 4907
rect 6933 4854 6947 4868
rect 6993 4854 7007 4868
rect 6873 4812 6887 4826
rect 6913 4812 6927 4826
rect 6853 4493 6867 4507
rect 7013 4813 7027 4827
rect 6993 4753 7007 4767
rect 7013 4673 7027 4687
rect 6953 4593 6967 4607
rect 6893 4533 6907 4547
rect 6873 4373 6887 4387
rect 6973 4512 6987 4526
rect 6893 4353 6907 4367
rect 6933 4473 6947 4487
rect 6973 4273 6987 4287
rect 7033 4553 7047 4567
rect 7133 5113 7147 5127
rect 7113 5053 7127 5067
rect 7133 5013 7147 5027
rect 7173 5253 7187 5267
rect 7173 5093 7187 5107
rect 7193 5052 7207 5066
rect 7113 4973 7127 4987
rect 7153 4993 7167 5007
rect 7133 4933 7147 4947
rect 7272 6453 7286 6467
rect 7293 6453 7307 6467
rect 7253 5933 7267 5947
rect 7433 6473 7447 6487
rect 7373 6453 7387 6467
rect 7353 6433 7367 6447
rect 7333 6414 7347 6428
rect 7353 6372 7367 6386
rect 7293 6333 7307 6347
rect 7493 6493 7507 6507
rect 7473 6373 7487 6387
rect 7393 6333 7407 6347
rect 7433 6333 7447 6347
rect 7353 6293 7367 6307
rect 7553 6453 7567 6467
rect 7513 6433 7527 6447
rect 7533 6414 7547 6428
rect 7513 6393 7527 6407
rect 7513 6293 7527 6307
rect 7493 6253 7507 6267
rect 7533 6253 7547 6267
rect 7393 6233 7407 6247
rect 7353 6153 7367 6167
rect 7692 6393 7706 6407
rect 7713 6394 7727 6408
rect 7573 6372 7587 6386
rect 7553 6193 7567 6207
rect 7553 6153 7567 6167
rect 7433 6114 7447 6128
rect 7493 6114 7507 6128
rect 7293 6093 7307 6107
rect 7333 6072 7347 6086
rect 7293 6033 7307 6047
rect 7413 6073 7427 6087
rect 7513 6073 7527 6087
rect 7372 6033 7386 6047
rect 7393 6033 7407 6047
rect 7333 5993 7347 6007
rect 7353 5953 7367 5967
rect 7313 5894 7327 5908
rect 7373 5894 7387 5908
rect 7253 5853 7267 5867
rect 7293 5852 7307 5866
rect 7273 5773 7287 5787
rect 7253 5653 7267 5667
rect 7353 5733 7367 5747
rect 7333 5713 7347 5727
rect 7293 5613 7307 5627
rect 7273 5573 7287 5587
rect 7393 5653 7407 5667
rect 7513 6033 7527 6047
rect 7673 6333 7687 6347
rect 7653 6233 7667 6247
rect 7613 6072 7627 6086
rect 7633 6013 7647 6027
rect 7493 5933 7507 5947
rect 7553 5894 7567 5908
rect 7513 5852 7527 5866
rect 7633 5933 7647 5947
rect 7613 5893 7627 5907
rect 7633 5853 7647 5867
rect 7613 5773 7627 5787
rect 7633 5753 7647 5767
rect 7573 5733 7587 5747
rect 7612 5713 7626 5727
rect 7633 5713 7647 5727
rect 7433 5613 7447 5627
rect 7493 5613 7507 5627
rect 7533 5653 7547 5667
rect 7513 5593 7527 5607
rect 7293 5393 7307 5407
rect 7333 5552 7347 5566
rect 7413 5553 7427 5567
rect 7373 5493 7387 5507
rect 7233 5273 7247 5287
rect 7293 5253 7307 5267
rect 7313 5233 7327 5247
rect 7353 5233 7367 5247
rect 7233 5193 7247 5207
rect 7633 5673 7647 5687
rect 7653 5653 7667 5667
rect 7553 5613 7567 5627
rect 7613 5613 7627 5627
rect 7653 5613 7667 5627
rect 7613 5552 7627 5566
rect 7553 5493 7567 5507
rect 7453 5453 7467 5467
rect 7353 5193 7367 5207
rect 7413 5193 7427 5207
rect 7313 5133 7327 5147
rect 7293 5113 7307 5127
rect 7253 4993 7267 5007
rect 7273 4933 7287 4947
rect 7233 4892 7247 4906
rect 7153 4873 7167 4887
rect 7213 4873 7227 4887
rect 7273 4854 7287 4868
rect 7113 4833 7127 4847
rect 7253 4834 7267 4848
rect 7193 4812 7207 4826
rect 7233 4713 7247 4727
rect 7133 4633 7147 4647
rect 7113 4554 7127 4568
rect 7153 4554 7167 4568
rect 7193 4554 7207 4568
rect 7233 4554 7247 4568
rect 7313 5013 7327 5027
rect 7333 4973 7347 4987
rect 7313 4933 7327 4947
rect 7473 5393 7487 5407
rect 7513 5374 7527 5388
rect 7653 5453 7667 5467
rect 7693 6153 7707 6167
rect 7693 6072 7707 6086
rect 7693 6013 7707 6027
rect 7793 6553 7807 6567
rect 7833 7093 7847 7107
rect 7933 7073 7947 7087
rect 7893 7013 7907 7027
rect 7953 6973 7967 6987
rect 7993 6953 8007 6967
rect 8033 6953 8047 6967
rect 7993 6873 8007 6887
rect 8033 6873 8047 6887
rect 7973 6853 7987 6867
rect 7933 6773 7947 6787
rect 7933 6634 7947 6648
rect 7973 6634 7987 6648
rect 7833 6513 7847 6527
rect 8013 6593 8027 6607
rect 7813 6493 7827 6507
rect 7913 6493 7927 6507
rect 7973 6393 7987 6407
rect 8033 6513 8047 6527
rect 7833 6373 7847 6387
rect 7753 6253 7767 6267
rect 7913 6253 7927 6267
rect 7733 6193 7747 6207
rect 7893 6193 7907 6207
rect 7853 6153 7867 6167
rect 7773 6114 7787 6128
rect 7813 6114 7827 6128
rect 7853 6114 7867 6128
rect 7753 6073 7767 6087
rect 7733 6053 7747 6067
rect 7753 5973 7767 5987
rect 7833 6013 7847 6027
rect 7833 5992 7847 6006
rect 7813 5953 7827 5967
rect 7793 5894 7807 5908
rect 7693 5852 7707 5866
rect 7733 5852 7747 5866
rect 7773 5833 7787 5847
rect 7853 5894 7867 5908
rect 7833 5833 7847 5847
rect 7813 5813 7827 5827
rect 7853 5813 7867 5827
rect 7693 5753 7707 5767
rect 7813 5733 7827 5747
rect 7753 5633 7767 5647
rect 7733 5552 7747 5566
rect 7692 5433 7706 5447
rect 7713 5433 7727 5447
rect 7673 5393 7687 5407
rect 7693 5373 7707 5387
rect 7473 5353 7487 5367
rect 7613 5332 7627 5346
rect 7673 5332 7687 5346
rect 7713 5332 7727 5346
rect 7853 5713 7867 5727
rect 7853 5673 7867 5687
rect 7873 5633 7887 5647
rect 7853 5594 7867 5608
rect 7753 5533 7767 5547
rect 7793 5533 7807 5547
rect 7893 5513 7907 5527
rect 7993 6353 8007 6367
rect 7953 6153 7967 6167
rect 8093 7533 8107 7547
rect 8173 7613 8187 7627
rect 8133 7593 8147 7607
rect 8153 7553 8167 7567
rect 8113 7513 8127 7527
rect 8073 7433 8087 7447
rect 8113 7453 8127 7467
rect 8073 7393 8087 7407
rect 8113 7393 8127 7407
rect 8093 7373 8107 7387
rect 8073 7113 8087 7127
rect 8113 7333 8127 7347
rect 8233 8013 8247 8027
rect 8213 7913 8227 7927
rect 8333 8593 8347 8607
rect 8313 8573 8327 8587
rect 8333 8533 8347 8547
rect 8393 8734 8407 8748
rect 8413 8693 8427 8707
rect 8833 10054 8847 10068
rect 8693 10012 8707 10026
rect 8753 10012 8767 10026
rect 8653 9953 8667 9967
rect 9633 11113 9647 11127
rect 9393 11094 9407 11108
rect 9472 11093 9486 11107
rect 9493 11093 9507 11107
rect 9593 11094 9607 11108
rect 9773 11094 9787 11108
rect 9833 11094 9847 11108
rect 9873 11094 9887 11108
rect 10053 11094 10067 11108
rect 10293 11094 10307 11108
rect 9113 11033 9127 11047
rect 9153 10953 9167 10967
rect 9373 11052 9387 11066
rect 9353 11033 9367 11047
rect 9193 10873 9207 10887
rect 9273 10873 9287 10887
rect 9233 10833 9247 10847
rect 9193 10794 9207 10808
rect 9113 10752 9127 10766
rect 9173 10752 9187 10766
rect 9213 10752 9227 10766
rect 9273 10752 9287 10766
rect 9233 10613 9247 10627
rect 9393 10873 9407 10887
rect 9433 10833 9447 10847
rect 9413 10813 9427 10827
rect 9413 10752 9427 10766
rect 9493 11052 9507 11066
rect 9653 11052 9667 11066
rect 9693 11052 9707 11066
rect 9613 10933 9627 10947
rect 9653 10893 9667 10907
rect 9573 10794 9587 10808
rect 9613 10794 9627 10808
rect 9753 10813 9767 10827
rect 9693 10773 9707 10787
rect 9633 10752 9647 10766
rect 9573 10633 9587 10647
rect 9373 10613 9387 10627
rect 9413 10613 9427 10627
rect 9473 10613 9487 10627
rect 9053 10574 9067 10588
rect 9093 10574 9107 10588
rect 9273 10574 9287 10588
rect 9053 10453 9067 10467
rect 9033 10313 9047 10327
rect 8873 10274 8887 10288
rect 8993 10274 9007 10288
rect 9073 10293 9087 10307
rect 9373 10532 9387 10546
rect 9253 10473 9267 10487
rect 8973 10232 8987 10246
rect 9053 10232 9067 10246
rect 8933 10093 8947 10107
rect 8973 10093 8987 10107
rect 8893 10054 8907 10068
rect 8853 10012 8867 10026
rect 8833 9833 8847 9847
rect 8893 9793 8907 9807
rect 8713 9773 8727 9787
rect 8673 9754 8687 9768
rect 8792 9753 8806 9767
rect 8813 9754 8827 9768
rect 8853 9754 8867 9768
rect 8913 9773 8927 9787
rect 8653 9693 8667 9707
rect 8713 9693 8727 9707
rect 8793 9693 8807 9707
rect 8773 9593 8787 9607
rect 8673 9533 8687 9547
rect 8733 9534 8747 9548
rect 8653 9492 8667 9506
rect 8633 9293 8647 9307
rect 8753 9492 8767 9506
rect 8873 9712 8887 9726
rect 8913 9693 8927 9707
rect 9033 9754 9047 9768
rect 9033 9713 9047 9727
rect 9153 10232 9167 10246
rect 9193 10193 9207 10207
rect 9233 10153 9247 10167
rect 9333 10433 9347 10447
rect 9313 10313 9327 10327
rect 9453 10574 9467 10588
rect 9493 10574 9507 10588
rect 9693 10574 9707 10588
rect 9473 10532 9487 10546
rect 9713 10532 9727 10546
rect 9753 10533 9767 10547
rect 9493 10413 9507 10427
rect 9373 10313 9387 10327
rect 9413 10313 9427 10327
rect 9473 10313 9487 10327
rect 9433 10293 9447 10307
rect 9413 10273 9427 10287
rect 9253 10133 9267 10147
rect 9293 10133 9307 10147
rect 9233 10093 9247 10107
rect 9073 10073 9087 10087
rect 9173 10073 9187 10087
rect 9093 10053 9107 10067
rect 9133 10054 9147 10068
rect 9073 9933 9087 9947
rect 9153 10012 9167 10026
rect 9293 10013 9307 10027
rect 9393 10192 9407 10206
rect 9353 10054 9367 10068
rect 9433 10173 9447 10187
rect 9313 9993 9327 10007
rect 9373 9993 9387 10007
rect 9413 9933 9427 9947
rect 9113 9873 9127 9887
rect 9313 9754 9327 9768
rect 9353 9754 9367 9768
rect 9333 9712 9347 9726
rect 9013 9693 9027 9707
rect 9053 9693 9067 9707
rect 9093 9693 9107 9707
rect 9153 9693 9167 9707
rect 8933 9673 8947 9687
rect 8973 9673 8987 9687
rect 8913 9633 8927 9647
rect 8913 9492 8927 9506
rect 8793 9453 8807 9467
rect 8833 9453 8847 9467
rect 8613 9234 8627 9248
rect 8613 9192 8627 9206
rect 8553 9093 8567 9107
rect 8533 9033 8547 9047
rect 8973 9652 8987 9666
rect 9013 9573 9027 9587
rect 9073 9553 9087 9567
rect 9013 9534 9027 9548
rect 8993 9492 9007 9506
rect 9033 9453 9047 9467
rect 8933 9273 8947 9287
rect 9013 9273 9027 9287
rect 8773 9234 8787 9248
rect 8913 9234 8927 9248
rect 8973 9234 8987 9248
rect 9053 9253 9067 9267
rect 8673 9192 8687 9206
rect 9053 9213 9067 9227
rect 8913 9173 8927 9187
rect 8673 9133 8687 9147
rect 8713 9133 8727 9147
rect 8653 9073 8667 9087
rect 8653 9033 8667 9047
rect 8453 8994 8467 9008
rect 8613 8994 8627 9008
rect 8493 8972 8507 8986
rect 8573 8933 8587 8947
rect 8613 8913 8627 8927
rect 8533 8873 8547 8887
rect 8453 8813 8467 8827
rect 8473 8793 8487 8807
rect 8453 8713 8467 8727
rect 8433 8673 8447 8687
rect 8433 8513 8447 8527
rect 8413 8493 8427 8507
rect 8453 8493 8467 8507
rect 8433 8474 8447 8488
rect 8313 8453 8327 8467
rect 8353 8452 8367 8466
rect 8393 8452 8407 8466
rect 8293 8133 8307 8147
rect 8293 8013 8307 8027
rect 8273 7973 8287 7987
rect 8513 8714 8527 8728
rect 8553 8714 8567 8728
rect 8593 8714 8607 8728
rect 8493 8673 8507 8687
rect 8533 8672 8547 8686
rect 8593 8653 8607 8667
rect 8513 8613 8527 8627
rect 8693 9073 8707 9087
rect 8693 8993 8707 9007
rect 8733 9093 8747 9107
rect 8873 8993 8887 9007
rect 8853 8973 8867 8987
rect 8713 8913 8727 8927
rect 8693 8853 8707 8867
rect 8673 8833 8687 8847
rect 8713 8833 8727 8847
rect 8693 8793 8707 8807
rect 8733 8753 8747 8767
rect 8773 8733 8787 8747
rect 8613 8613 8627 8627
rect 8993 9192 9007 9206
rect 8993 9153 9007 9167
rect 8973 9033 8987 9047
rect 9273 9573 9287 9587
rect 9233 9553 9247 9567
rect 9413 9553 9427 9567
rect 9473 9553 9487 9567
rect 9253 9492 9267 9506
rect 9213 9473 9227 9487
rect 9113 9433 9127 9447
rect 9093 9133 9107 9147
rect 9073 9053 9087 9067
rect 9053 9013 9067 9027
rect 8993 8993 9007 9007
rect 9193 9293 9207 9307
rect 10373 11093 10387 11107
rect 10353 11073 10367 11087
rect 9853 11033 9867 11047
rect 10073 11052 10087 11066
rect 10273 11052 10287 11066
rect 10313 11052 10327 11066
rect 9893 10993 9907 11007
rect 10293 10933 10307 10947
rect 9793 10893 9807 10907
rect 10093 10853 10107 10867
rect 9933 10833 9947 10847
rect 9853 10813 9867 10827
rect 9893 10794 9907 10808
rect 10053 10794 10067 10808
rect 10373 11052 10387 11066
rect 10513 11094 10527 11108
rect 10633 11093 10647 11107
rect 10673 11094 10687 11108
rect 10713 11094 10727 11108
rect 10753 11094 10767 11108
rect 10453 11033 10467 11047
rect 10533 11033 10547 11047
rect 10633 11033 10647 11047
rect 10493 10973 10507 10987
rect 10353 10913 10367 10927
rect 10653 10973 10667 10987
rect 10533 10873 10547 10887
rect 10513 10853 10527 10867
rect 10333 10794 10347 10808
rect 10373 10794 10387 10808
rect 10553 10833 10567 10847
rect 10553 10794 10567 10808
rect 9873 10752 9887 10766
rect 9933 10753 9947 10767
rect 10073 10752 10087 10766
rect 10113 10752 10127 10766
rect 9793 10713 9807 10727
rect 9833 10713 9847 10727
rect 10073 10653 10087 10667
rect 10053 10613 10067 10627
rect 9853 10574 9867 10588
rect 9893 10574 9907 10588
rect 10033 10574 10047 10588
rect 9913 10532 9927 10546
rect 10033 10533 10047 10547
rect 10133 10574 10147 10588
rect 10373 10753 10387 10767
rect 10813 11093 10827 11107
rect 10973 11094 10987 11108
rect 11133 11094 11147 11108
rect 11173 11094 11187 11108
rect 10773 11033 10787 11047
rect 10693 10973 10707 10987
rect 10733 10973 10747 10987
rect 10673 10913 10687 10927
rect 10533 10752 10547 10766
rect 10653 10752 10667 10766
rect 10413 10613 10427 10627
rect 10533 10613 10547 10627
rect 10673 10613 10687 10627
rect 10093 10532 10107 10546
rect 10053 10493 10067 10507
rect 10153 10493 10167 10507
rect 9853 10473 9867 10487
rect 9833 10353 9847 10367
rect 9773 10313 9787 10327
rect 9593 10293 9607 10307
rect 9673 10193 9687 10207
rect 9793 10273 9807 10287
rect 9733 10133 9747 10147
rect 9773 10133 9787 10147
rect 9573 10093 9587 10107
rect 9513 10053 9527 10067
rect 9613 10073 9627 10087
rect 9673 10054 9687 10068
rect 9513 9973 9527 9987
rect 9533 9813 9547 9827
rect 9573 9793 9587 9807
rect 10353 10574 10367 10588
rect 10333 10532 10347 10546
rect 10493 10573 10507 10587
rect 10573 10574 10587 10588
rect 10633 10553 10647 10567
rect 10493 10532 10507 10546
rect 10373 10513 10387 10527
rect 10413 10513 10427 10527
rect 10593 10532 10607 10546
rect 10553 10493 10567 10507
rect 10593 10433 10607 10447
rect 10293 10413 10307 10427
rect 10513 10353 10527 10367
rect 10593 10353 10607 10367
rect 9893 10274 9907 10288
rect 10053 10274 10067 10288
rect 10113 10274 10127 10288
rect 9853 10232 9867 10246
rect 9833 10193 9847 10207
rect 10093 10232 10107 10246
rect 9913 10173 9927 10187
rect 10013 10173 10027 10187
rect 10053 10173 10067 10187
rect 9893 10133 9907 10147
rect 9793 10073 9807 10087
rect 9853 10054 9867 10068
rect 9953 10053 9967 10067
rect 9793 10012 9807 10026
rect 9833 10012 9847 10026
rect 9873 9973 9887 9987
rect 9773 9933 9787 9947
rect 9933 9813 9947 9827
rect 9653 9754 9667 9768
rect 9693 9754 9707 9768
rect 9753 9754 9767 9768
rect 9793 9754 9807 9768
rect 10033 10133 10047 10147
rect 10133 10133 10147 10147
rect 10013 10012 10027 10026
rect 10353 10274 10367 10288
rect 10353 10213 10367 10227
rect 10333 10173 10347 10187
rect 10133 10093 10147 10107
rect 10193 10093 10207 10107
rect 10093 10054 10107 10068
rect 10313 10054 10327 10068
rect 10553 10313 10567 10327
rect 10573 10232 10587 10246
rect 10953 11052 10967 11066
rect 10993 11052 11007 11066
rect 10813 10933 10827 10947
rect 10733 10873 10747 10887
rect 10753 10853 10767 10867
rect 11193 11052 11207 11066
rect 11133 10833 11147 10847
rect 10813 10794 10827 10808
rect 10893 10794 10907 10808
rect 10753 10752 10767 10766
rect 10953 10793 10967 10807
rect 11013 10794 11027 10808
rect 11073 10793 11087 10807
rect 11213 10794 11227 10808
rect 10893 10733 10907 10747
rect 10833 10693 10847 10707
rect 10833 10613 10847 10627
rect 10793 10574 10807 10588
rect 10693 10532 10707 10546
rect 10653 10393 10667 10407
rect 10633 10193 10647 10207
rect 10373 10093 10387 10107
rect 10513 10093 10527 10107
rect 10593 10093 10607 10107
rect 10433 10053 10447 10067
rect 10493 10054 10507 10068
rect 10553 10054 10567 10068
rect 10113 10012 10127 10026
rect 9953 9793 9967 9807
rect 9993 9754 10007 9768
rect 10073 9973 10087 9987
rect 10293 9973 10307 9987
rect 10073 9933 10087 9947
rect 9553 9712 9567 9726
rect 9693 9713 9707 9727
rect 9933 9713 9947 9727
rect 9973 9712 9987 9726
rect 10013 9712 10027 9726
rect 9773 9673 9787 9687
rect 9573 9573 9587 9587
rect 9953 9573 9967 9587
rect 9493 9534 9507 9548
rect 9413 9492 9427 9506
rect 9512 9492 9526 9506
rect 9533 9493 9547 9507
rect 9413 9293 9427 9307
rect 9453 9293 9467 9307
rect 9313 9253 9327 9267
rect 9233 9234 9247 9248
rect 9373 9234 9387 9248
rect 9413 9234 9427 9248
rect 9473 9192 9487 9206
rect 9213 9173 9227 9187
rect 9373 9173 9387 9187
rect 9433 9173 9447 9187
rect 9133 9113 9147 9127
rect 9413 9113 9427 9127
rect 9173 9053 9187 9067
rect 9133 9013 9147 9027
rect 9073 8994 9087 9008
rect 9113 8994 9127 9008
rect 8953 8933 8967 8947
rect 9053 8953 9067 8967
rect 9013 8913 9027 8927
rect 8933 8853 8947 8867
rect 9053 8853 9067 8867
rect 8913 8714 8927 8728
rect 8913 8673 8927 8687
rect 8793 8633 8807 8647
rect 8853 8633 8867 8647
rect 8873 8593 8887 8607
rect 8593 8573 8607 8587
rect 8753 8573 8767 8587
rect 8533 8553 8547 8567
rect 8512 8473 8526 8487
rect 8533 8473 8547 8487
rect 8673 8472 8687 8486
rect 8533 8452 8547 8466
rect 8493 8373 8507 8387
rect 8473 8333 8487 8347
rect 8333 8293 8347 8307
rect 8453 8253 8467 8267
rect 8393 8194 8407 8208
rect 8333 7933 8347 7947
rect 8313 7913 8327 7927
rect 8373 8152 8387 8166
rect 8413 8093 8427 8107
rect 8373 8073 8387 8087
rect 8373 7973 8387 7987
rect 8353 7873 8367 7887
rect 8333 7833 8347 7847
rect 8293 7773 8307 7787
rect 8273 7733 8287 7747
rect 8253 7713 8267 7727
rect 8313 7753 8327 7767
rect 8293 7713 8307 7727
rect 8233 7633 8247 7647
rect 8213 7373 8227 7387
rect 8273 7593 8287 7607
rect 8253 7353 8267 7367
rect 8193 7313 8207 7327
rect 8133 7273 8147 7287
rect 8173 7273 8187 7287
rect 8113 7093 8127 7107
rect 8173 7233 8187 7247
rect 8213 7154 8227 7168
rect 8193 7112 8207 7126
rect 8233 7113 8247 7127
rect 8173 7093 8187 7107
rect 8133 6993 8147 7007
rect 8213 6993 8227 7007
rect 8173 6973 8187 6987
rect 8253 7093 8267 7107
rect 8293 7513 8307 7527
rect 8293 7353 8307 7367
rect 8233 6933 8247 6947
rect 8193 6892 8207 6906
rect 8093 6733 8107 6747
rect 8293 6993 8307 7007
rect 8273 6973 8287 6987
rect 8153 6634 8167 6648
rect 8093 6573 8107 6587
rect 8073 6473 8087 6487
rect 8053 6453 8067 6467
rect 8213 6613 8227 6627
rect 8193 6573 8207 6587
rect 8133 6553 8147 6567
rect 8113 6533 8127 6547
rect 8173 6533 8187 6547
rect 8133 6473 8147 6487
rect 8113 6413 8127 6427
rect 8113 6373 8127 6387
rect 8093 6313 8107 6327
rect 8073 6293 8087 6307
rect 8033 6253 8047 6267
rect 8113 6153 8127 6167
rect 8033 6114 8047 6128
rect 8073 6114 8087 6128
rect 8093 6072 8107 6086
rect 8053 6053 8067 6067
rect 7993 5953 8007 5967
rect 8033 5953 8047 5967
rect 8073 5953 8087 5967
rect 7933 5893 7947 5907
rect 7993 5894 8007 5908
rect 8033 5894 8047 5908
rect 8093 5894 8107 5908
rect 8013 5852 8027 5866
rect 8073 5852 8087 5866
rect 8033 5813 8047 5827
rect 7952 5773 7966 5787
rect 7973 5773 7987 5787
rect 7933 5713 7947 5727
rect 7933 5594 7947 5608
rect 7933 5553 7947 5567
rect 7853 5493 7867 5507
rect 7913 5493 7927 5507
rect 7833 5433 7847 5447
rect 7833 5392 7847 5406
rect 7573 5273 7587 5287
rect 7693 5273 7707 5287
rect 7733 5273 7747 5287
rect 7613 5233 7627 5247
rect 7653 5233 7667 5247
rect 7533 5193 7547 5207
rect 7592 5193 7606 5207
rect 7613 5193 7627 5207
rect 7453 5173 7467 5187
rect 7593 5113 7607 5127
rect 7493 5073 7507 5087
rect 7613 5052 7627 5066
rect 7793 5233 7807 5247
rect 7713 5073 7727 5087
rect 7753 5053 7767 5067
rect 7713 4993 7727 5007
rect 7533 4933 7547 4947
rect 7573 4933 7587 4947
rect 7693 4933 7707 4947
rect 7793 4933 7807 4947
rect 7413 4893 7427 4907
rect 7513 4893 7527 4907
rect 7373 4854 7387 4868
rect 7473 4834 7487 4848
rect 7333 4812 7347 4826
rect 7393 4812 7407 4826
rect 7313 4713 7327 4727
rect 7293 4673 7307 4687
rect 7453 4713 7467 4727
rect 7433 4653 7447 4667
rect 7293 4633 7307 4647
rect 7273 4593 7287 4607
rect 7093 4513 7107 4527
rect 7173 4512 7187 4526
rect 7113 4453 7127 4467
rect 7213 4453 7227 4467
rect 7193 4373 7207 4387
rect 7093 4353 7107 4367
rect 7173 4353 7187 4367
rect 7133 4334 7147 4348
rect 7033 4293 7047 4307
rect 6993 4233 7007 4247
rect 6853 4153 6867 4167
rect 6953 4153 6967 4167
rect 6933 4093 6947 4107
rect 6833 3992 6847 4006
rect 6913 3993 6927 4007
rect 6993 4093 7007 4107
rect 7073 4273 7087 4287
rect 7053 4253 7067 4267
rect 7153 4193 7167 4207
rect 7193 4213 7207 4227
rect 7173 4133 7187 4147
rect 7113 4113 7127 4127
rect 7153 4113 7167 4127
rect 7033 4073 7047 4087
rect 6973 4034 6987 4048
rect 7053 4034 7067 4048
rect 6953 3992 6967 4006
rect 6873 3953 6887 3967
rect 6913 3953 6927 3967
rect 6773 3893 6787 3907
rect 6813 3893 6827 3907
rect 6793 3873 6807 3887
rect 6773 3853 6787 3867
rect 6833 3853 6847 3867
rect 6853 3772 6867 3786
rect 6793 3733 6807 3747
rect 6773 3673 6787 3687
rect 6753 3633 6767 3647
rect 6813 3633 6827 3647
rect 6733 3613 6747 3627
rect 6713 3533 6727 3547
rect 6513 3453 6527 3467
rect 6533 3393 6547 3407
rect 6413 3373 6427 3387
rect 6313 3353 6327 3367
rect 6713 3494 6727 3508
rect 6573 3453 6587 3467
rect 6553 3333 6567 3347
rect 6593 3393 6607 3407
rect 6793 3393 6807 3407
rect 6313 3273 6327 3287
rect 6153 3233 6167 3247
rect 6093 3173 6107 3187
rect 6113 2994 6127 3008
rect 5993 2953 6007 2967
rect 5973 2913 5987 2927
rect 6093 2873 6107 2887
rect 6113 2853 6127 2867
rect 6113 2813 6127 2827
rect 5973 2773 5987 2787
rect 6013 2774 6027 2788
rect 6073 2774 6087 2788
rect 6133 2773 6147 2787
rect 6073 2733 6087 2747
rect 6013 2713 6027 2727
rect 6053 2713 6067 2727
rect 5993 2693 6007 2707
rect 6073 2453 6087 2467
rect 5933 2373 5947 2387
rect 6013 2393 6027 2407
rect 5993 2333 6007 2347
rect 5893 2254 5907 2268
rect 5933 2254 5947 2268
rect 5993 2253 6007 2267
rect 5853 2193 5867 2207
rect 5873 2093 5887 2107
rect 5713 1853 5727 1867
rect 5753 1852 5767 1866
rect 5733 1773 5747 1787
rect 5753 1753 5767 1767
rect 5773 1734 5787 1748
rect 5853 1813 5867 1827
rect 5793 1692 5807 1706
rect 5693 1673 5707 1687
rect 5673 1533 5687 1547
rect 5673 1453 5687 1467
rect 5713 1453 5727 1467
rect 5613 1393 5627 1407
rect 5653 1392 5667 1406
rect 5693 1392 5707 1406
rect 5673 1273 5687 1287
rect 5633 1214 5647 1228
rect 5773 1433 5787 1447
rect 5773 1392 5787 1406
rect 5653 1172 5667 1186
rect 5753 1173 5767 1187
rect 5713 1113 5727 1127
rect 5572 993 5586 1007
rect 5593 993 5607 1007
rect 5613 993 5627 1007
rect 5593 914 5607 928
rect 5513 872 5527 886
rect 5393 753 5407 767
rect 5493 753 5507 767
rect 5353 593 5367 607
rect 5653 733 5667 747
rect 5413 713 5427 727
rect 5573 713 5587 727
rect 5633 713 5647 727
rect 5473 694 5487 708
rect 5513 694 5527 708
rect 5553 693 5567 707
rect 5413 652 5427 666
rect 5453 652 5467 666
rect 5493 613 5507 627
rect 5493 433 5507 447
rect 5573 673 5587 687
rect 5573 633 5587 647
rect 5553 413 5567 427
rect 5393 333 5407 347
rect 5473 333 5487 347
rect 5533 353 5547 367
rect 5813 1093 5827 1107
rect 5773 914 5787 928
rect 5893 1953 5907 1967
rect 5893 1912 5907 1926
rect 5953 2193 5967 2207
rect 5953 2013 5967 2027
rect 5933 1993 5947 2007
rect 5913 1893 5927 1907
rect 6033 2093 6047 2107
rect 6693 3373 6707 3387
rect 6613 3333 6627 3347
rect 6413 3253 6427 3267
rect 6553 3253 6567 3267
rect 6253 3232 6267 3246
rect 6313 3232 6327 3246
rect 6213 3193 6227 3207
rect 6173 3053 6187 3067
rect 6313 3033 6327 3047
rect 6273 2994 6287 3008
rect 6233 2952 6247 2966
rect 6293 2952 6307 2966
rect 6233 2893 6247 2907
rect 6273 2774 6287 2788
rect 6253 2732 6267 2746
rect 6313 2633 6327 2647
rect 6173 2533 6187 2547
rect 6273 2533 6287 2547
rect 6153 2393 6167 2407
rect 6233 2513 6247 2527
rect 6253 2432 6267 2446
rect 6213 2353 6227 2367
rect 6133 2293 6147 2307
rect 6173 2293 6187 2307
rect 6173 2254 6187 2268
rect 6213 2254 6227 2268
rect 6153 2212 6167 2226
rect 6213 2213 6227 2227
rect 6073 2053 6087 2067
rect 6153 2053 6167 2067
rect 6033 2033 6047 2047
rect 6013 2013 6027 2027
rect 6073 1993 6087 2007
rect 6113 1993 6127 2007
rect 5953 1873 5967 1887
rect 5873 1734 5887 1748
rect 5853 1692 5867 1706
rect 5933 1793 5947 1807
rect 5913 1753 5927 1767
rect 5893 1493 5907 1507
rect 6073 1954 6087 1968
rect 6013 1912 6027 1926
rect 6053 1912 6067 1926
rect 6093 1873 6107 1887
rect 6013 1813 6027 1827
rect 6053 1813 6067 1827
rect 5993 1793 6007 1807
rect 5973 1753 5987 1767
rect 6013 1773 6027 1787
rect 6013 1692 6027 1706
rect 6133 1773 6147 1787
rect 6093 1672 6107 1686
rect 5973 1633 5987 1647
rect 5892 1453 5906 1467
rect 5913 1453 5927 1467
rect 5953 1453 5967 1467
rect 5913 1392 5927 1406
rect 5893 1293 5907 1307
rect 5853 1093 5867 1107
rect 5953 1172 5967 1186
rect 5993 1613 6007 1627
rect 6033 1573 6047 1587
rect 5993 1493 6007 1507
rect 5993 1392 6007 1406
rect 5973 1073 5987 1087
rect 5933 1053 5947 1067
rect 5913 953 5927 967
rect 5793 733 5807 747
rect 5713 694 5727 708
rect 5773 694 5787 708
rect 5673 573 5687 587
rect 5753 633 5767 647
rect 5773 613 5787 627
rect 5693 533 5707 547
rect 5753 533 5767 547
rect 5693 394 5707 408
rect 5653 352 5667 366
rect 5713 352 5727 366
rect 5533 313 5547 327
rect 5513 253 5527 267
rect 5473 233 5487 247
rect 5493 132 5507 146
rect 5873 913 5887 927
rect 5973 993 5987 1007
rect 6093 1434 6107 1448
rect 6113 1392 6127 1406
rect 6133 1313 6147 1327
rect 6073 1293 6087 1307
rect 6093 1233 6107 1247
rect 6173 1993 6187 2007
rect 6273 2173 6287 2187
rect 6213 1953 6227 1967
rect 6313 2373 6327 2387
rect 6593 3073 6607 3087
rect 6533 2994 6547 3008
rect 6413 2913 6427 2927
rect 6533 2813 6547 2827
rect 6413 2774 6427 2788
rect 6493 2774 6507 2788
rect 6393 2633 6407 2647
rect 6473 2732 6487 2746
rect 6533 2733 6547 2747
rect 6473 2653 6487 2667
rect 6413 2613 6427 2627
rect 6353 2293 6367 2307
rect 6293 2053 6307 2067
rect 6173 1913 6187 1927
rect 6213 1912 6227 1926
rect 6253 1912 6267 1926
rect 6293 1912 6307 1926
rect 6533 2493 6547 2507
rect 6433 2413 6447 2427
rect 6413 2053 6427 2067
rect 6373 1912 6387 1926
rect 6593 2433 6607 2447
rect 6713 3293 6727 3307
rect 6713 3253 6727 3267
rect 6693 3173 6707 3187
rect 6733 3033 6747 3047
rect 6633 2993 6647 3007
rect 6633 2952 6647 2966
rect 6713 2952 6727 2966
rect 6713 2913 6727 2927
rect 6753 2913 6767 2927
rect 6633 2774 6647 2788
rect 6673 2774 6687 2788
rect 6693 2732 6707 2746
rect 6733 2593 6747 2607
rect 6633 2533 6647 2547
rect 6713 2533 6727 2547
rect 6773 2513 6787 2527
rect 6873 3573 6887 3587
rect 6833 3492 6847 3506
rect 6873 3413 6887 3427
rect 6933 3533 6947 3547
rect 6913 3373 6927 3387
rect 6873 3353 6887 3367
rect 6813 3313 6827 3327
rect 6833 2813 6847 2827
rect 6873 3253 6887 3267
rect 6853 2732 6867 2746
rect 7073 3992 7087 4006
rect 7113 3992 7127 4006
rect 7033 3953 7047 3967
rect 7133 3873 7147 3887
rect 6993 3814 7007 3828
rect 7033 3814 7047 3828
rect 7073 3814 7087 3828
rect 7113 3814 7127 3828
rect 7133 3793 7147 3807
rect 7113 3773 7127 3787
rect 7173 4073 7187 4087
rect 6993 3753 7007 3767
rect 7133 3713 7147 3727
rect 7213 3993 7227 4007
rect 7273 4513 7287 4527
rect 7413 4593 7427 4607
rect 7373 4554 7387 4568
rect 7333 4493 7347 4507
rect 7433 4513 7447 4527
rect 7353 4453 7367 4467
rect 7393 4453 7407 4467
rect 7333 4393 7347 4407
rect 7393 4334 7407 4348
rect 7473 4673 7487 4687
rect 7352 4293 7366 4307
rect 7293 4213 7307 4227
rect 7273 4153 7287 4167
rect 7373 4292 7387 4306
rect 7433 4293 7447 4307
rect 7393 4273 7407 4287
rect 7373 4253 7387 4267
rect 7353 4133 7367 4147
rect 7313 3992 7327 4006
rect 7373 3993 7387 4007
rect 7273 3913 7287 3927
rect 7353 3913 7367 3927
rect 7253 3853 7267 3867
rect 7333 3873 7347 3887
rect 7393 3813 7407 3827
rect 7333 3793 7347 3807
rect 7233 3753 7247 3767
rect 6993 3673 7007 3687
rect 6973 3253 6987 3267
rect 6933 3153 6947 3167
rect 7073 3653 7087 3667
rect 7013 3573 7027 3587
rect 7173 3613 7187 3627
rect 7113 3514 7127 3528
rect 7153 3514 7167 3528
rect 7033 3493 7047 3507
rect 7033 3453 7047 3467
rect 7093 3453 7107 3467
rect 7153 3453 7167 3467
rect 7033 3393 7047 3407
rect 7033 3313 7047 3327
rect 7073 3294 7087 3308
rect 7133 3293 7147 3307
rect 7093 3252 7107 3266
rect 7133 3252 7147 3266
rect 7053 3213 7067 3227
rect 7073 3153 7087 3167
rect 6913 3033 6927 3047
rect 6993 3033 7007 3047
rect 6993 2913 7007 2927
rect 6933 2833 6947 2847
rect 7013 2753 7027 2767
rect 6953 2732 6967 2746
rect 6993 2732 7007 2746
rect 6873 2653 6887 2667
rect 7053 2673 7067 2687
rect 7153 3133 7167 3147
rect 7173 3073 7187 3087
rect 7213 3333 7227 3347
rect 7293 3713 7307 3727
rect 7333 3693 7347 3707
rect 7253 3553 7267 3567
rect 7293 3514 7307 3528
rect 7393 3653 7407 3667
rect 7353 3472 7367 3486
rect 7313 3393 7327 3407
rect 7353 3333 7367 3347
rect 7373 3313 7387 3327
rect 7313 3294 7327 3308
rect 7333 3252 7347 3266
rect 7293 3233 7307 3247
rect 7373 3233 7387 3247
rect 7233 3133 7247 3147
rect 7273 3133 7287 3147
rect 7253 2933 7267 2947
rect 7233 2853 7247 2867
rect 7013 2613 7027 2627
rect 7073 2613 7087 2627
rect 7053 2593 7067 2607
rect 6753 2494 6767 2508
rect 6913 2493 6927 2507
rect 6673 2413 6687 2427
rect 6813 2452 6827 2466
rect 6793 2333 6807 2347
rect 6893 2333 6907 2347
rect 7013 2333 7027 2347
rect 6633 2313 6647 2327
rect 6613 2293 6627 2307
rect 6493 2253 6507 2267
rect 6533 2253 6547 2267
rect 6473 2133 6487 2147
rect 6653 2273 6667 2287
rect 6553 2212 6567 2226
rect 6653 2213 6667 2227
rect 6593 2133 6607 2147
rect 6493 2073 6507 2087
rect 6613 2073 6627 2087
rect 6553 2053 6567 2067
rect 6453 2033 6467 2047
rect 6473 1993 6487 2007
rect 6513 1954 6527 1968
rect 6573 1954 6587 1968
rect 6433 1853 6447 1867
rect 6213 1813 6227 1827
rect 6333 1813 6347 1827
rect 6493 1813 6507 1827
rect 6293 1712 6307 1726
rect 6473 1712 6487 1726
rect 6453 1672 6467 1686
rect 6333 1493 6347 1507
rect 6293 1473 6307 1487
rect 6293 1434 6307 1448
rect 6473 1493 6487 1507
rect 6453 1473 6467 1487
rect 6313 1392 6327 1406
rect 6353 1392 6367 1406
rect 6433 1393 6447 1407
rect 6293 1293 6307 1307
rect 6193 1273 6207 1287
rect 6113 1172 6127 1186
rect 6093 1133 6107 1147
rect 6053 1033 6067 1047
rect 6033 953 6047 967
rect 6013 914 6027 928
rect 6133 1113 6147 1127
rect 6153 1093 6167 1107
rect 6133 1073 6147 1087
rect 6113 973 6127 987
rect 6093 893 6107 907
rect 5993 872 6007 886
rect 6033 872 6047 886
rect 5933 813 5947 827
rect 5953 713 5967 727
rect 6113 773 6127 787
rect 6213 1253 6227 1267
rect 6253 1153 6267 1167
rect 6213 1133 6227 1147
rect 6273 933 6287 947
rect 6253 914 6267 928
rect 6353 1233 6367 1247
rect 6333 1093 6347 1107
rect 6333 1053 6347 1067
rect 6373 933 6387 947
rect 6353 914 6367 928
rect 6193 872 6207 886
rect 6133 733 6147 747
rect 6213 813 6227 827
rect 6273 872 6287 886
rect 6313 853 6327 867
rect 6233 793 6247 807
rect 6313 793 6327 807
rect 6273 733 6287 747
rect 6033 673 6047 687
rect 5933 652 5947 666
rect 5993 653 6007 667
rect 5973 633 5987 647
rect 6013 633 6027 647
rect 5853 433 5867 447
rect 5953 433 5967 447
rect 5913 394 5927 408
rect 5993 394 6007 408
rect 5993 353 6007 367
rect 5933 313 5947 327
rect 5953 293 5967 307
rect 5893 253 5907 267
rect 5893 193 5907 207
rect 5693 174 5707 188
rect 5753 174 5767 188
rect 5853 174 5867 188
rect 5893 174 5907 188
rect 6193 652 6207 666
rect 6233 652 6247 666
rect 6273 652 6287 666
rect 6212 613 6226 627
rect 6233 613 6247 627
rect 6273 313 6287 327
rect 6133 193 6147 207
rect 6153 173 6167 187
rect 6353 733 6367 747
rect 6473 1273 6487 1287
rect 6473 1214 6487 1228
rect 6473 1093 6487 1107
rect 6513 1633 6527 1647
rect 6593 1913 6607 1927
rect 6553 1873 6567 1887
rect 6573 1733 6587 1747
rect 6553 1693 6567 1707
rect 6573 1593 6587 1607
rect 6533 1513 6547 1527
rect 6593 1293 6607 1307
rect 6733 2033 6747 2047
rect 6773 2133 6787 2147
rect 6753 1973 6767 1987
rect 6953 2293 6967 2307
rect 6933 2253 6947 2267
rect 6953 2234 6967 2248
rect 6993 2234 7007 2248
rect 6953 2133 6967 2147
rect 6913 2053 6927 2067
rect 6813 2033 6827 2047
rect 6673 1912 6687 1926
rect 6713 1912 6727 1926
rect 6753 1912 6767 1926
rect 6653 1773 6667 1787
rect 6893 2013 6907 2027
rect 6833 1973 6847 1987
rect 6873 1954 6887 1968
rect 6873 1913 6887 1927
rect 6833 1833 6847 1847
rect 6693 1753 6707 1767
rect 6813 1753 6827 1767
rect 7013 2013 7027 2027
rect 6993 1973 7007 1987
rect 6953 1954 6967 1968
rect 6913 1873 6927 1887
rect 6973 1833 6987 1847
rect 7013 1753 7027 1767
rect 6633 1693 6647 1707
rect 6673 1633 6687 1647
rect 6753 1533 6767 1547
rect 6913 1633 6927 1647
rect 6913 1612 6927 1626
rect 6793 1453 6807 1467
rect 6853 1453 6867 1467
rect 6893 1453 6907 1467
rect 6733 1392 6747 1406
rect 6813 1373 6827 1387
rect 6933 1553 6947 1567
rect 6773 1353 6787 1367
rect 6853 1353 6867 1367
rect 6633 1293 6647 1307
rect 6773 1293 6787 1307
rect 6533 1214 6547 1228
rect 6573 1214 6587 1228
rect 6613 1214 6627 1228
rect 6553 1153 6567 1167
rect 6653 1213 6667 1227
rect 6653 1173 6667 1187
rect 6793 1172 6807 1186
rect 6833 1172 6847 1186
rect 6753 1133 6767 1147
rect 6613 1073 6627 1087
rect 6613 973 6627 987
rect 6533 914 6547 928
rect 6593 914 6607 928
rect 6433 872 6447 886
rect 6473 872 6487 886
rect 6553 853 6567 867
rect 6553 793 6567 807
rect 6753 953 6767 967
rect 6793 914 6807 928
rect 6693 853 6707 867
rect 6613 793 6627 807
rect 6553 753 6567 767
rect 6593 753 6607 767
rect 6693 753 6707 767
rect 6433 694 6447 708
rect 6513 694 6527 708
rect 6373 652 6387 666
rect 6313 253 6327 267
rect 6413 394 6427 408
rect 6473 394 6487 408
rect 6533 393 6547 407
rect 6373 352 6387 366
rect 6433 352 6447 366
rect 6473 353 6487 367
rect 6353 273 6367 287
rect 6353 233 6367 247
rect 6333 193 6347 207
rect 6313 174 6327 188
rect 6413 173 6427 187
rect 5713 132 5727 146
rect 5853 133 5867 147
rect 5913 132 5927 146
rect 6013 133 6027 147
rect 6113 132 6127 146
rect 6273 133 6287 147
rect 6333 132 6347 146
rect 6373 132 6387 146
rect 6413 132 6427 146
rect 5653 113 5667 127
rect 6613 713 6627 727
rect 6653 694 6667 708
rect 6773 872 6787 886
rect 6773 813 6787 827
rect 6733 693 6747 707
rect 6633 652 6647 666
rect 6673 652 6687 666
rect 6593 533 6607 547
rect 6633 493 6647 507
rect 6593 394 6607 408
rect 6813 713 6827 727
rect 6813 673 6827 687
rect 6773 652 6787 666
rect 6853 1013 6867 1027
rect 6853 872 6867 886
rect 6993 1693 7007 1707
rect 7173 2732 7187 2746
rect 7213 2733 7227 2747
rect 7153 2593 7167 2607
rect 7153 2553 7167 2567
rect 7133 2533 7147 2547
rect 7093 2452 7107 2466
rect 7073 2393 7087 2407
rect 7093 2273 7107 2287
rect 7073 2253 7087 2267
rect 7073 1953 7087 1967
rect 7153 2452 7167 2466
rect 7213 2673 7227 2687
rect 7193 2493 7207 2507
rect 7133 2212 7147 2226
rect 7213 2452 7227 2466
rect 7313 2952 7327 2966
rect 7273 2913 7287 2927
rect 7273 2873 7287 2887
rect 7253 2432 7267 2446
rect 7233 2393 7247 2407
rect 7213 2353 7227 2367
rect 7253 2293 7267 2307
rect 7293 2593 7307 2607
rect 7453 4272 7467 4286
rect 7433 4233 7447 4247
rect 7573 4813 7587 4827
rect 7713 4813 7727 4827
rect 7553 4793 7567 4807
rect 7593 4653 7607 4667
rect 7553 4453 7567 4467
rect 7733 4793 7747 4807
rect 7993 5633 8007 5647
rect 7953 5453 7967 5467
rect 7873 5373 7887 5387
rect 8073 5733 8087 5747
rect 8113 5773 8127 5787
rect 8073 5633 8087 5647
rect 8033 5594 8047 5608
rect 8013 5553 8027 5567
rect 7993 5413 8007 5427
rect 8053 5552 8067 5566
rect 8093 5513 8107 5527
rect 8053 5473 8067 5487
rect 7893 5332 7907 5346
rect 7873 5233 7887 5247
rect 7833 5153 7847 5167
rect 7833 5093 7847 5107
rect 7853 5074 7867 5088
rect 8053 5374 8067 5388
rect 7993 5332 8007 5346
rect 7953 5293 7967 5307
rect 7933 5074 7947 5088
rect 7833 5033 7847 5047
rect 7913 5033 7927 5047
rect 7873 5013 7887 5027
rect 7933 5013 7947 5027
rect 7913 4973 7927 4987
rect 7912 4933 7926 4947
rect 7933 4933 7947 4947
rect 7873 4792 7887 4806
rect 7913 4792 7927 4806
rect 7813 4733 7827 4747
rect 7873 4713 7887 4727
rect 7813 4613 7827 4627
rect 7893 4693 7907 4707
rect 7873 4554 7887 4568
rect 7793 4493 7807 4507
rect 7673 4473 7687 4487
rect 7713 4473 7727 4487
rect 7853 4473 7867 4487
rect 7513 4393 7527 4407
rect 7613 4393 7627 4407
rect 7493 4373 7507 4387
rect 7533 4373 7547 4387
rect 7593 4334 7607 4348
rect 7633 4334 7647 4348
rect 7533 4292 7547 4306
rect 7573 4292 7587 4306
rect 7613 4292 7627 4306
rect 7613 4113 7627 4127
rect 7553 4073 7567 4087
rect 7513 4034 7527 4048
rect 7593 4034 7607 4048
rect 7533 3992 7547 4006
rect 7833 4373 7847 4387
rect 7693 4334 7707 4348
rect 7693 4293 7707 4307
rect 7813 4292 7827 4306
rect 7853 4292 7867 4306
rect 7973 4893 7987 4907
rect 7973 4593 7987 4607
rect 7953 4393 7967 4407
rect 7933 4293 7947 4307
rect 7893 4233 7907 4247
rect 7853 4213 7867 4227
rect 8033 5313 8047 5327
rect 8033 5292 8047 5306
rect 8013 5113 8027 5127
rect 8113 5473 8127 5487
rect 8113 5413 8127 5427
rect 8093 5213 8107 5227
rect 8073 5074 8087 5088
rect 8153 5973 8167 5987
rect 8213 6372 8227 6386
rect 8273 6653 8287 6667
rect 8253 6593 8267 6607
rect 8353 7773 8367 7787
rect 8333 7593 8347 7607
rect 8373 7633 8387 7647
rect 8433 7833 8447 7847
rect 8533 8273 8547 8287
rect 8493 8013 8507 8027
rect 8713 8333 8727 8347
rect 8673 8293 8687 8307
rect 8593 8213 8607 8227
rect 8633 8194 8647 8208
rect 8613 8152 8627 8166
rect 8653 8152 8667 8166
rect 8533 7974 8547 7988
rect 8573 7973 8587 7987
rect 8473 7833 8487 7847
rect 8453 7813 8467 7827
rect 8473 7793 8487 7807
rect 8533 7773 8547 7787
rect 8473 7693 8487 7707
rect 8513 7693 8527 7707
rect 8553 7673 8567 7687
rect 8493 7632 8507 7646
rect 8453 7613 8467 7627
rect 8373 7553 8387 7567
rect 8413 7553 8427 7567
rect 8513 7553 8527 7567
rect 8453 7493 8467 7507
rect 8373 7473 8387 7487
rect 8353 7454 8367 7468
rect 8393 7454 8407 7468
rect 8413 7393 8427 7407
rect 8373 7333 8387 7347
rect 8433 7333 8447 7347
rect 8413 7253 8427 7267
rect 8373 7153 8387 7167
rect 8433 7213 8447 7227
rect 8473 7453 8487 7467
rect 8473 7373 8487 7387
rect 8493 7132 8507 7146
rect 8333 7093 8347 7107
rect 8313 6893 8327 6907
rect 8493 7093 8507 7107
rect 8393 7053 8407 7067
rect 8493 7013 8507 7027
rect 8393 6953 8407 6967
rect 8573 7632 8587 7646
rect 8573 7573 8587 7587
rect 8833 8432 8847 8446
rect 8853 8413 8867 8427
rect 8893 8493 8907 8507
rect 9113 8833 9127 8847
rect 9013 8773 9027 8787
rect 8973 8714 8987 8728
rect 9313 8992 9327 9006
rect 9333 8873 9347 8887
rect 9173 8733 9187 8747
rect 9033 8672 9047 8686
rect 9193 8672 9207 8686
rect 9253 8672 9267 8686
rect 9033 8653 9047 8667
rect 8873 8373 8887 8387
rect 8853 8273 8867 8287
rect 8793 8233 8807 8247
rect 8913 8233 8927 8247
rect 8753 8213 8767 8227
rect 8753 8093 8767 8107
rect 8873 8194 8887 8208
rect 8993 8472 9007 8486
rect 9133 8472 9147 8486
rect 9293 8432 9307 8446
rect 9393 8853 9407 8867
rect 9353 8432 9367 8446
rect 9332 8393 9346 8407
rect 9353 8393 9367 8407
rect 9193 8313 9207 8327
rect 8993 8293 9007 8307
rect 8933 8193 8947 8207
rect 8953 8172 8967 8186
rect 8992 8172 9006 8186
rect 9013 8172 9027 8186
rect 9293 8213 9307 8227
rect 9533 9273 9547 9287
rect 9433 9093 9447 9107
rect 9513 9093 9527 9107
rect 9553 9233 9567 9247
rect 9553 9192 9567 9206
rect 9713 9553 9727 9567
rect 9773 9553 9787 9567
rect 9693 9433 9707 9447
rect 9633 9393 9647 9407
rect 9573 9093 9587 9107
rect 9473 8952 9487 8966
rect 9473 8913 9487 8927
rect 9453 8672 9467 8686
rect 9453 8651 9467 8665
rect 9433 8494 9447 8508
rect 9433 8293 9447 8307
rect 9393 8253 9407 8267
rect 8833 8152 8847 8166
rect 8853 8133 8867 8147
rect 9013 8153 9027 8167
rect 8893 8133 8907 8147
rect 8833 8113 8847 8127
rect 8913 8113 8927 8127
rect 8873 8073 8887 8087
rect 8793 8053 8807 8067
rect 8812 8013 8826 8027
rect 8833 8013 8847 8027
rect 8753 7974 8767 7988
rect 8833 7974 8847 7988
rect 8633 7933 8647 7947
rect 8593 7553 8607 7567
rect 8733 7913 8747 7927
rect 8773 7873 8787 7887
rect 8693 7674 8707 7688
rect 8713 7632 8727 7646
rect 8753 7553 8767 7567
rect 8633 7513 8647 7527
rect 8713 7493 8727 7507
rect 8553 7473 8567 7487
rect 8533 7453 8547 7467
rect 8613 7454 8627 7468
rect 8653 7454 8667 7468
rect 8693 7454 8707 7468
rect 8553 7412 8567 7426
rect 8593 7412 8607 7426
rect 8633 7393 8647 7407
rect 8713 7393 8727 7407
rect 8693 7293 8707 7307
rect 8613 7134 8627 7148
rect 8593 7033 8607 7047
rect 8573 7013 8587 7027
rect 8513 6933 8527 6947
rect 8593 6993 8607 7007
rect 8613 6934 8627 6948
rect 8413 6892 8427 6906
rect 8593 6892 8607 6906
rect 8633 6833 8647 6847
rect 8533 6813 8547 6827
rect 8333 6773 8347 6787
rect 8433 6614 8447 6628
rect 8733 6773 8747 6787
rect 8593 6713 8607 6727
rect 8633 6653 8647 6667
rect 8533 6553 8547 6567
rect 8573 6473 8587 6487
rect 8553 6434 8567 6448
rect 8273 6414 8287 6428
rect 8313 6414 8327 6428
rect 8333 6372 8347 6386
rect 8333 6233 8347 6247
rect 8233 6153 8247 6167
rect 8333 6114 8347 6128
rect 8213 5993 8227 6007
rect 8213 5894 8227 5908
rect 8333 6053 8347 6067
rect 8273 5953 8287 5967
rect 8313 5894 8327 5908
rect 8193 5853 8207 5867
rect 8193 5773 8207 5787
rect 8273 5852 8287 5866
rect 8233 5753 8247 5767
rect 8173 5673 8187 5687
rect 8273 5773 8287 5787
rect 8253 5633 8267 5647
rect 8153 5594 8167 5608
rect 8153 5513 8167 5527
rect 8033 5033 8047 5047
rect 8133 5032 8147 5046
rect 8093 4913 8107 4927
rect 8133 4913 8147 4927
rect 8073 4873 8087 4887
rect 8113 4873 8127 4887
rect 8153 4893 8167 4907
rect 8073 4733 8087 4747
rect 8013 4693 8027 4707
rect 8013 4553 8027 4567
rect 8153 4753 8167 4767
rect 8193 5613 8207 5627
rect 8233 5613 8247 5627
rect 8333 5753 8347 5767
rect 8193 5553 8207 5567
rect 8193 5513 8207 5527
rect 8293 5513 8307 5527
rect 8253 5413 8267 5427
rect 8293 5413 8307 5427
rect 8253 5374 8267 5388
rect 8313 5373 8327 5387
rect 8193 5293 8207 5307
rect 8193 5073 8207 5087
rect 8093 4593 8107 4607
rect 8113 4573 8127 4587
rect 8013 4512 8027 4526
rect 8053 4512 8067 4526
rect 7993 4473 8007 4487
rect 8053 4473 8067 4487
rect 8013 4334 8027 4348
rect 7993 4173 8007 4187
rect 8033 4173 8047 4187
rect 7833 4153 7847 4167
rect 7973 4153 7987 4167
rect 7813 4113 7827 4127
rect 7633 4053 7647 4067
rect 7673 4053 7687 4067
rect 7613 4013 7627 4027
rect 7553 3973 7567 3987
rect 7593 3973 7607 3987
rect 7473 3853 7487 3867
rect 7473 3814 7487 3828
rect 7513 3814 7527 3828
rect 7613 3913 7627 3927
rect 7593 3893 7607 3907
rect 7573 3814 7587 3828
rect 7433 3613 7447 3627
rect 7433 3393 7447 3407
rect 7433 3173 7447 3187
rect 7493 3772 7507 3786
rect 7553 3773 7567 3787
rect 7493 3713 7507 3727
rect 7473 3693 7487 3707
rect 7453 3153 7467 3167
rect 7493 3633 7507 3647
rect 7613 3813 7627 3827
rect 7593 3733 7607 3747
rect 7513 3573 7527 3587
rect 7573 3573 7587 3587
rect 7553 3514 7567 3528
rect 7593 3514 7607 3528
rect 7533 3472 7547 3486
rect 7533 3433 7547 3447
rect 7593 3373 7607 3387
rect 7533 3294 7547 3308
rect 7593 3293 7607 3307
rect 7553 3252 7567 3266
rect 7593 3233 7607 3247
rect 7513 3213 7527 3227
rect 7493 3153 7507 3167
rect 7473 3073 7487 3087
rect 7473 3013 7487 3027
rect 7433 2952 7447 2966
rect 7453 2913 7467 2927
rect 7413 2873 7427 2887
rect 7393 2793 7407 2807
rect 7353 2774 7367 2788
rect 7453 2754 7467 2768
rect 7353 2713 7367 2727
rect 7333 2613 7347 2627
rect 7313 2573 7327 2587
rect 7313 2433 7327 2447
rect 7293 2293 7307 2307
rect 7193 2212 7207 2226
rect 7233 2212 7247 2226
rect 7153 2173 7167 2187
rect 7213 2173 7227 2187
rect 7173 1993 7187 2007
rect 7293 2073 7307 2087
rect 7253 1993 7267 2007
rect 7213 1954 7227 1968
rect 7133 1913 7147 1927
rect 7193 1912 7207 1926
rect 7133 1873 7147 1887
rect 7113 1833 7127 1847
rect 7293 1973 7307 1987
rect 7253 1853 7267 1867
rect 7253 1793 7267 1807
rect 7193 1773 7207 1787
rect 7253 1753 7267 1767
rect 7113 1692 7127 1706
rect 7053 1613 7067 1627
rect 6993 1493 7007 1507
rect 7033 1453 7047 1467
rect 7073 1434 7087 1448
rect 6953 1413 6967 1427
rect 7013 1373 7027 1387
rect 7053 1353 7067 1367
rect 6993 1233 7007 1247
rect 7053 1233 7067 1247
rect 6933 1133 6947 1147
rect 6973 1113 6987 1127
rect 7013 1073 7027 1087
rect 7153 1593 7167 1607
rect 7273 1553 7287 1567
rect 7413 2732 7427 2746
rect 7433 2713 7447 2727
rect 7373 2693 7387 2707
rect 7413 2693 7427 2707
rect 7393 2432 7407 2446
rect 7453 2573 7467 2587
rect 7433 2513 7447 2527
rect 7333 2293 7347 2307
rect 7333 2173 7347 2187
rect 7333 2133 7347 2147
rect 7373 2173 7387 2187
rect 7353 2073 7367 2087
rect 7373 2053 7387 2067
rect 7433 2353 7447 2367
rect 7613 3133 7627 3147
rect 7553 3073 7567 3087
rect 7513 2933 7527 2947
rect 7513 2833 7527 2847
rect 7453 2293 7467 2307
rect 7433 2212 7447 2226
rect 7393 2033 7407 2047
rect 7413 2013 7427 2027
rect 7493 1933 7507 1947
rect 7313 1733 7327 1747
rect 7393 1912 7407 1926
rect 7393 1734 7407 1748
rect 7493 1813 7507 1827
rect 7473 1734 7487 1748
rect 7333 1633 7347 1647
rect 7433 1692 7447 1706
rect 7473 1693 7487 1707
rect 7373 1553 7387 1567
rect 7253 1513 7267 1527
rect 7293 1513 7307 1527
rect 7153 1453 7167 1467
rect 7253 1453 7267 1467
rect 7133 1433 7147 1447
rect 7233 1434 7247 1448
rect 7293 1433 7307 1447
rect 7413 1434 7427 1448
rect 7153 1333 7167 1347
rect 7233 1333 7247 1347
rect 7133 1313 7147 1327
rect 7173 1313 7187 1327
rect 7093 1253 7107 1267
rect 7233 1253 7247 1267
rect 7253 1253 7267 1267
rect 7193 1214 7207 1228
rect 7273 1214 7287 1228
rect 7073 1153 7087 1167
rect 7273 1173 7287 1187
rect 7173 1073 7187 1087
rect 7213 1073 7227 1087
rect 6993 933 7007 947
rect 7053 933 7067 947
rect 6753 593 6767 607
rect 6833 593 6847 607
rect 6813 553 6827 567
rect 6793 493 6807 507
rect 6773 473 6787 487
rect 6733 453 6747 467
rect 6553 353 6567 367
rect 6613 352 6627 366
rect 6913 652 6927 666
rect 6993 753 7007 767
rect 6973 694 6987 708
rect 6873 394 6887 408
rect 6793 352 6807 366
rect 6833 352 6847 366
rect 6773 313 6787 327
rect 6793 293 6807 307
rect 6853 233 6867 247
rect 6573 174 6587 188
rect 6793 174 6807 188
rect 6633 133 6647 147
rect 6773 132 6787 146
rect 6553 93 6567 107
rect 6433 73 6447 87
rect 6853 132 6867 146
rect 6813 53 6827 67
rect 6913 394 6927 408
rect 6913 353 6927 367
rect 7073 873 7087 887
rect 7153 813 7167 827
rect 7013 733 7027 747
rect 7093 694 7107 708
rect 7153 653 7167 667
rect 7113 633 7127 647
rect 7053 573 7067 587
rect 6993 513 7007 527
rect 7013 433 7027 447
rect 6953 393 6967 407
rect 6953 273 6967 287
rect 6953 173 6967 187
rect 7133 433 7147 447
rect 7093 394 7107 408
rect 7113 352 7127 366
rect 7073 313 7087 327
rect 7093 253 7107 267
rect 7053 174 7067 188
rect 6953 132 6967 146
rect 6993 132 7007 146
rect 6933 93 6947 107
rect 7433 1373 7447 1387
rect 7313 1333 7327 1347
rect 7293 1013 7307 1027
rect 7213 953 7227 967
rect 7293 953 7307 967
rect 7213 914 7227 928
rect 7233 872 7247 886
rect 7413 1214 7427 1228
rect 7533 2474 7547 2488
rect 7773 4034 7787 4048
rect 7813 4033 7827 4047
rect 7653 3853 7667 3867
rect 7693 4013 7707 4027
rect 7793 3992 7807 4006
rect 7753 3913 7767 3927
rect 7813 3853 7827 3867
rect 7693 3813 7707 3827
rect 7753 3794 7767 3808
rect 7793 3794 7807 3808
rect 7953 4133 7967 4147
rect 7853 4073 7867 4087
rect 7953 4073 7967 4087
rect 7673 3513 7687 3527
rect 7833 3793 7847 3807
rect 7793 3653 7807 3667
rect 7833 3573 7847 3587
rect 7713 3514 7727 3528
rect 7793 3514 7807 3528
rect 7692 3473 7706 3487
rect 7713 3473 7727 3487
rect 7773 3472 7787 3486
rect 7793 3453 7807 3467
rect 7712 3433 7726 3447
rect 7733 3433 7747 3447
rect 7733 3393 7747 3407
rect 7793 3373 7807 3387
rect 7673 3353 7687 3367
rect 7773 3353 7787 3367
rect 7713 3313 7727 3327
rect 7753 3294 7767 3308
rect 7793 3293 7807 3307
rect 8133 4334 8147 4348
rect 8113 4273 8127 4287
rect 8113 4213 8127 4227
rect 8133 4133 8147 4147
rect 8033 4053 8047 4067
rect 8113 4053 8127 4067
rect 7973 3992 7987 4006
rect 8073 3993 8087 4007
rect 8173 4613 8187 4627
rect 8013 3953 8027 3967
rect 8153 3953 8167 3967
rect 8153 3813 8167 3827
rect 8013 3793 8027 3807
rect 8213 4613 8227 4627
rect 8253 5253 8267 5267
rect 8353 5673 8367 5687
rect 8373 5594 8387 5608
rect 8353 5533 8367 5547
rect 8333 5313 8347 5327
rect 8473 6414 8487 6428
rect 8513 6414 8527 6428
rect 8553 6413 8567 6427
rect 8593 6433 8607 6447
rect 8473 6373 8487 6387
rect 8473 6313 8487 6327
rect 8553 6153 8567 6167
rect 8453 6053 8467 6067
rect 8533 6053 8547 6067
rect 8493 5993 8507 6007
rect 8473 5733 8487 5747
rect 8413 5713 8427 5727
rect 8413 5653 8427 5667
rect 8393 5513 8407 5527
rect 8393 5433 8407 5447
rect 8373 5413 8387 5427
rect 8393 5193 8407 5207
rect 8373 5153 8387 5167
rect 8353 5093 8367 5107
rect 8313 5074 8327 5088
rect 8333 5032 8347 5046
rect 8313 4993 8327 5007
rect 8273 4933 8287 4947
rect 8353 4854 8367 4868
rect 8253 4813 8267 4827
rect 8253 4753 8267 4767
rect 8233 4573 8247 4587
rect 8193 4353 8207 4367
rect 8193 4233 8207 4247
rect 8333 4812 8347 4826
rect 8533 5773 8547 5787
rect 8493 5713 8507 5727
rect 8553 5653 8567 5667
rect 8513 5594 8527 5608
rect 8813 7933 8827 7947
rect 8793 7633 8807 7647
rect 8893 8053 8907 8067
rect 8873 7853 8887 7867
rect 8833 7613 8847 7627
rect 8833 7493 8847 7507
rect 8853 7453 8867 7467
rect 8813 7412 8827 7426
rect 8813 7353 8827 7367
rect 8773 7333 8787 7347
rect 8793 7073 8807 7087
rect 8833 7253 8847 7267
rect 8813 6973 8827 6987
rect 9193 8013 9207 8027
rect 8913 7974 8927 7988
rect 8973 7974 8987 7988
rect 9013 7974 9027 7988
rect 9093 7973 9107 7987
rect 9233 7974 9247 7988
rect 8953 7932 8967 7946
rect 9053 7913 9067 7927
rect 8993 7893 9007 7907
rect 9053 7873 9067 7887
rect 9033 7853 9047 7867
rect 9033 7793 9047 7807
rect 8993 7713 9007 7727
rect 8893 7673 8907 7687
rect 8953 7674 8967 7688
rect 8933 7632 8947 7646
rect 8913 7613 8927 7627
rect 8893 7454 8907 7468
rect 8893 7333 8907 7347
rect 8813 6934 8827 6948
rect 8833 6892 8847 6906
rect 9033 7673 9047 7687
rect 8993 7593 9007 7607
rect 8933 7573 8947 7587
rect 8913 7093 8927 7107
rect 8853 6833 8867 6847
rect 8813 6634 8827 6648
rect 8793 6592 8807 6606
rect 8893 6553 8907 6567
rect 8833 6473 8847 6487
rect 8833 6433 8847 6447
rect 8773 6414 8787 6428
rect 8813 6414 8827 6428
rect 8673 6373 8687 6387
rect 8873 6413 8887 6427
rect 8713 6372 8727 6386
rect 8753 6372 8767 6386
rect 8793 6372 8807 6386
rect 8833 6372 8847 6386
rect 9073 7673 9087 7687
rect 9053 7633 9067 7647
rect 9033 7533 9047 7547
rect 8973 7493 8987 7507
rect 9253 7932 9267 7946
rect 9393 8193 9407 8207
rect 9293 7913 9307 7927
rect 9393 8113 9407 8127
rect 9373 8093 9387 8107
rect 9413 8093 9427 8107
rect 9553 8992 9567 9006
rect 9593 8994 9607 9008
rect 9653 9234 9667 9248
rect 9753 9493 9767 9507
rect 9853 9533 9867 9547
rect 9913 9534 9927 9548
rect 10033 9534 10047 9548
rect 9853 9492 9867 9506
rect 9933 9492 9947 9506
rect 9793 9453 9807 9467
rect 9993 9453 10007 9467
rect 10093 9913 10107 9927
rect 10433 10012 10447 10026
rect 10333 9833 10347 9847
rect 10213 9813 10227 9827
rect 10653 10033 10667 10047
rect 10533 10012 10547 10026
rect 10613 10012 10627 10026
rect 10573 9973 10587 9987
rect 10493 9913 10507 9927
rect 10653 9913 10667 9927
rect 10813 10532 10827 10546
rect 10733 10493 10747 10507
rect 10713 9933 10727 9947
rect 10613 9813 10627 9827
rect 10473 9773 10487 9787
rect 10253 9754 10267 9768
rect 10433 9754 10447 9768
rect 10513 9753 10527 9767
rect 10093 9733 10107 9747
rect 10113 9534 10127 9548
rect 10173 9534 10187 9548
rect 10453 9712 10467 9726
rect 10233 9673 10247 9687
rect 10253 9633 10267 9647
rect 10093 9493 10107 9507
rect 10073 9473 10087 9487
rect 10153 9492 10167 9506
rect 10233 9534 10247 9548
rect 10113 9393 10127 9407
rect 9733 9313 9747 9327
rect 9913 9313 9927 9327
rect 10033 9313 10047 9327
rect 9873 9273 9887 9287
rect 9993 9234 10007 9248
rect 9893 9192 9907 9206
rect 9993 9193 10007 9207
rect 10453 9593 10467 9607
rect 10393 9393 10407 9407
rect 10313 9313 10327 9327
rect 10073 9234 10087 9248
rect 10113 9234 10127 9248
rect 10253 9234 10267 9248
rect 10033 9192 10047 9206
rect 10053 9153 10067 9167
rect 9713 9133 9727 9147
rect 9893 9133 9907 9147
rect 9693 9093 9707 9107
rect 10033 9113 10047 9127
rect 9933 8952 9947 8966
rect 9773 8913 9787 8927
rect 9633 8853 9647 8867
rect 9973 8873 9987 8887
rect 9933 8833 9947 8847
rect 9593 8733 9607 8747
rect 9573 8672 9587 8686
rect 9513 8653 9527 8667
rect 9533 8513 9547 8527
rect 9573 8513 9587 8527
rect 9493 8494 9507 8508
rect 9513 8452 9527 8466
rect 9573 8413 9587 8427
rect 9493 8393 9507 8407
rect 9513 8373 9527 8387
rect 9493 8313 9507 8327
rect 9473 8153 9487 8167
rect 9473 8053 9487 8067
rect 9453 8033 9467 8047
rect 9413 7993 9427 8007
rect 9333 7974 9347 7988
rect 9373 7974 9387 7988
rect 9453 7974 9467 7988
rect 9373 7933 9387 7947
rect 9333 7913 9347 7927
rect 9433 7893 9447 7907
rect 10053 8994 10067 9008
rect 10133 9192 10147 9206
rect 10353 9133 10367 9147
rect 10353 9093 10367 9107
rect 10433 9153 10447 9167
rect 10333 9053 10347 9067
rect 10233 8992 10247 9006
rect 10333 8992 10347 9006
rect 10093 8913 10107 8927
rect 10133 8833 10147 8847
rect 10033 8793 10047 8807
rect 9633 8734 9647 8748
rect 9713 8734 9727 8748
rect 9773 8713 9787 8727
rect 9873 8713 9887 8727
rect 9613 8693 9627 8707
rect 9753 8692 9767 8706
rect 9753 8653 9767 8667
rect 10053 8633 10067 8647
rect 9752 8593 9766 8607
rect 9773 8593 9787 8607
rect 9953 8593 9967 8607
rect 9673 8573 9687 8587
rect 9753 8513 9767 8527
rect 9613 8493 9627 8507
rect 9713 8494 9727 8508
rect 9893 8494 9907 8508
rect 9993 8533 10007 8547
rect 9993 8494 10007 8508
rect 10113 8494 10127 8508
rect 9593 8313 9607 8327
rect 9733 8452 9747 8466
rect 9773 8452 9787 8466
rect 9873 8452 9887 8466
rect 9813 8313 9827 8327
rect 9853 8313 9867 8327
rect 9613 8293 9627 8307
rect 9653 8174 9667 8188
rect 9753 8174 9767 8188
rect 9773 8153 9787 8167
rect 9693 8073 9707 8087
rect 9753 8073 9767 8087
rect 9793 8073 9807 8087
rect 9593 8013 9607 8027
rect 9573 7974 9587 7988
rect 9513 7873 9527 7887
rect 9313 7793 9327 7807
rect 9573 7773 9587 7787
rect 9253 7733 9267 7747
rect 9233 7693 9247 7707
rect 9153 7674 9167 7688
rect 9133 7632 9147 7646
rect 9193 7632 9207 7646
rect 9093 7573 9107 7587
rect 9073 7473 9087 7487
rect 9013 7454 9027 7468
rect 9053 7454 9067 7468
rect 9073 7412 9087 7426
rect 8953 7293 8967 7307
rect 8973 7253 8987 7267
rect 9033 7253 9047 7267
rect 8953 6793 8967 6807
rect 9053 7233 9067 7247
rect 9173 7573 9187 7587
rect 9133 7473 9147 7487
rect 9113 7173 9127 7187
rect 9173 7453 9187 7467
rect 9093 7154 9107 7168
rect 9133 7154 9147 7168
rect 9153 7132 9167 7146
rect 9092 7093 9106 7107
rect 9113 7093 9127 7107
rect 9073 7053 9087 7067
rect 9073 6973 9087 6987
rect 9173 7053 9187 7067
rect 9213 7533 9227 7547
rect 9313 7693 9327 7707
rect 9653 7974 9667 7988
rect 9753 8052 9767 8066
rect 9613 7694 9627 7708
rect 9673 7893 9687 7907
rect 9693 7873 9707 7887
rect 9293 7654 9307 7668
rect 9273 7533 9287 7547
rect 9453 7654 9467 7668
rect 9573 7652 9587 7666
rect 9313 7613 9327 7627
rect 9593 7613 9607 7627
rect 9533 7553 9547 7567
rect 9393 7533 9407 7547
rect 9253 7473 9267 7487
rect 9313 7513 9327 7527
rect 9213 7412 9227 7426
rect 9293 7412 9307 7426
rect 9493 7473 9507 7487
rect 9513 7412 9527 7426
rect 9553 7412 9567 7426
rect 9493 7213 9507 7227
rect 9553 7213 9567 7227
rect 9393 7173 9407 7187
rect 9213 7132 9227 7146
rect 9253 7134 9267 7148
rect 9393 7134 9407 7148
rect 9253 7093 9267 7107
rect 9213 7073 9227 7087
rect 9093 6934 9107 6948
rect 9153 6934 9167 6948
rect 9073 6892 9087 6906
rect 8993 6733 9007 6747
rect 9113 6733 9127 6747
rect 9033 6693 9047 6707
rect 9113 6693 9127 6707
rect 9053 6634 9067 6648
rect 8993 6592 9007 6606
rect 9033 6592 9047 6606
rect 9073 6553 9087 6567
rect 8973 6533 8987 6547
rect 9053 6533 9067 6547
rect 9033 6473 9047 6487
rect 8973 6433 8987 6447
rect 8913 6333 8927 6347
rect 8893 6313 8907 6327
rect 8813 6233 8827 6247
rect 8753 6193 8767 6207
rect 8733 6013 8747 6027
rect 8693 5993 8707 6007
rect 8633 5953 8647 5967
rect 8773 5953 8787 5967
rect 8733 5913 8747 5927
rect 8673 5894 8687 5908
rect 8733 5894 8747 5908
rect 8693 5852 8707 5866
rect 8753 5852 8767 5866
rect 8673 5833 8687 5847
rect 8733 5713 8747 5727
rect 8612 5593 8626 5607
rect 8633 5594 8647 5608
rect 8673 5594 8687 5608
rect 8753 5613 8767 5627
rect 8453 5533 8467 5547
rect 8533 5553 8547 5567
rect 8573 5553 8587 5567
rect 8613 5553 8627 5567
rect 8493 5493 8507 5507
rect 8453 5473 8467 5487
rect 8553 5513 8567 5527
rect 8533 5433 8547 5447
rect 8493 5413 8507 5427
rect 8473 5313 8487 5327
rect 8513 5273 8527 5287
rect 8433 5213 8447 5227
rect 8413 4973 8427 4987
rect 8413 4893 8427 4907
rect 8413 4773 8427 4787
rect 8593 5373 8607 5387
rect 8553 5193 8567 5207
rect 8553 5093 8567 5107
rect 8633 5493 8647 5507
rect 8713 5374 8727 5388
rect 8613 5273 8627 5287
rect 8653 5133 8667 5147
rect 8533 5013 8547 5027
rect 8453 4973 8467 4987
rect 8293 4693 8307 4707
rect 8353 4693 8367 4707
rect 8333 4573 8347 4587
rect 8353 4553 8367 4567
rect 8373 4532 8387 4546
rect 8353 4513 8367 4527
rect 8253 4473 8267 4487
rect 8313 4473 8327 4487
rect 8273 4413 8287 4427
rect 8253 4373 8267 4387
rect 8273 4353 8287 4367
rect 8293 4213 8307 4227
rect 8253 4173 8267 4187
rect 8233 4053 8247 4067
rect 8333 4213 8347 4227
rect 8333 4113 8347 4127
rect 8233 3992 8247 4006
rect 8213 3813 8227 3827
rect 8253 3813 8267 3827
rect 7993 3753 8007 3767
rect 7893 3633 7907 3647
rect 7873 3533 7887 3547
rect 7853 3293 7867 3307
rect 7973 3593 7987 3607
rect 7913 3553 7927 3567
rect 7893 3353 7907 3367
rect 7693 3253 7707 3267
rect 7653 3193 7667 3207
rect 7773 3252 7787 3266
rect 7733 3233 7747 3247
rect 7793 3233 7807 3247
rect 7693 3173 7707 3187
rect 7633 3013 7647 3027
rect 7653 2952 7667 2966
rect 7773 3053 7787 3067
rect 7773 3013 7787 3027
rect 7713 2853 7727 2867
rect 7693 2633 7707 2647
rect 7753 2613 7767 2627
rect 7832 3193 7846 3207
rect 7853 3193 7867 3207
rect 7873 3073 7887 3087
rect 7933 3514 7947 3528
rect 8153 3733 8167 3747
rect 8093 3693 8107 3707
rect 7993 3553 8007 3567
rect 8013 3514 8027 3528
rect 7933 3473 7947 3487
rect 8033 3472 8047 3486
rect 7993 3453 8007 3467
rect 8093 3453 8107 3467
rect 8053 3253 8067 3267
rect 8073 3233 8087 3247
rect 8173 3713 8187 3727
rect 8253 3773 8267 3787
rect 8313 3993 8327 4007
rect 8373 4093 8387 4107
rect 8353 3933 8367 3947
rect 8313 3913 8327 3927
rect 8433 4753 8447 4767
rect 8473 4913 8487 4927
rect 8453 4573 8467 4587
rect 8453 4533 8467 4547
rect 8433 4453 8447 4467
rect 8433 4373 8447 4387
rect 8413 4253 8427 4267
rect 8613 5033 8627 5047
rect 8733 5273 8747 5287
rect 8853 6173 8867 6187
rect 8833 6013 8847 6027
rect 8813 5894 8827 5908
rect 8793 5852 8807 5866
rect 8813 5653 8827 5667
rect 8953 6273 8967 6287
rect 8953 6153 8967 6167
rect 9053 6273 9067 6287
rect 9453 7013 9467 7027
rect 9293 6993 9307 7007
rect 9333 6973 9347 6987
rect 9393 6933 9407 6947
rect 9313 6892 9327 6906
rect 9373 6892 9387 6906
rect 9353 6873 9367 6887
rect 9353 6793 9367 6807
rect 9273 6634 9287 6648
rect 9173 6593 9187 6607
rect 9453 6893 9467 6907
rect 9393 6873 9407 6887
rect 9613 7293 9627 7307
rect 9673 7653 9687 7667
rect 9673 7513 9687 7527
rect 9733 7693 9747 7707
rect 9733 7593 9747 7607
rect 9973 8452 9987 8466
rect 9893 8373 9907 8387
rect 9893 8213 9907 8227
rect 9973 8293 9987 8307
rect 9953 8153 9967 8167
rect 9913 8133 9927 8147
rect 9872 8073 9886 8087
rect 9893 8073 9907 8087
rect 9913 8053 9927 8067
rect 9853 8013 9867 8027
rect 9933 7993 9947 8007
rect 9813 7974 9827 7988
rect 9853 7974 9867 7988
rect 9813 7713 9827 7727
rect 9953 7913 9967 7927
rect 9933 7833 9947 7847
rect 10013 8293 10027 8307
rect 10013 8233 10027 8247
rect 9993 8193 10007 8207
rect 10053 8194 10067 8208
rect 10093 8194 10107 8208
rect 10033 8152 10047 8166
rect 10073 8152 10087 8166
rect 10273 8714 10287 8728
rect 10233 8593 10247 8607
rect 10233 8533 10247 8547
rect 10193 8494 10207 8508
rect 10373 8813 10387 8827
rect 10473 9533 10487 9547
rect 10613 9553 10627 9567
rect 10573 9534 10587 9548
rect 10673 9712 10687 9726
rect 10593 9492 10607 9506
rect 10513 9473 10527 9487
rect 10553 9473 10567 9487
rect 10493 9234 10507 9248
rect 10533 9234 10547 9248
rect 10713 9633 10727 9647
rect 10813 10393 10827 10407
rect 10853 10393 10867 10407
rect 10773 10353 10787 10367
rect 10753 10073 10767 10087
rect 10773 10053 10787 10067
rect 10813 10073 10827 10087
rect 10793 10012 10807 10026
rect 10833 10012 10847 10026
rect 10933 10613 10947 10627
rect 10913 10573 10927 10587
rect 10913 10532 10927 10546
rect 10913 10273 10927 10287
rect 10913 10012 10927 10026
rect 10813 9953 10827 9967
rect 10893 9953 10907 9967
rect 10753 9773 10767 9787
rect 10753 9712 10767 9726
rect 10733 9593 10747 9607
rect 10913 9813 10927 9827
rect 10873 9754 10887 9768
rect 10993 10752 11007 10766
rect 11073 10752 11087 10766
rect 11033 10733 11047 10747
rect 11233 10693 11247 10707
rect 11033 10613 11047 10627
rect 10953 10574 10967 10588
rect 10993 10574 11007 10588
rect 11153 10573 11167 10587
rect 11233 10574 11247 10588
rect 11013 10532 11027 10546
rect 11053 10532 11067 10546
rect 11133 10532 11147 10546
rect 10953 10433 10967 10447
rect 11013 10274 11027 10288
rect 10993 10232 11007 10246
rect 11033 10193 11047 10207
rect 10993 10133 11007 10147
rect 10973 10053 10987 10067
rect 10953 10012 10967 10026
rect 10893 9712 10907 9726
rect 10853 9633 10867 9647
rect 10853 9553 10867 9567
rect 10833 9492 10847 9506
rect 10793 9453 10807 9467
rect 10713 9413 10727 9427
rect 10513 9153 10527 9167
rect 10593 9153 10607 9167
rect 10973 9754 10987 9768
rect 11033 10093 11047 10107
rect 11073 10054 11087 10068
rect 11093 10012 11107 10026
rect 11053 9973 11067 9987
rect 11053 9952 11067 9966
rect 11133 9953 11147 9967
rect 10993 9712 11007 9726
rect 10973 9593 10987 9607
rect 11213 10532 11227 10546
rect 11333 10532 11347 10546
rect 11253 10493 11267 10507
rect 11253 10133 11267 10147
rect 11293 10093 11307 10107
rect 11193 9973 11207 9987
rect 11153 9813 11167 9827
rect 11213 9813 11227 9827
rect 11073 9712 11087 9726
rect 11033 9413 11047 9427
rect 10913 9353 10927 9367
rect 10953 9353 10967 9367
rect 10773 9254 10787 9268
rect 10733 9173 10747 9187
rect 10673 9113 10687 9127
rect 10713 9113 10727 9127
rect 10633 9053 10647 9067
rect 10593 9014 10607 9028
rect 10693 9033 10707 9047
rect 10473 8972 10487 8986
rect 10613 8972 10627 8986
rect 10653 8972 10667 8986
rect 10693 8972 10707 8986
rect 10453 8833 10467 8847
rect 10633 8833 10647 8847
rect 10433 8773 10447 8787
rect 10373 8734 10387 8748
rect 10313 8714 10327 8728
rect 10293 8673 10307 8687
rect 10393 8653 10407 8667
rect 11113 9492 11127 9506
rect 11153 9493 11167 9507
rect 11013 9333 11027 9347
rect 11073 9333 11087 9347
rect 10853 9033 10867 9047
rect 11073 9254 11087 9268
rect 11033 9193 11047 9207
rect 11013 9014 11027 9028
rect 11053 9014 11067 9028
rect 11093 9014 11107 9028
rect 10873 8972 10887 8986
rect 10953 8973 10967 8987
rect 10833 8893 10847 8907
rect 10833 8872 10847 8886
rect 10793 8734 10807 8748
rect 10753 8692 10767 8706
rect 10453 8633 10467 8647
rect 10453 8573 10467 8587
rect 10533 8573 10547 8587
rect 10453 8513 10467 8527
rect 10333 8494 10347 8508
rect 10413 8494 10427 8508
rect 10213 8452 10227 8466
rect 10173 8393 10187 8407
rect 10233 8233 10247 8247
rect 10173 8193 10187 8207
rect 10213 8173 10227 8187
rect 10193 8153 10207 8167
rect 10053 8133 10067 8147
rect 10013 8093 10027 8107
rect 10073 8093 10087 8107
rect 10193 8093 10207 8107
rect 10053 8073 10067 8087
rect 10073 8053 10087 8067
rect 10113 7974 10127 7988
rect 10173 7954 10187 7968
rect 10013 7873 10027 7887
rect 9993 7833 10007 7847
rect 9973 7753 9987 7767
rect 10153 7933 10167 7947
rect 10133 7913 10147 7927
rect 10013 7793 10027 7807
rect 10093 7793 10107 7807
rect 10013 7653 10027 7667
rect 9852 7593 9866 7607
rect 9873 7593 9887 7607
rect 9993 7593 10007 7607
rect 9753 7533 9767 7547
rect 9653 7093 9667 7107
rect 9593 7013 9607 7027
rect 9533 6934 9547 6948
rect 9573 6934 9587 6948
rect 9553 6892 9567 6906
rect 9713 7493 9727 7507
rect 9793 7493 9807 7507
rect 9693 7453 9707 7467
rect 9753 7454 9767 7468
rect 10133 7632 10147 7646
rect 10193 7873 10207 7887
rect 10193 7793 10207 7807
rect 10493 8474 10507 8488
rect 10573 8513 10587 8527
rect 10593 8493 10607 8507
rect 10473 8453 10487 8467
rect 10473 8393 10487 8407
rect 10393 8293 10407 8307
rect 10513 8233 10527 8247
rect 10573 8473 10587 8487
rect 10733 8453 10747 8467
rect 10933 8694 10947 8708
rect 10913 8633 10927 8647
rect 10853 8573 10867 8587
rect 10853 8493 10867 8507
rect 10693 8353 10707 8367
rect 10833 8353 10847 8367
rect 10633 8313 10647 8327
rect 10533 8213 10547 8227
rect 10373 8073 10387 8087
rect 10533 8152 10547 8166
rect 10573 8152 10587 8166
rect 10513 8133 10527 8147
rect 10313 8053 10327 8067
rect 10353 8053 10367 8067
rect 10493 8053 10507 8067
rect 10273 7953 10287 7967
rect 10413 7833 10427 7847
rect 10313 7793 10327 7807
rect 10473 7793 10487 7807
rect 10193 7713 10207 7727
rect 10053 7573 10067 7587
rect 10093 7573 10107 7587
rect 9893 7553 9907 7567
rect 9893 7453 9907 7467
rect 9853 7433 9867 7447
rect 9693 7412 9707 7426
rect 9693 7353 9707 7367
rect 9673 6934 9687 6948
rect 9573 6833 9587 6847
rect 9493 6793 9507 6807
rect 9573 6793 9587 6807
rect 9473 6753 9487 6767
rect 9513 6753 9527 6767
rect 9553 6733 9567 6747
rect 9473 6693 9487 6707
rect 9373 6673 9387 6687
rect 9253 6493 9267 6507
rect 9213 6433 9227 6447
rect 9173 6414 9187 6428
rect 9193 6372 9207 6386
rect 9533 6613 9547 6627
rect 9513 6593 9527 6607
rect 9493 6553 9507 6567
rect 9453 6513 9467 6527
rect 9413 6453 9427 6467
rect 9453 6433 9467 6447
rect 9373 6373 9387 6387
rect 9433 6372 9447 6386
rect 9473 6372 9487 6386
rect 9353 6313 9367 6327
rect 9413 6313 9427 6327
rect 9253 6293 9267 6307
rect 9133 6233 9147 6247
rect 9233 6233 9247 6247
rect 9113 6193 9127 6207
rect 9093 6173 9107 6187
rect 9033 6153 9047 6167
rect 8993 6114 9007 6128
rect 9033 6092 9047 6106
rect 8893 6033 8907 6047
rect 8853 5993 8867 6007
rect 8873 5953 8887 5967
rect 8873 5813 8887 5827
rect 8853 5773 8867 5787
rect 8993 6053 9007 6067
rect 8973 5953 8987 5967
rect 9113 6094 9127 6108
rect 9113 6053 9127 6067
rect 9093 6033 9107 6047
rect 9413 6273 9427 6287
rect 9493 6353 9507 6367
rect 9433 6253 9447 6267
rect 9473 6233 9487 6247
rect 9253 6193 9267 6207
rect 9433 6134 9447 6148
rect 9473 6134 9487 6148
rect 9273 6094 9287 6108
rect 9373 6093 9387 6107
rect 9373 6033 9387 6047
rect 9133 5973 9147 5987
rect 8913 5913 8927 5927
rect 8933 5894 8947 5908
rect 9053 5913 9067 5927
rect 9053 5873 9067 5887
rect 8953 5852 8967 5866
rect 9033 5832 9047 5846
rect 8993 5813 9007 5827
rect 9193 5872 9207 5886
rect 9333 5872 9347 5886
rect 9193 5832 9207 5846
rect 9093 5713 9107 5727
rect 9213 5713 9227 5727
rect 9313 5713 9327 5727
rect 8893 5613 8907 5627
rect 9193 5614 9207 5628
rect 8793 5572 8807 5586
rect 8833 5572 8847 5586
rect 8813 5533 8827 5547
rect 8713 5253 8727 5267
rect 8773 5253 8787 5267
rect 8693 5074 8707 5088
rect 8673 5013 8687 5027
rect 8653 4933 8667 4947
rect 8573 4913 8587 4927
rect 8533 4873 8547 4887
rect 8493 4854 8507 4868
rect 9033 5574 9047 5588
rect 9253 5614 9267 5628
rect 9153 5572 9167 5586
rect 9233 5573 9247 5587
rect 9133 5553 9147 5567
rect 8853 5533 8867 5547
rect 8893 5533 8907 5547
rect 8833 5374 8847 5388
rect 8873 5453 8887 5467
rect 8853 5333 8867 5347
rect 8953 5433 8967 5447
rect 8913 5374 8927 5388
rect 9233 5513 9247 5527
rect 9173 5433 9187 5447
rect 9113 5333 9127 5347
rect 8933 5313 8947 5327
rect 8873 5233 8887 5247
rect 9033 5193 9047 5207
rect 8893 5173 8907 5187
rect 8773 5074 8787 5088
rect 8713 5013 8727 5027
rect 8813 5013 8827 5027
rect 8793 4993 8807 5007
rect 8713 4973 8727 4987
rect 8693 4853 8707 4867
rect 8753 4854 8767 4868
rect 8493 4813 8507 4827
rect 8553 4812 8567 4826
rect 8693 4813 8707 4827
rect 8493 4713 8507 4727
rect 8613 4534 8627 4548
rect 8733 4773 8747 4787
rect 8773 4773 8787 4787
rect 8733 4532 8747 4546
rect 8713 4493 8727 4507
rect 8773 4493 8787 4507
rect 8713 4453 8727 4467
rect 8513 4433 8527 4447
rect 8553 4433 8567 4447
rect 8533 4413 8547 4427
rect 8513 4393 8527 4407
rect 8553 4373 8567 4387
rect 8533 4353 8547 4367
rect 8493 4292 8507 4306
rect 8433 4153 8447 4167
rect 8493 4113 8507 4127
rect 8513 4053 8527 4067
rect 8393 4034 8407 4048
rect 8473 4034 8487 4048
rect 8333 3873 8347 3887
rect 8373 3873 8387 3887
rect 8293 3853 8307 3867
rect 8273 3653 8287 3667
rect 8253 3573 8267 3587
rect 8453 3973 8467 3987
rect 8453 3933 8467 3947
rect 8393 3853 8407 3867
rect 8373 3814 8387 3828
rect 8473 3813 8487 3827
rect 8353 3772 8367 3786
rect 8313 3713 8327 3727
rect 8293 3533 8307 3547
rect 8212 3433 8226 3447
rect 8233 3433 8247 3447
rect 8213 3393 8227 3407
rect 8273 3353 8287 3367
rect 8173 3313 8187 3327
rect 8253 3313 8267 3327
rect 8173 3274 8187 3288
rect 8193 3233 8207 3247
rect 8233 3233 8247 3247
rect 8033 3033 8047 3047
rect 7913 2993 7927 3007
rect 7973 2993 7987 3007
rect 8013 2994 8027 3008
rect 7893 2952 7907 2966
rect 7933 2833 7947 2847
rect 7893 2793 7907 2807
rect 7833 2753 7847 2767
rect 7913 2753 7927 2767
rect 7893 2732 7907 2746
rect 7853 2712 7867 2726
rect 7873 2693 7887 2707
rect 7853 2673 7867 2687
rect 7733 2593 7747 2607
rect 7693 2533 7707 2547
rect 7633 2493 7647 2507
rect 7593 2474 7607 2488
rect 7693 2473 7707 2487
rect 7533 2333 7547 2347
rect 7533 2233 7547 2247
rect 7653 2432 7667 2446
rect 7693 2432 7707 2446
rect 7613 2393 7627 2407
rect 7633 2293 7647 2307
rect 7573 2173 7587 2187
rect 7653 2153 7667 2167
rect 7713 2093 7727 2107
rect 7673 2033 7687 2047
rect 7653 1893 7667 1907
rect 7573 1773 7587 1787
rect 7513 1734 7527 1748
rect 7613 1734 7627 1748
rect 7753 2233 7767 2247
rect 7813 2474 7827 2488
rect 7953 2773 7967 2787
rect 7953 2633 7967 2647
rect 7933 2533 7947 2547
rect 7913 2513 7927 2527
rect 7853 2473 7867 2487
rect 7893 2453 7907 2467
rect 7833 2432 7847 2446
rect 7873 2433 7887 2447
rect 7953 2454 7967 2468
rect 7953 2393 7967 2407
rect 7913 2313 7927 2327
rect 7953 2313 7967 2327
rect 7913 2254 7927 2268
rect 7773 2213 7787 2227
rect 7853 2212 7867 2226
rect 7833 2053 7847 2067
rect 7933 2073 7947 2087
rect 7913 1913 7927 1927
rect 7953 1993 7967 2007
rect 7933 1893 7947 1907
rect 7733 1813 7747 1827
rect 7813 1813 7827 1827
rect 7853 1813 7867 1827
rect 8093 2994 8107 3008
rect 8133 2994 8147 3008
rect 8033 2953 8047 2967
rect 8113 2933 8127 2947
rect 8073 2893 8087 2907
rect 8113 2893 8127 2907
rect 8073 2774 8087 2788
rect 8113 2774 8127 2788
rect 8153 2774 8167 2788
rect 8053 2732 8067 2746
rect 8093 2732 8107 2746
rect 8013 2673 8027 2687
rect 8193 2933 8207 2947
rect 8193 2853 8207 2867
rect 8293 3333 8307 3347
rect 8273 3073 8287 3087
rect 8213 2833 8227 2847
rect 8193 2813 8207 2827
rect 8173 2673 8187 2687
rect 8213 2673 8227 2687
rect 8193 2633 8207 2647
rect 8153 2593 8167 2607
rect 8113 2454 8127 2468
rect 8253 2833 8267 2847
rect 8313 3233 8327 3247
rect 8453 3773 8467 3787
rect 8393 3733 8407 3747
rect 8373 3653 8387 3667
rect 8353 3213 8367 3227
rect 8313 3193 8327 3207
rect 8293 2993 8307 3007
rect 8513 3893 8527 3907
rect 8533 3853 8547 3867
rect 8533 3772 8547 3786
rect 8513 3733 8527 3747
rect 8493 3593 8507 3607
rect 8473 3573 8487 3587
rect 8433 3553 8447 3567
rect 8533 3553 8547 3567
rect 8633 4334 8647 4348
rect 8673 4334 8687 4348
rect 8853 4813 8867 4827
rect 8833 4633 8847 4647
rect 8833 4413 8847 4427
rect 8853 4373 8867 4387
rect 8633 4293 8647 4307
rect 8733 4292 8747 4306
rect 8773 4293 8787 4307
rect 8813 4293 8827 4307
rect 8633 4213 8647 4227
rect 8693 4213 8707 4227
rect 8593 4193 8607 4207
rect 8593 4073 8607 4087
rect 8613 4053 8627 4067
rect 8653 4153 8667 4167
rect 8633 3893 8647 3907
rect 8713 4093 8727 4107
rect 8793 4213 8807 4227
rect 8733 4053 8747 4067
rect 8753 4034 8767 4048
rect 8813 4034 8827 4048
rect 8853 4034 8867 4048
rect 8693 3992 8707 4006
rect 8733 3992 8747 4006
rect 8793 3992 8807 4006
rect 8653 3873 8667 3887
rect 8953 5074 8967 5088
rect 8993 5074 9007 5088
rect 9033 5074 9047 5088
rect 9073 5052 9087 5066
rect 9153 5313 9167 5327
rect 9433 5973 9447 5987
rect 9473 5833 9487 5847
rect 9353 5653 9367 5667
rect 9333 5553 9347 5567
rect 9533 6433 9547 6447
rect 9573 6453 9587 6467
rect 9553 6233 9567 6247
rect 9533 6173 9547 6187
rect 9573 5973 9587 5987
rect 9533 5873 9547 5887
rect 9513 5733 9527 5747
rect 9453 5613 9467 5627
rect 9493 5613 9507 5627
rect 9413 5594 9427 5608
rect 9393 5552 9407 5566
rect 9353 5513 9367 5527
rect 9493 5552 9507 5566
rect 9433 5513 9447 5527
rect 9413 5473 9427 5487
rect 9633 6693 9647 6707
rect 9613 6633 9627 6647
rect 9613 6453 9627 6467
rect 9733 7273 9747 7287
rect 9833 7392 9847 7406
rect 9873 7373 9887 7387
rect 9853 7333 9867 7347
rect 9793 7313 9807 7327
rect 9853 7273 9867 7287
rect 9773 7253 9787 7267
rect 9813 7213 9827 7227
rect 9773 7173 9787 7187
rect 9753 7154 9767 7168
rect 9713 7093 9727 7107
rect 9773 7093 9787 7107
rect 9733 7053 9747 7067
rect 9853 7173 9867 7187
rect 9773 6973 9787 6987
rect 9813 6973 9827 6987
rect 9973 7433 9987 7447
rect 10193 7593 10207 7607
rect 10213 7533 10227 7547
rect 10173 7453 10187 7467
rect 10393 7673 10407 7687
rect 10333 7632 10347 7646
rect 10293 7573 10307 7587
rect 10373 7533 10387 7547
rect 10293 7513 10307 7527
rect 10253 7473 10267 7487
rect 10133 7373 10147 7387
rect 10293 7453 10307 7467
rect 10253 7373 10267 7387
rect 10253 7333 10267 7347
rect 10093 7293 10107 7307
rect 10193 7293 10207 7307
rect 9913 7252 9927 7266
rect 10033 7213 10047 7227
rect 9913 7173 9927 7187
rect 9933 7153 9947 7167
rect 9953 7173 9967 7187
rect 10033 7153 10047 7167
rect 10653 8273 10667 8287
rect 10753 8273 10767 8287
rect 10553 8013 10567 8027
rect 10593 8013 10607 8027
rect 10532 7954 10546 7968
rect 10553 7953 10567 7967
rect 10573 7912 10587 7926
rect 10593 7813 10607 7827
rect 10633 8233 10647 8247
rect 10673 8213 10687 8227
rect 10713 8194 10727 8208
rect 10793 8253 10807 8267
rect 10873 8233 10887 8247
rect 10832 8172 10846 8186
rect 10853 8173 10867 8187
rect 10693 8152 10707 8166
rect 10733 8152 10747 8166
rect 10673 8113 10687 8127
rect 10653 7953 10667 7967
rect 10653 7913 10667 7927
rect 10633 7853 10647 7867
rect 10473 7633 10487 7647
rect 10453 7553 10467 7567
rect 10612 7673 10626 7687
rect 10633 7674 10647 7688
rect 10533 7573 10547 7587
rect 10493 7533 10507 7547
rect 10453 7473 10467 7487
rect 10533 7473 10547 7487
rect 10393 7353 10407 7367
rect 10293 7213 10307 7227
rect 10153 7193 10167 7207
rect 9913 7093 9927 7107
rect 10013 7112 10027 7126
rect 10053 7073 10067 7087
rect 9973 7013 9987 7027
rect 10253 7013 10267 7027
rect 10313 7013 10327 7027
rect 10133 6973 10147 6987
rect 9873 6933 9887 6947
rect 9853 6913 9867 6927
rect 9753 6833 9767 6847
rect 9713 6693 9727 6707
rect 9713 6672 9727 6686
rect 9693 6653 9707 6667
rect 9673 6634 9687 6648
rect 9753 6653 9767 6667
rect 9653 6592 9667 6606
rect 9693 6553 9707 6567
rect 9653 6513 9667 6527
rect 9713 6473 9727 6487
rect 9693 6414 9707 6428
rect 9613 6353 9627 6367
rect 9733 6333 9747 6347
rect 9633 6153 9647 6167
rect 9713 6153 9727 6167
rect 9673 6133 9687 6147
rect 9613 6072 9627 6086
rect 9653 6072 9667 6086
rect 9693 6072 9707 6086
rect 9733 6073 9747 6087
rect 9653 6033 9667 6047
rect 9692 6033 9706 6047
rect 9713 6033 9727 6047
rect 9673 6013 9687 6027
rect 9673 5933 9687 5947
rect 9693 5913 9707 5927
rect 9713 5874 9727 5888
rect 9673 5852 9687 5866
rect 9633 5813 9647 5827
rect 9593 5713 9607 5727
rect 9593 5673 9607 5687
rect 9633 5653 9647 5667
rect 9713 5653 9727 5667
rect 9653 5594 9667 5608
rect 9633 5552 9647 5566
rect 9573 5513 9587 5527
rect 9673 5513 9687 5527
rect 9713 5513 9727 5527
rect 9813 6813 9827 6827
rect 9793 6634 9807 6648
rect 9853 6873 9867 6887
rect 9833 6733 9847 6747
rect 9993 6912 10007 6926
rect 10033 6793 10047 6807
rect 9913 6673 9927 6687
rect 10013 6653 10027 6667
rect 9813 6593 9827 6607
rect 9793 6473 9807 6487
rect 9793 6413 9807 6427
rect 9773 6313 9787 6327
rect 9813 6313 9827 6327
rect 9773 6273 9787 6287
rect 9813 6133 9827 6147
rect 9773 6093 9787 6107
rect 9793 5773 9807 5787
rect 9513 5433 9527 5447
rect 9533 5413 9547 5427
rect 9513 5354 9527 5368
rect 9313 5293 9327 5307
rect 9253 5273 9267 5287
rect 9613 5353 9627 5367
rect 9413 5293 9427 5307
rect 9373 5233 9387 5247
rect 8973 5033 8987 5047
rect 9013 5032 9027 5046
rect 9173 5054 9187 5068
rect 9313 5054 9327 5068
rect 8953 5013 8967 5027
rect 9093 5013 9107 5027
rect 9133 5013 9147 5027
rect 9033 4913 9047 4927
rect 8933 4854 8947 4868
rect 8993 4853 9007 4867
rect 8893 4793 8907 4807
rect 8953 4793 8967 4807
rect 9053 4834 9067 4848
rect 8893 4673 8907 4687
rect 8973 4653 8987 4667
rect 8993 4593 9007 4607
rect 8933 4533 8947 4547
rect 8893 4493 8907 4507
rect 8933 4393 8947 4407
rect 9013 4433 9027 4447
rect 8973 4334 8987 4348
rect 8893 4233 8907 4247
rect 8873 3972 8887 3986
rect 8853 3913 8867 3927
rect 8813 3853 8827 3867
rect 8613 3814 8627 3828
rect 8553 3533 8567 3547
rect 8653 3772 8667 3786
rect 8813 3772 8827 3786
rect 8813 3733 8827 3747
rect 8833 3713 8847 3727
rect 8853 3693 8867 3707
rect 8833 3633 8847 3647
rect 8513 3492 8527 3506
rect 8453 3453 8467 3467
rect 8513 3413 8527 3427
rect 8493 3393 8507 3407
rect 8493 3353 8507 3367
rect 8413 3333 8427 3347
rect 8453 3313 8467 3327
rect 8553 3393 8567 3407
rect 8553 3313 8567 3327
rect 8513 3274 8527 3288
rect 8593 3494 8607 3508
rect 8373 3073 8387 3087
rect 8473 3252 8487 3266
rect 8513 3213 8527 3227
rect 8433 3173 8447 3187
rect 8453 3113 8467 3127
rect 8353 3053 8367 3067
rect 8413 3053 8427 3067
rect 8413 2972 8427 2986
rect 8333 2952 8347 2966
rect 8373 2952 8387 2966
rect 8453 2953 8467 2967
rect 8353 2913 8367 2927
rect 8353 2873 8367 2887
rect 8333 2853 8347 2867
rect 8453 2853 8467 2867
rect 8273 2774 8287 2788
rect 8593 3273 8607 3287
rect 8753 3494 8767 3508
rect 8913 4213 8927 4227
rect 8953 4193 8967 4207
rect 9033 4253 9047 4267
rect 8973 4173 8987 4187
rect 8933 4034 8947 4048
rect 8973 4034 8987 4048
rect 8953 3992 8967 4006
rect 8973 3893 8987 3907
rect 8933 3853 8947 3867
rect 8933 3733 8947 3747
rect 8913 3693 8927 3707
rect 8913 3633 8927 3647
rect 8893 3533 8907 3547
rect 8953 3533 8967 3547
rect 8873 3492 8887 3506
rect 8853 3313 8867 3327
rect 8773 3273 8787 3287
rect 8753 3253 8767 3267
rect 8553 3113 8567 3127
rect 8613 3113 8627 3127
rect 8653 2974 8667 2988
rect 8973 3453 8987 3467
rect 8973 3313 8987 3327
rect 8953 3253 8967 3267
rect 8893 3233 8907 3247
rect 9013 3673 9027 3687
rect 9013 3593 9027 3607
rect 9013 3572 9027 3586
rect 9013 3453 9027 3467
rect 9013 3432 9027 3446
rect 8813 3053 8827 3067
rect 8773 2972 8787 2986
rect 8853 2973 8867 2987
rect 8913 3113 8927 3127
rect 8893 2893 8907 2907
rect 8993 3233 9007 3247
rect 8993 3193 9007 3207
rect 8973 3173 8987 3187
rect 8953 3132 8967 3146
rect 8933 3093 8947 3107
rect 8473 2833 8487 2847
rect 8453 2813 8467 2827
rect 8373 2774 8387 2788
rect 8453 2773 8467 2787
rect 8313 2732 8327 2746
rect 8253 2693 8267 2707
rect 8253 2653 8267 2667
rect 8233 2553 8247 2567
rect 8353 2673 8367 2687
rect 8333 2553 8347 2567
rect 8313 2532 8327 2546
rect 8233 2452 8247 2466
rect 8213 2413 8227 2427
rect 8273 2413 8287 2427
rect 8253 2373 8267 2387
rect 7993 2353 8007 2367
rect 8233 2333 8247 2347
rect 8033 2313 8047 2327
rect 8093 2313 8107 2327
rect 8013 2293 8027 2307
rect 8013 2272 8027 2286
rect 8053 2273 8067 2287
rect 8173 2293 8187 2307
rect 8133 2254 8147 2268
rect 8213 2233 8227 2247
rect 8253 2233 8267 2247
rect 8013 2213 8027 2227
rect 7993 2173 8007 2187
rect 8113 2212 8127 2226
rect 8173 2113 8187 2127
rect 8073 2013 8087 2027
rect 8133 2013 8147 2027
rect 8093 1993 8107 2007
rect 8053 1973 8067 1987
rect 8033 1893 8047 1907
rect 7993 1833 8007 1847
rect 7713 1753 7727 1767
rect 7653 1733 7667 1747
rect 7593 1692 7607 1706
rect 7553 1653 7567 1667
rect 7573 1633 7587 1647
rect 7653 1633 7667 1647
rect 7553 1593 7567 1607
rect 7513 1493 7527 1507
rect 7813 1712 7827 1726
rect 7793 1553 7807 1567
rect 7573 1473 7587 1487
rect 7493 1453 7507 1467
rect 7873 1493 7887 1507
rect 7613 1434 7627 1448
rect 7653 1434 7667 1448
rect 7753 1434 7767 1448
rect 7793 1434 7807 1448
rect 7833 1434 7847 1448
rect 7493 1393 7507 1407
rect 7633 1392 7647 1406
rect 7653 1214 7667 1228
rect 7433 1172 7447 1186
rect 7493 1172 7507 1186
rect 7633 1172 7647 1186
rect 7673 1172 7687 1186
rect 7513 1153 7527 1167
rect 7453 1033 7467 1047
rect 7293 833 7307 847
rect 7293 793 7307 807
rect 7233 753 7247 767
rect 7193 393 7207 407
rect 7193 313 7207 327
rect 7473 872 7487 886
rect 7433 813 7447 827
rect 7313 753 7327 767
rect 7333 694 7347 708
rect 7353 633 7367 647
rect 7553 1073 7567 1087
rect 7533 913 7547 927
rect 7533 872 7547 886
rect 7513 713 7527 727
rect 7453 694 7467 708
rect 7693 973 7707 987
rect 7673 872 7687 886
rect 7593 694 7607 708
rect 7533 652 7547 666
rect 7432 613 7446 627
rect 7453 613 7467 627
rect 7353 513 7367 527
rect 7573 513 7587 527
rect 7613 513 7627 527
rect 7533 493 7547 507
rect 7313 473 7327 487
rect 7353 473 7367 487
rect 7333 394 7347 408
rect 7393 393 7407 407
rect 7573 394 7587 408
rect 7393 352 7407 366
rect 7553 352 7567 366
rect 7613 353 7627 367
rect 7773 1053 7787 1067
rect 7973 1793 7987 1807
rect 8053 1753 8067 1767
rect 8113 1893 8127 1907
rect 8113 1853 8127 1867
rect 8153 1933 8167 1947
rect 8133 1673 8147 1687
rect 8153 1613 8167 1627
rect 8113 1473 8127 1487
rect 8013 1433 8027 1447
rect 7893 1392 7907 1406
rect 7953 1392 7967 1406
rect 8013 1353 8027 1367
rect 7853 1313 7867 1327
rect 7813 1253 7827 1267
rect 7813 1013 7827 1027
rect 7793 973 7807 987
rect 7873 993 7887 1007
rect 7953 1213 7967 1227
rect 7993 1213 8007 1227
rect 7893 953 7907 967
rect 7913 933 7927 947
rect 7953 933 7967 947
rect 7873 914 7887 928
rect 7813 873 7827 887
rect 7853 813 7867 827
rect 7773 753 7787 767
rect 7953 873 7967 887
rect 7973 853 7987 867
rect 7893 793 7907 807
rect 7933 793 7947 807
rect 7893 753 7907 767
rect 7833 694 7847 708
rect 7913 653 7927 667
rect 7793 613 7807 627
rect 7753 553 7767 567
rect 7893 553 7907 567
rect 7813 433 7827 447
rect 7753 394 7767 408
rect 7673 352 7687 366
rect 7733 352 7747 366
rect 7773 352 7787 366
rect 7813 352 7827 366
rect 7353 313 7367 327
rect 7673 313 7687 327
rect 7853 313 7867 327
rect 7433 253 7447 267
rect 7313 213 7327 227
rect 7233 174 7247 188
rect 7313 173 7327 187
rect 8073 1433 8087 1447
rect 8113 1434 8127 1448
rect 8133 1392 8147 1406
rect 8133 1373 8147 1387
rect 8133 1333 8147 1347
rect 8053 1273 8067 1287
rect 8093 1273 8107 1287
rect 8033 1214 8047 1228
rect 8093 1214 8107 1228
rect 8013 1172 8027 1186
rect 8033 953 8047 967
rect 8133 1093 8147 1107
rect 8133 953 8147 967
rect 8033 793 8047 807
rect 7993 773 8007 787
rect 7953 653 7967 667
rect 7953 593 7967 607
rect 7953 493 7967 507
rect 7933 473 7947 487
rect 8113 872 8127 886
rect 8153 873 8167 887
rect 8153 833 8167 847
rect 8353 2493 8367 2507
rect 8333 2373 8347 2387
rect 8533 2873 8547 2887
rect 8573 2873 8587 2887
rect 8753 2873 8767 2887
rect 8913 2873 8927 2887
rect 8613 2813 8627 2827
rect 8493 2733 8507 2747
rect 8553 2732 8567 2746
rect 8553 2673 8567 2687
rect 8473 2512 8487 2526
rect 8553 2453 8567 2467
rect 8513 2413 8527 2427
rect 8493 2373 8507 2387
rect 8313 2333 8327 2347
rect 8433 2333 8447 2347
rect 8413 2173 8427 2187
rect 8653 2653 8667 2667
rect 8633 2553 8647 2567
rect 8613 2474 8627 2488
rect 8593 2413 8607 2427
rect 8573 2192 8587 2206
rect 8513 2133 8527 2147
rect 8273 2113 8287 2127
rect 8553 2113 8567 2127
rect 8553 2053 8567 2067
rect 8573 2033 8587 2047
rect 8213 2013 8227 2027
rect 8493 2013 8507 2027
rect 8233 1993 8247 2007
rect 8213 1973 8227 1987
rect 8293 1954 8307 1968
rect 8453 1954 8467 1968
rect 8573 1993 8587 2007
rect 8553 1973 8567 1987
rect 8233 1912 8247 1926
rect 8273 1912 8287 1926
rect 8473 1912 8487 1926
rect 8553 1873 8567 1887
rect 8293 1853 8307 1867
rect 8513 1853 8527 1867
rect 8213 1734 8227 1748
rect 8253 1734 8267 1748
rect 8493 1734 8507 1748
rect 8573 1773 8587 1787
rect 8193 1613 8207 1627
rect 8213 1593 8227 1607
rect 8413 1673 8427 1687
rect 8273 1553 8287 1567
rect 8233 1473 8247 1487
rect 8313 1434 8327 1448
rect 8273 1392 8287 1406
rect 8333 1373 8347 1387
rect 8273 1273 8287 1287
rect 8393 1273 8407 1287
rect 8233 1173 8247 1187
rect 8293 1172 8307 1186
rect 8373 1013 8387 1027
rect 8213 953 8227 967
rect 8333 914 8347 928
rect 8353 872 8367 886
rect 8313 853 8327 867
rect 8193 813 8207 827
rect 8173 713 8187 727
rect 8113 694 8127 708
rect 8173 673 8187 687
rect 8053 652 8067 666
rect 8093 652 8107 666
rect 8033 613 8047 627
rect 7993 433 8007 447
rect 7993 394 8007 408
rect 7913 353 7927 367
rect 7973 352 7987 366
rect 7913 293 7927 307
rect 7933 233 7947 247
rect 7913 213 7927 227
rect 7473 174 7487 188
rect 7513 174 7527 188
rect 7653 174 7667 188
rect 7853 174 7867 188
rect 7893 174 7907 188
rect 7173 132 7187 146
rect 7253 132 7267 146
rect 7093 53 7107 67
rect 7453 53 7467 67
rect 7633 132 7647 146
rect 7833 133 7847 147
rect 7873 132 7887 146
rect 7933 133 7947 147
rect 8093 593 8107 607
rect 8052 533 8066 547
rect 8073 533 8087 547
rect 8113 433 8127 447
rect 8113 352 8127 366
rect 8173 593 8187 607
rect 8173 493 8187 507
rect 8313 713 8327 727
rect 8353 694 8367 708
rect 8513 1692 8527 1706
rect 8593 1733 8607 1747
rect 8573 1653 8587 1667
rect 8413 693 8427 707
rect 8553 1453 8567 1467
rect 8713 2593 8727 2607
rect 8733 2593 8747 2607
rect 8793 2533 8807 2547
rect 8773 2493 8787 2507
rect 8693 2474 8707 2488
rect 8653 2192 8667 2206
rect 8633 2153 8647 2167
rect 8653 2053 8667 2067
rect 8713 2413 8727 2427
rect 8733 2313 8747 2327
rect 8693 2273 8707 2287
rect 8693 2113 8707 2127
rect 8633 2013 8647 2027
rect 8673 2013 8687 2027
rect 8613 1593 8627 1607
rect 8673 1954 8687 1968
rect 8873 2613 8887 2627
rect 8813 2393 8827 2407
rect 8793 2273 8807 2287
rect 8813 2254 8827 2268
rect 8913 2573 8927 2587
rect 9173 4993 9187 5007
rect 9533 5313 9547 5327
rect 9633 5313 9647 5327
rect 9473 5273 9487 5287
rect 9653 5233 9667 5247
rect 9473 5094 9487 5108
rect 9433 5052 9447 5066
rect 9513 5053 9527 5067
rect 9713 5094 9727 5108
rect 9473 4933 9487 4947
rect 9413 4913 9427 4927
rect 9433 4873 9447 4887
rect 9193 4693 9207 4707
rect 9233 4693 9247 4707
rect 9273 4693 9287 4707
rect 9133 4653 9147 4667
rect 9233 4554 9247 4568
rect 9393 4753 9407 4767
rect 9293 4554 9307 4568
rect 9453 4834 9467 4848
rect 9473 4813 9487 4827
rect 9453 4793 9467 4807
rect 9593 4753 9607 4767
rect 9613 4713 9627 4727
rect 9513 4653 9527 4667
rect 9453 4593 9467 4607
rect 9133 4512 9147 4526
rect 9173 4512 9187 4526
rect 9213 4512 9227 4526
rect 9273 4513 9287 4527
rect 9233 4433 9247 4447
rect 9093 4393 9107 4407
rect 9113 4373 9127 4387
rect 9153 4334 9167 4348
rect 9133 4292 9147 4306
rect 9133 4034 9147 4048
rect 9173 4034 9187 4048
rect 9193 3953 9207 3967
rect 9153 3913 9167 3927
rect 9173 3873 9187 3887
rect 9113 3814 9127 3828
rect 9133 3772 9147 3786
rect 9073 3693 9087 3707
rect 9133 3733 9147 3747
rect 9053 3633 9067 3647
rect 9053 3493 9067 3507
rect 9053 3393 9067 3407
rect 9093 3513 9107 3527
rect 9273 4073 9287 4087
rect 9253 4034 9267 4048
rect 9273 3993 9287 4007
rect 9273 3813 9287 3827
rect 9473 4512 9487 4526
rect 9433 4473 9447 4487
rect 9413 4373 9427 4387
rect 9473 4373 9487 4387
rect 9373 4334 9387 4348
rect 9393 4292 9407 4306
rect 9333 4233 9347 4247
rect 9473 4334 9487 4348
rect 9413 4213 9427 4227
rect 9393 4073 9407 4087
rect 9433 4034 9447 4048
rect 9333 3993 9347 4007
rect 9373 3992 9387 4006
rect 9413 3873 9427 3887
rect 9553 4433 9567 4447
rect 9693 4673 9707 4687
rect 9653 4554 9667 4568
rect 9953 6634 9967 6648
rect 9893 6592 9907 6606
rect 9933 6592 9947 6606
rect 10012 6593 10026 6607
rect 10173 6953 10187 6967
rect 10233 6914 10247 6928
rect 10273 6953 10287 6967
rect 10293 6913 10307 6927
rect 10273 6853 10287 6867
rect 10293 6833 10307 6847
rect 10453 7193 10467 7207
rect 10433 7173 10447 7187
rect 10433 7133 10447 7147
rect 10413 7073 10427 7087
rect 10333 6973 10347 6987
rect 10393 6973 10407 6987
rect 10313 6813 10327 6827
rect 10253 6793 10267 6807
rect 10153 6773 10167 6787
rect 10133 6733 10147 6747
rect 10273 6733 10287 6747
rect 10193 6653 10207 6667
rect 10273 6654 10287 6668
rect 10073 6613 10087 6627
rect 10033 6592 10047 6606
rect 10033 6553 10047 6567
rect 9973 6473 9987 6487
rect 9893 6453 9907 6467
rect 9933 6414 9947 6428
rect 10013 6453 10027 6467
rect 9873 6353 9887 6367
rect 9893 6313 9907 6327
rect 9853 6173 9867 6187
rect 9833 6113 9847 6127
rect 9893 6153 9907 6167
rect 9973 6133 9987 6147
rect 9913 6072 9927 6086
rect 10233 6612 10247 6626
rect 10273 6614 10287 6628
rect 10133 6592 10147 6606
rect 10173 6533 10187 6547
rect 10272 6533 10286 6547
rect 10293 6533 10307 6547
rect 10573 7553 10587 7567
rect 10633 7473 10647 7487
rect 10693 8093 10707 8107
rect 10773 8093 10787 8107
rect 10713 8073 10727 8087
rect 10853 8073 10867 8087
rect 10693 8013 10707 8027
rect 10693 7813 10707 7827
rect 10693 7753 10707 7767
rect 11013 8972 11027 8986
rect 11073 8953 11087 8967
rect 11173 9013 11187 9027
rect 11153 8953 11167 8967
rect 11113 8873 11127 8887
rect 11173 8833 11187 8847
rect 11273 9733 11287 9747
rect 11273 9593 11287 9607
rect 11253 9453 11267 9467
rect 11273 9333 11287 9347
rect 11253 9193 11267 9207
rect 11313 9133 11327 9147
rect 11093 8694 11107 8708
rect 11133 8593 11147 8607
rect 11053 8573 11067 8587
rect 11053 8494 11067 8508
rect 11093 8494 11107 8508
rect 10913 8213 10927 8227
rect 10913 8173 10927 8187
rect 10893 8113 10907 8127
rect 11113 8313 11127 8327
rect 11253 8734 11267 8748
rect 11293 8734 11307 8748
rect 11213 8692 11227 8706
rect 11313 8693 11327 8707
rect 11233 8673 11247 8687
rect 11293 8673 11307 8687
rect 11293 8652 11307 8666
rect 11333 8653 11347 8667
rect 11073 8213 11087 8227
rect 11073 8174 11087 8188
rect 10933 8133 10947 8147
rect 10913 8093 10927 8107
rect 10893 8073 10907 8087
rect 10873 8033 10887 8047
rect 10773 7993 10787 8007
rect 10873 7993 10887 8007
rect 10813 7974 10827 7988
rect 10793 7932 10807 7946
rect 10833 7913 10847 7927
rect 10813 7833 10827 7847
rect 10733 7674 10747 7688
rect 10873 7793 10887 7807
rect 10933 8033 10947 8047
rect 10813 7673 10827 7687
rect 10833 7652 10847 7666
rect 10693 7632 10707 7646
rect 10673 7593 10687 7607
rect 10673 7513 10687 7527
rect 10753 7632 10767 7646
rect 10673 7353 10687 7367
rect 10713 7353 10727 7367
rect 10593 7313 10607 7327
rect 10753 7313 10767 7327
rect 10913 7654 10927 7668
rect 10893 7593 10907 7607
rect 10873 7553 10887 7567
rect 10893 7533 10907 7547
rect 10833 7513 10847 7527
rect 10893 7512 10907 7526
rect 10853 7473 10867 7487
rect 10873 7393 10887 7407
rect 10753 7273 10767 7287
rect 10793 7273 10807 7287
rect 10613 7253 10627 7267
rect 10593 7173 10607 7187
rect 10493 7113 10507 7127
rect 10533 7113 10547 7127
rect 10493 7013 10507 7027
rect 10453 6973 10467 6987
rect 10393 6952 10407 6966
rect 10433 6953 10447 6967
rect 10533 6913 10547 6927
rect 10393 6892 10407 6906
rect 10433 6892 10447 6906
rect 10593 7133 10607 7147
rect 10593 6993 10607 7007
rect 10593 6972 10607 6986
rect 10593 6892 10607 6906
rect 10573 6853 10587 6867
rect 10573 6773 10587 6787
rect 10473 6693 10487 6707
rect 10473 6614 10487 6628
rect 10493 6513 10507 6527
rect 11053 7993 11067 8007
rect 11013 7974 11027 7988
rect 11033 7873 11047 7887
rect 11073 7833 11087 7847
rect 11073 7654 11087 7668
rect 10953 7553 10967 7567
rect 10893 7073 10907 7087
rect 10713 6993 10727 7007
rect 10753 6993 10767 7007
rect 10853 6993 10867 7007
rect 10673 6934 10687 6948
rect 10653 6892 10667 6906
rect 10733 6893 10747 6907
rect 10693 6773 10707 6787
rect 10613 6733 10627 6747
rect 10633 6654 10647 6668
rect 10693 6733 10707 6747
rect 10593 6612 10607 6626
rect 10673 6613 10687 6627
rect 10593 6553 10607 6567
rect 10473 6473 10487 6487
rect 10213 6392 10227 6406
rect 10213 6313 10227 6327
rect 10173 6273 10187 6287
rect 10073 6193 10087 6207
rect 10133 6133 10147 6147
rect 10053 6114 10067 6128
rect 10093 6114 10107 6128
rect 10193 6153 10207 6167
rect 10173 6113 10187 6127
rect 10033 6073 10047 6087
rect 9973 6033 9987 6047
rect 10013 6033 10027 6047
rect 10153 6033 10167 6047
rect 10113 5913 10127 5927
rect 10053 5894 10067 5908
rect 9953 5872 9967 5886
rect 9813 5753 9827 5767
rect 9973 5753 9987 5767
rect 9953 5693 9967 5707
rect 9873 5633 9887 5647
rect 9913 5613 9927 5627
rect 9893 5533 9907 5547
rect 9913 5513 9927 5527
rect 9853 5413 9867 5427
rect 9793 5373 9807 5387
rect 9813 5273 9827 5287
rect 9793 4893 9807 4907
rect 9613 4513 9627 4527
rect 9673 4512 9687 4526
rect 9693 4413 9707 4427
rect 9593 4393 9607 4407
rect 9673 4393 9687 4407
rect 9593 4372 9607 4386
rect 9513 4293 9527 4307
rect 9613 4292 9627 4306
rect 9573 4233 9587 4247
rect 9553 4093 9567 4107
rect 9413 3852 9427 3866
rect 9473 3853 9487 3867
rect 9333 3814 9347 3828
rect 9373 3814 9387 3828
rect 9333 3773 9347 3787
rect 9273 3753 9287 3767
rect 9253 3693 9267 3707
rect 9393 3753 9407 3767
rect 9433 3713 9447 3727
rect 9353 3673 9367 3687
rect 9493 3673 9507 3687
rect 9253 3633 9267 3647
rect 9233 3553 9247 3567
rect 9213 3493 9227 3507
rect 9353 3573 9367 3587
rect 9333 3553 9347 3567
rect 9333 3493 9347 3507
rect 9093 3433 9107 3447
rect 9113 3413 9127 3427
rect 9153 3413 9167 3427
rect 9253 3453 9267 3467
rect 9133 3294 9147 3308
rect 9173 3294 9187 3308
rect 9213 3292 9227 3306
rect 9073 3233 9087 3247
rect 9173 3233 9187 3247
rect 9153 3212 9167 3226
rect 9033 3173 9047 3187
rect 9113 3173 9127 3187
rect 9013 3053 9027 3067
rect 8973 2993 8987 3007
rect 9013 2994 9027 3008
rect 9053 2952 9067 2966
rect 9053 2853 9067 2867
rect 8993 2833 9007 2847
rect 8973 2753 8987 2767
rect 9013 2813 9027 2827
rect 9053 2773 9067 2787
rect 9053 2754 9067 2768
rect 9013 2733 9027 2747
rect 9033 2713 9047 2727
rect 9033 2533 9047 2547
rect 9093 3053 9107 3067
rect 9093 2533 9107 2547
rect 9033 2493 9047 2507
rect 8953 2473 8967 2487
rect 8893 2433 8907 2447
rect 8973 2432 8987 2446
rect 8933 2393 8947 2407
rect 9033 2453 9047 2467
rect 9013 2353 9027 2367
rect 8933 2313 8947 2327
rect 8893 2173 8907 2187
rect 8913 2133 8927 2147
rect 8813 2013 8827 2027
rect 8753 1954 8767 1968
rect 8653 1913 8667 1927
rect 8693 1893 8707 1907
rect 8733 1893 8747 1907
rect 8653 1753 8667 1767
rect 8753 1833 8767 1847
rect 8733 1734 8747 1748
rect 8793 1733 8807 1747
rect 8753 1673 8767 1687
rect 8713 1633 8727 1647
rect 8833 1954 8847 1968
rect 8813 1673 8827 1687
rect 8753 1613 8767 1627
rect 8793 1613 8807 1627
rect 8633 1553 8647 1567
rect 8733 1533 8747 1547
rect 8673 1453 8687 1467
rect 8653 1413 8667 1427
rect 8533 1233 8547 1247
rect 8493 1214 8507 1228
rect 8513 1172 8527 1186
rect 8613 1392 8627 1406
rect 8673 1393 8687 1407
rect 8652 1353 8666 1367
rect 8673 1353 8687 1367
rect 8613 1233 8627 1247
rect 8713 1273 8727 1287
rect 8713 1234 8727 1248
rect 8793 1573 8807 1587
rect 8973 2273 8987 2287
rect 9013 2273 9027 2287
rect 8953 2253 8967 2267
rect 9133 3013 9147 3027
rect 9133 2953 9147 2967
rect 9133 2893 9147 2907
rect 9133 2793 9147 2807
rect 9273 3333 9287 3347
rect 9253 3252 9267 3266
rect 9213 3213 9227 3227
rect 9193 3193 9207 3207
rect 9233 3013 9247 3027
rect 9193 2993 9207 3007
rect 9413 3313 9427 3327
rect 9293 3293 9307 3307
rect 9373 3294 9387 3308
rect 9353 3252 9367 3266
rect 9513 3493 9527 3507
rect 9533 3473 9547 3487
rect 9513 3253 9527 3267
rect 9513 3133 9527 3147
rect 9493 3093 9507 3107
rect 9513 3073 9527 3087
rect 9633 4253 9647 4267
rect 9633 4213 9647 4227
rect 9613 4054 9627 4068
rect 9633 3973 9647 3987
rect 9593 3953 9607 3967
rect 9633 3814 9647 3828
rect 9673 3772 9687 3786
rect 9613 3753 9627 3767
rect 9613 3713 9627 3727
rect 9613 3514 9627 3528
rect 9633 3473 9647 3487
rect 9673 3413 9687 3427
rect 9573 3373 9587 3387
rect 9633 3353 9647 3367
rect 9653 3333 9667 3347
rect 9573 3313 9587 3327
rect 9613 3294 9627 3308
rect 9593 3252 9607 3266
rect 9613 3213 9627 3227
rect 9633 3193 9647 3207
rect 9593 3113 9607 3127
rect 9553 3093 9567 3107
rect 9373 3033 9387 3047
rect 9533 3033 9547 3047
rect 9273 2993 9287 3007
rect 9213 2952 9227 2966
rect 9253 2952 9267 2966
rect 9313 2973 9327 2987
rect 9293 2933 9307 2947
rect 9173 2913 9187 2927
rect 9273 2913 9287 2927
rect 9213 2873 9227 2887
rect 9173 2853 9187 2867
rect 9153 2753 9167 2767
rect 9133 2613 9147 2627
rect 9193 2573 9207 2587
rect 9173 2553 9187 2567
rect 9313 2893 9327 2907
rect 9233 2713 9247 2727
rect 9253 2713 9267 2727
rect 9213 2513 9227 2527
rect 9293 2673 9307 2687
rect 9293 2573 9307 2587
rect 9273 2553 9287 2567
rect 9273 2453 9287 2467
rect 9353 2972 9367 2986
rect 9393 2974 9407 2988
rect 9533 2974 9547 2988
rect 9673 3153 9687 3167
rect 9673 3093 9687 3107
rect 9733 4353 9747 4367
rect 9713 4213 9727 4227
rect 9713 4033 9727 4047
rect 9713 3493 9727 3507
rect 9733 3413 9747 3427
rect 9733 3373 9747 3387
rect 9713 3293 9727 3307
rect 9693 3053 9707 3067
rect 9713 3013 9727 3027
rect 9653 2972 9667 2986
rect 9633 2913 9647 2927
rect 9573 2873 9587 2887
rect 9413 2853 9427 2867
rect 9533 2833 9547 2847
rect 9493 2774 9507 2788
rect 9473 2732 9487 2746
rect 9413 2633 9427 2647
rect 9393 2613 9407 2627
rect 9413 2474 9427 2488
rect 9173 2432 9187 2446
rect 9213 2432 9227 2446
rect 9293 2432 9307 2446
rect 9333 2432 9347 2446
rect 9393 2432 9407 2446
rect 9113 2413 9127 2427
rect 9193 2373 9207 2387
rect 9173 2353 9187 2367
rect 9073 2333 9087 2347
rect 9053 2313 9067 2327
rect 9173 2293 9187 2307
rect 9433 2413 9447 2427
rect 9453 2373 9467 2387
rect 9513 2373 9527 2387
rect 9393 2353 9407 2367
rect 9433 2353 9447 2367
rect 9193 2253 9207 2267
rect 8973 2212 8987 2226
rect 8953 2093 8967 2107
rect 8933 2033 8947 2047
rect 8953 1993 8967 2007
rect 8913 1954 8927 1968
rect 8953 1954 8967 1968
rect 8893 1913 8907 1927
rect 8853 1873 8867 1887
rect 8933 1912 8947 1926
rect 8973 1893 8987 1907
rect 8853 1693 8867 1707
rect 8792 1473 8806 1487
rect 8813 1473 8827 1487
rect 8833 1453 8847 1467
rect 8853 1393 8867 1407
rect 8813 1333 8827 1347
rect 8753 1253 8767 1267
rect 8833 1253 8847 1267
rect 8673 1214 8687 1228
rect 8713 1213 8727 1227
rect 8653 1172 8667 1186
rect 8573 1113 8587 1127
rect 8513 1053 8527 1067
rect 8473 993 8487 1007
rect 8453 953 8467 967
rect 8373 652 8387 666
rect 8413 652 8427 666
rect 8473 873 8487 887
rect 8453 633 8467 647
rect 8333 613 8347 627
rect 8293 493 8307 507
rect 8193 433 8207 447
rect 8173 352 8187 366
rect 8133 293 8147 307
rect 8113 253 8127 267
rect 8093 233 8107 247
rect 8213 233 8227 247
rect 8393 394 8407 408
rect 8373 293 8387 307
rect 8153 174 8167 188
rect 8073 113 8087 127
rect 8033 93 8047 107
rect 8433 253 8447 267
rect 8153 113 8167 127
rect 8413 113 8427 127
rect 8553 1013 8567 1027
rect 8733 1133 8747 1147
rect 8773 1133 8787 1147
rect 8693 1033 8707 1047
rect 8593 914 8607 928
rect 8652 914 8666 928
rect 8673 914 8687 928
rect 8573 872 8587 886
rect 8613 853 8627 867
rect 8593 793 8607 807
rect 8593 753 8607 767
rect 8633 793 8647 807
rect 8633 693 8647 707
rect 8613 613 8627 627
rect 8553 533 8567 547
rect 8573 473 8587 487
rect 8613 413 8627 427
rect 8653 393 8667 407
rect 8513 293 8527 307
rect 8633 352 8647 366
rect 8613 293 8627 307
rect 8593 253 8607 267
rect 8493 233 8507 247
rect 8513 174 8527 188
rect 8433 93 8447 107
rect 8573 132 8587 146
rect 8533 53 8547 67
rect 7833 33 7847 47
rect 8113 33 8127 47
rect 8573 33 8587 47
rect 8713 973 8727 987
rect 8693 694 8707 708
rect 8673 313 8687 327
rect 8893 1734 8907 1748
rect 8933 1734 8947 1748
rect 8953 1692 8967 1706
rect 9013 2212 9027 2226
rect 9073 2193 9087 2207
rect 9013 2173 9027 2187
rect 9033 1954 9047 1968
rect 9013 1913 9027 1927
rect 9093 2153 9107 2167
rect 9293 2093 9307 2107
rect 9313 2073 9327 2087
rect 9133 2053 9147 2067
rect 9113 2033 9127 2047
rect 9313 2013 9327 2027
rect 9113 1993 9127 2007
rect 9253 1993 9267 2007
rect 9393 1993 9407 2007
rect 9193 1973 9207 1987
rect 9093 1954 9107 1968
rect 9153 1954 9167 1968
rect 9033 1893 9047 1907
rect 9133 1912 9147 1926
rect 9173 1893 9187 1907
rect 9233 1893 9247 1907
rect 9133 1853 9147 1867
rect 9213 1773 9227 1787
rect 9193 1753 9207 1767
rect 9173 1734 9187 1748
rect 9213 1733 9227 1747
rect 9373 1912 9387 1926
rect 9453 2293 9467 2307
rect 9493 2293 9507 2307
rect 9473 2253 9487 2267
rect 9453 2033 9467 2047
rect 9293 1853 9307 1867
rect 9433 1853 9447 1867
rect 9253 1793 9267 1807
rect 9273 1773 9287 1787
rect 9153 1692 9167 1706
rect 9093 1673 9107 1687
rect 9153 1673 9167 1687
rect 8993 1633 9007 1647
rect 9173 1633 9187 1647
rect 9133 1553 9147 1567
rect 8892 1533 8906 1547
rect 8913 1533 8927 1547
rect 9093 1533 9107 1547
rect 8893 1473 8907 1487
rect 8853 1213 8867 1227
rect 8853 1173 8867 1187
rect 8853 1133 8867 1147
rect 8913 1453 8927 1467
rect 8913 1413 8927 1427
rect 8973 1434 8987 1448
rect 9033 1434 9047 1448
rect 8953 1353 8967 1367
rect 9113 1433 9127 1447
rect 9053 1392 9067 1406
rect 9073 1373 9087 1387
rect 9013 1353 9027 1367
rect 8972 1333 8986 1347
rect 8993 1333 9007 1347
rect 9073 1333 9087 1347
rect 8913 1273 8927 1287
rect 9013 1273 9027 1287
rect 9053 1253 9067 1267
rect 8973 1233 8987 1247
rect 8853 1053 8867 1067
rect 8893 1053 8907 1067
rect 8833 1033 8847 1047
rect 8793 993 8807 1007
rect 8993 1013 9007 1027
rect 8833 933 8847 947
rect 8833 914 8847 928
rect 8953 913 8967 927
rect 9153 1533 9167 1547
rect 9153 1393 9167 1407
rect 9133 1333 9147 1347
rect 9273 1593 9287 1607
rect 9233 1473 9247 1487
rect 9313 1793 9327 1807
rect 9253 1434 9267 1448
rect 9293 1434 9307 1448
rect 9213 1393 9227 1407
rect 9133 1293 9147 1307
rect 9173 1293 9187 1307
rect 9113 993 9127 1007
rect 9093 913 9107 927
rect 8933 893 8947 907
rect 8733 873 8747 887
rect 8733 773 8747 787
rect 8813 853 8827 867
rect 8773 733 8787 747
rect 8773 694 8787 708
rect 8793 633 8807 647
rect 8753 553 8767 567
rect 8873 693 8887 707
rect 8953 833 8967 847
rect 8993 833 9007 847
rect 9093 853 9107 867
rect 8993 753 9007 767
rect 9033 753 9047 767
rect 9013 694 9027 708
rect 9033 652 9047 666
rect 9073 652 9087 666
rect 9113 653 9127 667
rect 8933 613 8947 627
rect 8993 613 9007 627
rect 8873 573 8887 587
rect 8853 493 8867 507
rect 8993 433 9007 447
rect 8793 394 8807 408
rect 8873 393 8887 407
rect 8953 394 8967 408
rect 9033 394 9047 408
rect 8753 353 8767 367
rect 8813 352 8827 366
rect 8733 333 8747 347
rect 8813 333 8827 347
rect 8853 333 8867 347
rect 8853 253 8867 267
rect 8713 193 8727 207
rect 8753 174 8767 188
rect 9013 352 9027 366
rect 8953 293 8967 307
rect 9253 1353 9267 1367
rect 9153 1214 9167 1228
rect 9213 1214 9227 1228
rect 9193 1172 9207 1186
rect 9233 1173 9247 1187
rect 9233 1033 9247 1047
rect 9173 1013 9187 1027
rect 9293 1214 9307 1228
rect 9293 1133 9307 1147
rect 9273 973 9287 987
rect 9193 873 9207 887
rect 9173 793 9187 807
rect 9213 853 9227 867
rect 9273 793 9287 807
rect 9193 753 9207 767
rect 9233 753 9247 767
rect 9173 694 9187 708
rect 9253 694 9267 708
rect 9333 1773 9347 1787
rect 9353 1734 9367 1748
rect 9393 1734 9407 1748
rect 9373 1692 9387 1706
rect 9373 1613 9387 1627
rect 9373 1592 9387 1606
rect 9413 1593 9427 1607
rect 9353 1493 9367 1507
rect 9333 1172 9347 1186
rect 9313 613 9327 627
rect 9253 533 9267 547
rect 9233 513 9247 527
rect 9173 493 9187 507
rect 9153 393 9167 407
rect 9293 493 9307 507
rect 9553 2774 9567 2788
rect 9553 2653 9567 2667
rect 9553 2473 9567 2487
rect 9773 4554 9787 4568
rect 9773 4513 9787 4527
rect 9873 5354 9887 5368
rect 9853 5233 9867 5247
rect 9833 5053 9847 5067
rect 9833 5013 9847 5027
rect 9813 4853 9827 4867
rect 9793 4413 9807 4427
rect 9793 4392 9807 4406
rect 9833 4812 9847 4826
rect 9833 4593 9847 4607
rect 9933 5374 9947 5388
rect 9933 5273 9947 5287
rect 9913 5173 9927 5187
rect 9993 5733 10007 5747
rect 9973 5293 9987 5307
rect 9953 5074 9967 5088
rect 9933 5032 9947 5046
rect 9893 4953 9907 4967
rect 9913 4933 9927 4947
rect 9913 4812 9927 4826
rect 10113 5832 10127 5846
rect 10013 5693 10027 5707
rect 10093 5633 10107 5647
rect 10173 5893 10187 5907
rect 10193 5852 10207 5866
rect 10133 5613 10147 5627
rect 10153 5593 10167 5607
rect 10033 5552 10047 5566
rect 10073 5552 10087 5566
rect 10113 5552 10127 5566
rect 10153 5552 10167 5566
rect 10113 5533 10127 5547
rect 10153 5433 10167 5447
rect 10093 5393 10107 5407
rect 10093 5374 10107 5388
rect 10133 5374 10147 5388
rect 10193 5552 10207 5566
rect 10193 5373 10207 5387
rect 10033 5333 10047 5347
rect 10073 5332 10087 5346
rect 10113 5293 10127 5307
rect 10073 5273 10087 5287
rect 10153 5273 10167 5287
rect 10033 5253 10047 5267
rect 10013 5233 10027 5247
rect 10013 5093 10027 5107
rect 10013 5032 10027 5046
rect 10013 4853 10027 4867
rect 10013 4813 10027 4827
rect 9953 4793 9967 4807
rect 9993 4793 10007 4807
rect 9933 4733 9947 4747
rect 9813 4353 9827 4367
rect 9853 4554 9867 4568
rect 9893 4554 9907 4568
rect 10013 4633 10027 4647
rect 9973 4554 9987 4568
rect 9853 4433 9867 4447
rect 9893 4393 9907 4407
rect 9873 4333 9887 4347
rect 9813 4292 9827 4306
rect 9853 4292 9867 4306
rect 9813 4253 9827 4267
rect 9833 4034 9847 4048
rect 9953 4512 9967 4526
rect 9933 4333 9947 4347
rect 9913 4293 9927 4307
rect 9853 3992 9867 4006
rect 9893 3992 9907 4006
rect 9773 3913 9787 3927
rect 9813 3813 9827 3827
rect 9893 3873 9907 3887
rect 10013 4453 10027 4467
rect 10053 5173 10067 5187
rect 10053 4913 10067 4927
rect 10273 6253 10287 6267
rect 10213 5253 10227 5267
rect 10193 5193 10207 5207
rect 10133 5093 10147 5107
rect 10093 5073 10107 5087
rect 10093 4993 10107 5007
rect 10253 6113 10267 6127
rect 10253 5813 10267 5827
rect 10253 5713 10267 5727
rect 10333 6394 10347 6408
rect 10433 6393 10447 6407
rect 10373 6352 10387 6366
rect 10373 6233 10387 6247
rect 10473 6153 10487 6167
rect 10313 6113 10327 6127
rect 10353 6114 10367 6128
rect 10393 6113 10407 6127
rect 10333 6072 10347 6086
rect 10353 5913 10367 5927
rect 10313 5894 10327 5908
rect 10393 5893 10407 5907
rect 10333 5852 10347 5866
rect 10373 5852 10387 5866
rect 10273 5693 10287 5707
rect 10313 5594 10327 5608
rect 10353 5593 10367 5607
rect 10373 5572 10387 5586
rect 10453 6113 10467 6127
rect 10453 6073 10467 6087
rect 10453 5993 10467 6007
rect 10473 5852 10487 5866
rect 10473 5793 10487 5807
rect 10573 6493 10587 6507
rect 10553 6473 10567 6487
rect 10533 6413 10547 6427
rect 10693 6493 10707 6507
rect 10693 6453 10707 6467
rect 10593 6433 10607 6447
rect 10613 6414 10627 6428
rect 10513 6373 10527 6387
rect 10513 6313 10527 6327
rect 10693 6393 10707 6407
rect 10733 6513 10747 6527
rect 10913 6853 10927 6867
rect 10853 6634 10867 6648
rect 10833 6553 10847 6567
rect 10933 6633 10947 6647
rect 10933 6592 10947 6606
rect 10913 6533 10927 6547
rect 10973 7513 10987 7527
rect 11053 7493 11067 7507
rect 11013 7473 11027 7487
rect 11053 7454 11067 7468
rect 11093 7454 11107 7468
rect 11013 7412 11027 7426
rect 11073 7412 11087 7426
rect 11033 6892 11047 6906
rect 10973 6853 10987 6867
rect 10993 6813 11007 6827
rect 10973 6633 10987 6647
rect 10953 6513 10967 6527
rect 10733 6453 10747 6467
rect 10733 6414 10747 6428
rect 10533 6293 10547 6307
rect 10613 6253 10627 6267
rect 10673 6352 10687 6366
rect 10713 6313 10727 6327
rect 10653 6193 10667 6207
rect 10633 6113 10647 6127
rect 10553 6072 10567 6086
rect 10553 6013 10567 6027
rect 10513 5913 10527 5927
rect 10593 5993 10607 6007
rect 10673 6033 10687 6047
rect 10653 5913 10667 5927
rect 10593 5894 10607 5908
rect 10653 5892 10667 5906
rect 10573 5852 10587 5866
rect 10513 5813 10527 5827
rect 10613 5813 10627 5827
rect 10673 5753 10687 5767
rect 10493 5713 10507 5727
rect 10613 5713 10627 5727
rect 10653 5713 10667 5727
rect 10473 5693 10487 5707
rect 10293 5552 10307 5566
rect 10273 5513 10287 5527
rect 10333 5513 10347 5527
rect 10333 5473 10347 5487
rect 10333 5393 10347 5407
rect 10833 6273 10847 6287
rect 10873 6273 10887 6287
rect 10813 6133 10827 6147
rect 10753 6073 10767 6087
rect 10733 5953 10747 5967
rect 10713 5653 10727 5667
rect 10473 5473 10487 5487
rect 10833 6072 10847 6086
rect 10773 6033 10787 6047
rect 10933 6193 10947 6207
rect 10913 6072 10927 6086
rect 10913 6033 10927 6047
rect 10833 5913 10847 5927
rect 10893 5913 10907 5927
rect 10773 5832 10787 5846
rect 10853 5852 10867 5866
rect 10813 5793 10827 5807
rect 10773 5733 10787 5747
rect 10753 5613 10767 5627
rect 10913 5853 10927 5867
rect 10813 5613 10827 5627
rect 10853 5613 10867 5627
rect 10713 5393 10727 5407
rect 10393 5373 10407 5387
rect 10433 5373 10447 5387
rect 10473 5373 10487 5387
rect 10853 5573 10867 5587
rect 10853 5413 10867 5427
rect 10813 5393 10827 5407
rect 10373 5354 10387 5368
rect 10413 5354 10427 5368
rect 10273 5333 10287 5347
rect 10313 5332 10327 5346
rect 10353 5333 10367 5347
rect 10353 5293 10367 5307
rect 10293 5253 10307 5267
rect 10613 5313 10627 5327
rect 10613 5253 10627 5267
rect 10473 5213 10487 5227
rect 10533 5213 10547 5227
rect 10413 5193 10427 5207
rect 10433 5133 10447 5147
rect 10253 5113 10267 5127
rect 10293 5113 10307 5127
rect 10253 5052 10267 5066
rect 10253 5033 10267 5047
rect 10433 5073 10447 5087
rect 10833 5354 10847 5368
rect 10753 5313 10767 5327
rect 10813 5313 10827 5327
rect 10853 5273 10867 5287
rect 10773 5233 10787 5247
rect 10753 5213 10767 5227
rect 10613 5193 10627 5207
rect 10593 5094 10607 5108
rect 10713 5094 10727 5108
rect 10553 5052 10567 5066
rect 10633 5053 10647 5067
rect 10533 5033 10547 5047
rect 10653 5033 10667 5047
rect 10293 4933 10307 4947
rect 10233 4893 10247 4907
rect 10113 4854 10127 4868
rect 10173 4854 10187 4868
rect 10213 4854 10227 4868
rect 10273 4854 10287 4868
rect 10073 4733 10087 4747
rect 10133 4673 10147 4687
rect 10193 4812 10207 4826
rect 10233 4812 10247 4826
rect 10233 4653 10247 4667
rect 10153 4633 10167 4647
rect 10213 4633 10227 4647
rect 10473 4913 10487 4927
rect 10433 4854 10447 4868
rect 10413 4812 10427 4826
rect 10453 4713 10467 4727
rect 10673 4713 10687 4727
rect 10533 4673 10547 4687
rect 10293 4633 10307 4647
rect 10233 4613 10247 4627
rect 10273 4613 10287 4627
rect 10113 4513 10127 4527
rect 9973 4193 9987 4207
rect 9993 4033 10007 4047
rect 9993 3973 10007 3987
rect 10073 4393 10087 4407
rect 10113 4373 10127 4387
rect 10033 4292 10047 4306
rect 10033 4253 10047 4267
rect 10093 4253 10107 4267
rect 10213 4554 10227 4568
rect 10193 4393 10207 4407
rect 10173 4273 10187 4287
rect 10133 4253 10147 4267
rect 10113 4233 10127 4247
rect 10173 4213 10187 4227
rect 10093 4173 10107 4187
rect 10593 4574 10607 4588
rect 10653 4574 10667 4588
rect 10753 5093 10767 5107
rect 10793 5093 10807 5107
rect 10313 4532 10327 4546
rect 10353 4534 10367 4548
rect 10493 4534 10507 4548
rect 10253 4493 10267 4507
rect 10273 4453 10287 4467
rect 10313 4393 10327 4407
rect 10313 4334 10327 4348
rect 10293 4253 10307 4267
rect 10333 4193 10347 4207
rect 10233 4173 10247 4187
rect 10713 4573 10727 4587
rect 10613 4532 10627 4546
rect 10653 4513 10667 4527
rect 10473 4413 10487 4427
rect 10593 4413 10607 4427
rect 10453 4333 10467 4347
rect 10453 4233 10467 4247
rect 10573 4373 10587 4387
rect 10533 4334 10547 4348
rect 10573 4334 10587 4348
rect 10913 5613 10927 5627
rect 10913 5573 10927 5587
rect 10893 5373 10907 5387
rect 10953 6114 10967 6128
rect 11113 7393 11127 7407
rect 11113 7293 11127 7307
rect 11153 7154 11167 7168
rect 11153 6893 11167 6907
rect 11073 6653 11087 6667
rect 11113 6653 11127 6667
rect 11053 6634 11067 6648
rect 11073 6592 11087 6606
rect 11093 6553 11107 6567
rect 11013 6533 11027 6547
rect 11033 6513 11047 6527
rect 11093 6253 11107 6267
rect 11033 6173 11047 6187
rect 11093 6173 11107 6187
rect 11033 6133 11047 6147
rect 10993 6114 11007 6128
rect 11013 6072 11027 6086
rect 10973 6033 10987 6047
rect 10953 6013 10967 6027
rect 10993 5973 11007 5987
rect 10973 5953 10987 5967
rect 10953 5894 10967 5908
rect 10953 5853 10967 5867
rect 11073 5973 11087 5987
rect 11113 5973 11127 5987
rect 11053 5933 11067 5947
rect 11033 5894 11047 5908
rect 11093 5933 11107 5947
rect 11113 5893 11127 5907
rect 11053 5852 11067 5866
rect 10993 5833 11007 5847
rect 11073 5733 11087 5747
rect 11073 5712 11087 5726
rect 11153 6633 11167 6647
rect 11133 5733 11147 5747
rect 11113 5713 11127 5727
rect 11153 5713 11167 5727
rect 11093 5693 11107 5707
rect 11093 5633 11107 5647
rect 11073 5593 11087 5607
rect 10933 5433 10947 5447
rect 10913 5354 10927 5368
rect 10913 5313 10927 5327
rect 10873 5033 10887 5047
rect 10893 4993 10907 5007
rect 11233 8233 11247 8247
rect 11193 8172 11207 8186
rect 11313 8173 11327 8187
rect 11193 8133 11207 8147
rect 11293 8133 11307 8147
rect 11253 8113 11267 8127
rect 11213 8033 11227 8047
rect 11293 8053 11307 8067
rect 11193 7893 11207 7907
rect 11273 7893 11287 7907
rect 11253 7853 11267 7867
rect 11193 7652 11207 7666
rect 11293 7653 11307 7667
rect 11193 7453 11207 7467
rect 11233 7154 11247 7168
rect 11193 6712 11207 6726
rect 11273 6892 11287 6906
rect 11313 7453 11327 7467
rect 11313 7353 11327 7367
rect 11293 6713 11307 6727
rect 11273 6634 11287 6648
rect 11313 6633 11327 6647
rect 11233 6593 11247 6607
rect 11213 6573 11227 6587
rect 11253 6573 11267 6587
rect 11233 6313 11247 6327
rect 11233 6213 11247 6227
rect 11333 6573 11347 6587
rect 11293 6553 11307 6567
rect 11253 6193 11267 6207
rect 11253 6072 11267 6086
rect 11193 6033 11207 6047
rect 11213 6013 11227 6027
rect 11293 6013 11307 6027
rect 11193 5813 11207 5827
rect 11193 5713 11207 5727
rect 11253 5894 11267 5908
rect 11273 5852 11287 5866
rect 11313 5833 11327 5847
rect 11213 5653 11227 5667
rect 11193 5633 11207 5647
rect 11273 5813 11287 5827
rect 11333 5733 11347 5747
rect 11313 5653 11327 5667
rect 11233 5614 11247 5628
rect 11273 5612 11287 5626
rect 11193 5572 11207 5586
rect 11253 5533 11267 5547
rect 11173 5373 11187 5387
rect 11073 5352 11087 5366
rect 10953 5213 10967 5227
rect 11253 5353 11267 5367
rect 11213 5313 11227 5327
rect 10993 5193 11007 5207
rect 11173 5172 11187 5186
rect 11153 5133 11167 5147
rect 11027 5093 11041 5107
rect 11033 5074 11047 5088
rect 10953 5033 10967 5047
rect 10933 4993 10947 5007
rect 10853 4933 10867 4947
rect 10873 4873 10887 4887
rect 10913 4873 10927 4887
rect 10873 4554 10887 4568
rect 10853 4453 10867 4467
rect 10673 4413 10687 4427
rect 10753 4413 10767 4427
rect 10513 4292 10527 4306
rect 10553 4253 10567 4267
rect 10473 4193 10487 4207
rect 10533 4193 10547 4207
rect 10613 4193 10627 4207
rect 10233 4113 10247 4127
rect 10373 4113 10387 4127
rect 10133 3993 10147 4007
rect 9933 3813 9947 3827
rect 9953 3794 9967 3808
rect 9873 3772 9887 3786
rect 9913 3772 9927 3786
rect 9973 3733 9987 3747
rect 9953 3573 9967 3587
rect 9813 3553 9827 3567
rect 9893 3553 9907 3567
rect 9793 3514 9807 3528
rect 9833 3514 9847 3528
rect 9793 3453 9807 3467
rect 9773 3373 9787 3387
rect 9773 3352 9787 3366
rect 9833 3433 9847 3447
rect 9813 3353 9827 3367
rect 9793 3293 9807 3307
rect 9853 3333 9867 3347
rect 9873 3313 9887 3327
rect 9913 3514 9927 3528
rect 9913 3453 9927 3467
rect 9953 3513 9967 3527
rect 9933 3433 9947 3447
rect 9913 3313 9927 3327
rect 9893 3293 9907 3307
rect 9793 3253 9807 3267
rect 9933 3293 9947 3307
rect 9793 3193 9807 3207
rect 9753 3012 9767 3026
rect 9593 2853 9607 2867
rect 9733 2853 9747 2867
rect 9633 2793 9647 2807
rect 9673 2793 9687 2807
rect 9613 2573 9627 2587
rect 9593 2473 9607 2487
rect 9753 2773 9767 2787
rect 9693 2732 9707 2746
rect 9673 2513 9687 2527
rect 9593 2413 9607 2427
rect 9573 2293 9587 2307
rect 9533 2253 9547 2267
rect 9513 2193 9527 2207
rect 9493 1933 9507 1947
rect 9473 1912 9487 1926
rect 9473 1653 9487 1667
rect 9453 1553 9467 1567
rect 9553 2113 9567 2127
rect 9573 2053 9587 2067
rect 9533 1993 9547 2007
rect 9593 2033 9607 2047
rect 9653 2433 9667 2447
rect 9633 2213 9647 2227
rect 9653 2193 9667 2207
rect 9693 2333 9707 2347
rect 9753 2693 9767 2707
rect 9733 2653 9747 2667
rect 9733 2333 9747 2347
rect 9733 2293 9747 2307
rect 9773 2433 9787 2447
rect 9753 2273 9767 2287
rect 9753 2212 9767 2226
rect 9673 2133 9687 2147
rect 9653 2093 9667 2107
rect 9613 1993 9627 2007
rect 9613 1954 9627 1968
rect 9673 1954 9687 1968
rect 9553 1873 9567 1887
rect 9533 1833 9547 1847
rect 9533 1734 9547 1748
rect 9493 1453 9507 1467
rect 9413 1434 9427 1448
rect 9453 1434 9467 1448
rect 9473 1392 9487 1406
rect 9413 1353 9427 1367
rect 9473 1353 9487 1367
rect 9413 1313 9427 1327
rect 9373 1233 9387 1247
rect 9393 1172 9407 1186
rect 9393 1113 9407 1127
rect 9433 1073 9447 1087
rect 9473 1033 9487 1047
rect 9673 1913 9687 1927
rect 9613 1873 9627 1887
rect 9593 1813 9607 1827
rect 9653 1833 9667 1847
rect 9553 1692 9567 1706
rect 9553 1653 9567 1667
rect 9493 993 9507 1007
rect 9533 993 9547 1007
rect 9433 914 9447 928
rect 9513 933 9527 947
rect 9493 893 9507 907
rect 9353 873 9367 887
rect 9413 872 9427 886
rect 9473 853 9487 867
rect 9453 793 9467 807
rect 9533 793 9547 807
rect 9513 713 9527 727
rect 9333 473 9347 487
rect 9293 413 9307 427
rect 9333 413 9347 427
rect 9213 352 9227 366
rect 9253 352 9267 366
rect 9173 293 9187 307
rect 9133 273 9147 287
rect 9453 493 9467 507
rect 9453 394 9467 408
rect 9393 373 9407 387
rect 9433 333 9447 347
rect 9393 293 9407 307
rect 9393 253 9407 267
rect 9453 253 9467 267
rect 9333 233 9347 247
rect 8913 193 8927 207
rect 8893 173 8907 187
rect 8733 132 8747 146
rect 8773 132 8787 146
rect 8873 132 8887 146
rect 8633 73 8647 87
rect 8873 73 8887 87
rect 8613 53 8627 67
rect 8733 53 8747 67
rect 8973 174 8987 188
rect 9133 173 9147 187
rect 9193 174 9207 188
rect 8913 132 8927 146
rect 8953 132 8967 146
rect 8993 93 9007 107
rect 9433 193 9447 207
rect 9393 174 9407 188
rect 9313 132 9327 146
rect 9413 132 9427 146
rect 9453 132 9467 146
rect 9173 113 9187 127
rect 9213 113 9227 127
rect 9333 93 9347 107
rect 8973 73 8987 87
rect 9133 73 9147 87
rect 9313 73 9327 87
rect 8893 33 8907 47
rect 9593 1692 9607 1706
rect 9593 1533 9607 1547
rect 9593 1433 9607 1447
rect 9573 1393 9587 1407
rect 9633 1593 9647 1607
rect 9633 1553 9647 1567
rect 9633 1473 9647 1487
rect 9613 1313 9627 1327
rect 9713 2013 9727 2027
rect 9913 3233 9927 3247
rect 9873 3113 9887 3127
rect 9853 3053 9867 3067
rect 9833 2992 9847 3006
rect 9813 2973 9827 2987
rect 9833 2913 9847 2927
rect 9833 2833 9847 2847
rect 9813 2693 9827 2707
rect 9813 2553 9827 2567
rect 10013 3913 10027 3927
rect 10053 3973 10067 3987
rect 10573 4133 10587 4147
rect 10533 4093 10547 4107
rect 10533 4054 10547 4068
rect 10373 4014 10387 4028
rect 10473 4014 10487 4028
rect 10233 3993 10247 4007
rect 10173 3913 10187 3927
rect 10293 3913 10307 3927
rect 10053 3873 10067 3887
rect 10013 3794 10027 3808
rect 10493 3993 10507 4007
rect 10473 3833 10487 3847
rect 10053 3733 10067 3747
rect 10173 3653 10187 3667
rect 10153 3613 10167 3627
rect 10133 3553 10147 3567
rect 9993 3513 10007 3527
rect 10073 3533 10087 3547
rect 10053 3472 10067 3486
rect 10033 3413 10047 3427
rect 10013 3373 10027 3387
rect 9993 3293 10007 3307
rect 9973 3153 9987 3167
rect 9913 2933 9927 2947
rect 9873 2813 9887 2827
rect 9953 2813 9967 2827
rect 9853 2493 9867 2507
rect 9853 2432 9867 2446
rect 9833 2273 9847 2287
rect 9853 2113 9867 2127
rect 9833 2073 9847 2087
rect 9833 1993 9847 2007
rect 9713 1773 9727 1787
rect 9713 1734 9727 1748
rect 9733 1473 9747 1487
rect 9693 1433 9707 1447
rect 9733 1434 9747 1448
rect 9793 1953 9807 1967
rect 9813 1912 9827 1926
rect 9773 1813 9787 1827
rect 9913 2774 9927 2788
rect 9893 2613 9907 2627
rect 9893 2493 9907 2507
rect 10173 3493 10187 3507
rect 10353 3673 10367 3687
rect 10293 3653 10307 3667
rect 10213 3514 10227 3528
rect 10313 3593 10327 3607
rect 10413 3593 10427 3607
rect 10273 3514 10287 3528
rect 10353 3553 10367 3567
rect 10353 3513 10367 3527
rect 10372 3492 10386 3506
rect 10393 3493 10407 3507
rect 10212 3473 10226 3487
rect 10233 3473 10247 3487
rect 10253 3453 10267 3467
rect 10193 3433 10207 3447
rect 10153 3413 10167 3427
rect 10133 3373 10147 3387
rect 10053 3333 10067 3347
rect 10093 3333 10107 3347
rect 10093 3294 10107 3308
rect 10193 3393 10207 3407
rect 10233 3393 10247 3407
rect 10013 3253 10027 3267
rect 9993 3113 10007 3127
rect 9973 2593 9987 2607
rect 9973 2533 9987 2547
rect 9953 2373 9967 2387
rect 9973 2293 9987 2307
rect 9933 2254 9947 2268
rect 9973 2254 9987 2268
rect 9913 2213 9927 2227
rect 9893 2173 9907 2187
rect 9893 1953 9907 1967
rect 9893 1913 9907 1927
rect 9873 1853 9887 1867
rect 9933 2193 9947 2207
rect 10033 2893 10047 2907
rect 10113 3252 10127 3266
rect 10073 3193 10087 3207
rect 10073 3033 10087 3047
rect 10093 2994 10107 3008
rect 10093 2933 10107 2947
rect 10053 2774 10067 2788
rect 10113 2893 10127 2907
rect 10213 3353 10227 3367
rect 10333 3453 10347 3467
rect 10373 3453 10387 3467
rect 10293 3433 10307 3447
rect 10333 3413 10347 3427
rect 10473 3793 10487 3807
rect 10453 3533 10467 3547
rect 10513 3933 10527 3947
rect 10773 4233 10787 4247
rect 10933 4753 10947 4767
rect 10953 4553 10967 4567
rect 11053 5032 11067 5046
rect 11093 4993 11107 5007
rect 11013 4953 11027 4967
rect 11053 4933 11067 4947
rect 11153 5032 11167 5046
rect 11073 4812 11087 4826
rect 11153 4812 11167 4826
rect 11013 4793 11027 4807
rect 11253 5313 11267 5327
rect 11233 5233 11247 5247
rect 11293 5573 11307 5587
rect 11273 5233 11287 5247
rect 11293 5173 11307 5187
rect 11093 4753 11107 4767
rect 10993 4633 11007 4647
rect 11053 4533 11067 4547
rect 11013 4333 11027 4347
rect 10973 4292 10987 4306
rect 11053 4273 11067 4287
rect 10973 4193 10987 4207
rect 10693 4093 10707 4107
rect 10633 4053 10647 4067
rect 10673 4053 10687 4067
rect 10593 3993 10607 4007
rect 10513 3893 10527 3907
rect 10573 3893 10587 3907
rect 10653 3813 10667 3827
rect 10513 3772 10527 3786
rect 10553 3772 10567 3786
rect 10493 3733 10507 3747
rect 10593 3733 10607 3747
rect 10633 3733 10647 3747
rect 10833 4014 10847 4028
rect 10813 3873 10827 3887
rect 10853 3833 10867 3847
rect 10793 3753 10807 3767
rect 10873 3772 10887 3786
rect 10773 3673 10787 3687
rect 10413 3433 10427 3447
rect 10613 3494 10627 3508
rect 10453 3473 10467 3487
rect 10393 3413 10407 3427
rect 10433 3413 10447 3427
rect 10373 3393 10387 3407
rect 10473 3433 10487 3447
rect 10453 3393 10467 3407
rect 10433 3373 10447 3387
rect 10253 3333 10267 3347
rect 10253 3233 10267 3247
rect 10193 2933 10207 2947
rect 10193 2873 10207 2887
rect 10033 2733 10047 2747
rect 10093 2733 10107 2747
rect 10133 2732 10147 2746
rect 10073 2573 10087 2587
rect 10033 2432 10047 2446
rect 10033 2373 10047 2387
rect 9953 2153 9967 2167
rect 9933 2133 9947 2147
rect 9933 2053 9947 2067
rect 9953 1973 9967 1987
rect 9933 1893 9947 1907
rect 10013 2133 10027 2147
rect 10113 2693 10127 2707
rect 10093 2093 10107 2107
rect 10013 2073 10027 2087
rect 10073 1954 10087 1968
rect 10173 2593 10187 2607
rect 10133 2453 10147 2467
rect 10233 2974 10247 2988
rect 10233 2873 10247 2887
rect 10213 2813 10227 2827
rect 10513 3393 10527 3407
rect 10593 3393 10607 3407
rect 10493 3173 10507 3187
rect 10393 3153 10407 3167
rect 10413 3033 10427 3047
rect 10392 2974 10406 2988
rect 10413 2973 10427 2987
rect 10373 2813 10387 2827
rect 10333 2774 10347 2788
rect 10313 2713 10327 2727
rect 10253 2573 10267 2587
rect 10253 2513 10267 2527
rect 10353 2513 10367 2527
rect 10293 2474 10307 2488
rect 10193 2413 10207 2427
rect 10173 2254 10187 2268
rect 10193 2212 10207 2226
rect 10313 2432 10327 2446
rect 10273 2413 10287 2427
rect 10353 2413 10367 2427
rect 10273 2333 10287 2347
rect 10253 2293 10267 2307
rect 10153 2193 10167 2207
rect 10193 2173 10207 2187
rect 9953 1833 9967 1847
rect 9913 1793 9927 1807
rect 9893 1734 9907 1748
rect 9973 1734 9987 1748
rect 9773 1693 9787 1707
rect 9813 1613 9827 1627
rect 9673 1392 9687 1406
rect 9713 1392 9727 1406
rect 9753 1353 9767 1367
rect 9653 1333 9667 1347
rect 9693 1333 9707 1347
rect 9633 1293 9647 1307
rect 9573 1233 9587 1247
rect 9553 493 9567 507
rect 9613 1214 9627 1228
rect 9653 1214 9667 1228
rect 9633 1133 9647 1147
rect 9593 1073 9607 1087
rect 9653 993 9667 1007
rect 9593 933 9607 947
rect 9593 872 9607 886
rect 9633 872 9647 886
rect 9713 1293 9727 1307
rect 9733 1053 9747 1067
rect 9733 872 9747 886
rect 9713 833 9727 847
rect 9693 753 9707 767
rect 9673 652 9687 666
rect 9713 613 9727 627
rect 9573 433 9587 447
rect 9653 413 9667 427
rect 9673 333 9687 347
rect 9573 293 9587 307
rect 9553 193 9567 207
rect 9653 273 9667 287
rect 9593 233 9607 247
rect 9573 173 9587 187
rect 9593 153 9607 167
rect 9753 413 9767 427
rect 9733 333 9747 347
rect 9733 253 9747 267
rect 9633 132 9647 146
rect 9553 73 9567 87
rect 9533 53 9547 67
rect 9713 133 9727 147
rect 9673 73 9687 87
rect 9693 53 9707 67
rect 9793 1434 9807 1448
rect 9853 1653 9867 1667
rect 9853 1573 9867 1587
rect 9833 1553 9847 1567
rect 9813 1392 9827 1406
rect 9973 1533 9987 1547
rect 9873 1493 9887 1507
rect 9933 1473 9947 1487
rect 9853 1392 9867 1406
rect 9913 1392 9927 1406
rect 9953 1392 9967 1406
rect 9833 1253 9847 1267
rect 9913 1253 9927 1267
rect 9833 1214 9847 1228
rect 9873 1214 9887 1228
rect 9853 1172 9867 1186
rect 9853 993 9867 1007
rect 9973 1253 9987 1267
rect 9953 1214 9967 1228
rect 9933 1093 9947 1107
rect 9933 1033 9947 1047
rect 9913 953 9927 967
rect 9853 933 9867 947
rect 9793 913 9807 927
rect 9973 1013 9987 1027
rect 9953 913 9967 927
rect 9833 872 9847 886
rect 9873 872 9887 886
rect 9913 872 9927 886
rect 9913 833 9927 847
rect 9853 753 9867 767
rect 9852 653 9866 667
rect 9873 652 9887 666
rect 9973 652 9987 666
rect 9793 573 9807 587
rect 9793 493 9807 507
rect 9913 493 9927 507
rect 9813 393 9827 407
rect 9873 394 9887 408
rect 9813 352 9827 366
rect 9853 352 9867 366
rect 9933 353 9947 367
rect 9893 333 9907 347
rect 9853 313 9867 327
rect 9793 132 9807 146
rect 9873 132 9887 146
rect 10113 1913 10127 1927
rect 10153 1913 10167 1927
rect 10053 1893 10067 1907
rect 10093 1873 10107 1887
rect 10133 1873 10147 1887
rect 10033 1853 10047 1867
rect 10013 1833 10027 1847
rect 10013 1393 10027 1407
rect 10093 1793 10107 1807
rect 10113 1734 10127 1748
rect 10053 1693 10067 1707
rect 10093 1553 10107 1567
rect 10073 1533 10087 1547
rect 10073 1353 10087 1367
rect 10153 1493 10167 1507
rect 10133 1473 10147 1487
rect 10253 2212 10267 2226
rect 10553 3213 10567 3227
rect 10513 3053 10527 3067
rect 10833 3733 10847 3747
rect 10813 3673 10827 3687
rect 10793 3533 10807 3547
rect 10753 3494 10767 3508
rect 10733 3473 10747 3487
rect 10613 3313 10627 3327
rect 10613 3213 10627 3227
rect 10593 3013 10607 3027
rect 10513 2972 10527 2986
rect 10593 2973 10607 2987
rect 10633 2974 10647 2988
rect 10613 2933 10627 2947
rect 10593 2873 10607 2887
rect 10633 2893 10647 2907
rect 10633 2872 10647 2886
rect 10613 2853 10627 2867
rect 10453 2793 10467 2807
rect 10493 2793 10507 2807
rect 10433 2474 10447 2488
rect 10433 2433 10447 2447
rect 10573 2774 10587 2788
rect 10553 2732 10567 2746
rect 10513 2713 10527 2727
rect 10573 2593 10587 2607
rect 10473 2573 10487 2587
rect 10533 2493 10547 2507
rect 10493 2474 10507 2488
rect 10473 2433 10487 2447
rect 10453 2373 10467 2387
rect 10333 2273 10347 2287
rect 10373 2273 10387 2287
rect 10433 2273 10447 2287
rect 10313 2173 10327 2187
rect 10313 2133 10327 2147
rect 10393 2254 10407 2268
rect 10353 2213 10367 2227
rect 10333 1993 10347 2007
rect 10293 1873 10307 1887
rect 10273 1793 10287 1807
rect 10213 1653 10227 1667
rect 10213 1613 10227 1627
rect 10153 1453 10167 1467
rect 10193 1453 10207 1467
rect 10253 1753 10267 1767
rect 10553 2433 10567 2447
rect 10513 2413 10527 2427
rect 10513 2373 10527 2387
rect 10493 2273 10507 2287
rect 10473 2193 10487 2207
rect 10413 2173 10427 2187
rect 10393 2133 10407 2147
rect 10373 2113 10387 2127
rect 10373 1953 10387 1967
rect 10353 1893 10367 1907
rect 10333 1753 10347 1767
rect 10293 1692 10307 1706
rect 10273 1653 10287 1667
rect 10293 1493 10307 1507
rect 10233 1453 10247 1467
rect 10093 1253 10107 1267
rect 10093 1214 10107 1228
rect 10073 1172 10087 1186
rect 10073 1133 10087 1147
rect 10133 1173 10147 1187
rect 10113 1093 10127 1107
rect 10133 1053 10147 1067
rect 10053 993 10067 1007
rect 10133 993 10147 1007
rect 10093 914 10107 928
rect 10133 914 10147 928
rect 10073 872 10087 886
rect 10053 733 10067 747
rect 10013 473 10027 487
rect 10013 433 10027 447
rect 10193 1293 10207 1307
rect 10173 1214 10187 1228
rect 10173 1113 10187 1127
rect 10173 993 10187 1007
rect 10093 652 10107 666
rect 10153 652 10167 666
rect 10153 573 10167 587
rect 10073 433 10087 447
rect 10093 394 10107 408
rect 10073 353 10087 367
rect 10113 352 10127 366
rect 10053 333 10067 347
rect 10213 1172 10227 1186
rect 10213 973 10227 987
rect 10193 813 10207 827
rect 10193 694 10207 708
rect 10213 652 10227 666
rect 10193 613 10207 627
rect 10213 473 10227 487
rect 10133 154 10147 168
rect 10173 154 10187 168
rect 10213 152 10227 166
rect 10013 132 10027 146
rect 10053 132 10067 146
rect 10253 1392 10267 1406
rect 10253 1333 10267 1347
rect 10293 1233 10307 1247
rect 10273 1214 10287 1228
rect 10333 1473 10347 1487
rect 10413 1954 10427 1968
rect 10393 1913 10407 1927
rect 10413 1853 10427 1867
rect 10413 1813 10427 1827
rect 10393 1753 10407 1767
rect 10373 1513 10387 1527
rect 10413 1693 10427 1707
rect 10393 1493 10407 1507
rect 10393 1434 10407 1448
rect 10373 1392 10387 1406
rect 10393 1373 10407 1387
rect 10293 1172 10307 1186
rect 10333 1153 10347 1167
rect 10353 1133 10367 1147
rect 10253 1113 10267 1127
rect 10293 1073 10307 1087
rect 10333 914 10347 928
rect 10273 872 10287 886
rect 10273 793 10287 807
rect 10333 773 10347 787
rect 10313 694 10327 708
rect 10413 1233 10427 1247
rect 10413 1172 10427 1186
rect 10413 1073 10427 1087
rect 10413 833 10427 847
rect 10533 2233 10547 2247
rect 10553 2212 10567 2226
rect 10533 2153 10547 2167
rect 10493 2133 10507 2147
rect 10473 1954 10487 1968
rect 10513 1954 10527 1968
rect 10453 1913 10467 1927
rect 10533 1893 10547 1907
rect 10493 1873 10507 1887
rect 10453 1773 10467 1787
rect 10493 1734 10507 1748
rect 10553 1813 10567 1827
rect 10473 1653 10487 1667
rect 10473 1533 10487 1547
rect 10453 1433 10467 1447
rect 10513 1613 10527 1627
rect 10533 1493 10547 1507
rect 10513 1373 10527 1387
rect 10493 1293 10507 1307
rect 10593 2493 10607 2507
rect 10793 3493 10807 3507
rect 10793 3393 10807 3407
rect 10793 3333 10807 3347
rect 10833 3553 10847 3567
rect 10913 3733 10927 3747
rect 10853 3493 10867 3507
rect 10833 3453 10847 3467
rect 10813 3313 10827 3327
rect 10833 3294 10847 3308
rect 10893 3553 10907 3567
rect 10913 3533 10927 3547
rect 10893 3473 10907 3487
rect 10873 3233 10887 3247
rect 10913 3393 10927 3407
rect 10893 3213 10907 3227
rect 10773 3193 10787 3207
rect 10853 3193 10867 3207
rect 10913 3193 10927 3207
rect 10753 3173 10767 3187
rect 10733 3113 10747 3127
rect 10913 3153 10927 3167
rect 10773 3013 10787 3027
rect 10773 2974 10787 2988
rect 10873 2873 10887 2887
rect 10713 2853 10727 2867
rect 10773 2833 10787 2847
rect 10733 2774 10747 2788
rect 10813 2793 10827 2807
rect 10713 2653 10727 2667
rect 10673 2593 10687 2607
rect 10793 2693 10807 2707
rect 10813 2474 10827 2488
rect 10613 2433 10627 2447
rect 10593 2333 10607 2347
rect 10633 2254 10647 2268
rect 10753 2393 10767 2407
rect 10753 2313 10767 2327
rect 10613 2212 10627 2226
rect 10613 2173 10627 2187
rect 10593 1954 10607 1968
rect 10693 2213 10707 2227
rect 10853 2333 10867 2347
rect 10773 2253 10787 2267
rect 10893 2773 10907 2787
rect 10873 2213 10887 2227
rect 10752 2173 10766 2187
rect 10773 2173 10787 2187
rect 10653 2153 10667 2167
rect 10653 2093 10667 2107
rect 10633 1993 10647 2007
rect 10613 1873 10627 1887
rect 10613 1773 10627 1787
rect 10593 1733 10607 1747
rect 10673 2013 10687 2027
rect 10733 1954 10747 1968
rect 10773 1954 10787 1968
rect 10673 1912 10687 1926
rect 10713 1912 10727 1926
rect 10793 1913 10807 1927
rect 10653 1873 10667 1887
rect 10753 1873 10767 1887
rect 10733 1833 10747 1847
rect 10673 1733 10687 1747
rect 10833 2153 10847 2167
rect 10813 1833 10827 1847
rect 10773 1734 10787 1748
rect 10673 1692 10687 1706
rect 10713 1692 10727 1706
rect 10753 1653 10767 1667
rect 10733 1633 10747 1647
rect 10713 1593 10727 1607
rect 10633 1533 10647 1547
rect 10593 1473 10607 1487
rect 10573 1453 10587 1467
rect 10673 1453 10687 1467
rect 10633 1434 10647 1448
rect 10573 1333 10587 1347
rect 10533 1233 10547 1247
rect 10513 1214 10527 1228
rect 10533 1113 10547 1127
rect 10493 1093 10507 1107
rect 10473 1073 10487 1087
rect 10453 953 10467 967
rect 10633 1233 10647 1247
rect 10613 1053 10627 1067
rect 10593 973 10607 987
rect 10553 953 10567 967
rect 10493 933 10507 947
rect 10473 914 10487 928
rect 10513 914 10527 928
rect 10493 872 10507 886
rect 10533 833 10547 847
rect 10453 793 10467 807
rect 10393 733 10407 747
rect 10433 713 10447 727
rect 10293 652 10307 666
rect 10333 633 10347 647
rect 10333 553 10347 567
rect 10273 453 10287 467
rect 10353 493 10367 507
rect 10433 673 10447 687
rect 10393 453 10407 467
rect 10333 413 10347 427
rect 10393 394 10407 408
rect 10493 694 10507 708
rect 10533 694 10547 708
rect 10553 633 10567 647
rect 10653 1133 10667 1147
rect 10633 572 10647 586
rect 10493 433 10507 447
rect 10473 394 10487 408
rect 10593 433 10607 447
rect 10293 313 10307 327
rect 10373 352 10387 366
rect 10413 352 10427 366
rect 10453 352 10467 366
rect 10333 293 10347 307
rect 10473 253 10487 267
rect 10373 152 10387 166
rect 10613 352 10627 366
rect 10093 113 10107 127
rect 10233 113 10247 127
rect 10853 1893 10867 1907
rect 10873 1673 10887 1687
rect 10853 1653 10867 1667
rect 10833 1613 10847 1627
rect 10813 1593 10827 1607
rect 10773 1434 10787 1448
rect 10873 1434 10887 1448
rect 10993 4093 11007 4107
rect 11033 4053 11047 4067
rect 10953 4012 10967 4026
rect 11073 4253 11087 4267
rect 11053 4033 11067 4047
rect 11033 3993 11047 4007
rect 10953 3973 10967 3987
rect 11013 3953 11027 3967
rect 10993 3913 11007 3927
rect 10953 3853 10967 3867
rect 10953 3772 10967 3786
rect 11113 4553 11127 4567
rect 11113 4133 11127 4147
rect 11253 5074 11267 5088
rect 11273 5032 11287 5046
rect 11233 4953 11247 4967
rect 11153 4593 11167 4607
rect 11193 4593 11207 4607
rect 11193 4554 11207 4568
rect 11273 4673 11287 4687
rect 11213 4493 11227 4507
rect 11233 4334 11247 4348
rect 11213 4292 11227 4306
rect 11153 4073 11167 4087
rect 11173 4034 11187 4048
rect 11253 4073 11267 4087
rect 11233 4013 11247 4027
rect 11093 3953 11107 3967
rect 11073 3913 11087 3927
rect 11093 3853 11107 3867
rect 10953 3733 10967 3747
rect 11193 3992 11207 4006
rect 11153 3753 11167 3767
rect 11073 3693 11087 3707
rect 11113 3693 11127 3707
rect 11233 3673 11247 3687
rect 11072 3494 11086 3508
rect 11173 3533 11187 3547
rect 11253 3533 11267 3547
rect 11093 3493 11107 3507
rect 11033 3393 11047 3407
rect 11072 3393 11086 3407
rect 11113 3393 11127 3407
rect 10973 3294 10987 3308
rect 10993 3252 11007 3266
rect 10933 3013 10947 3027
rect 10973 3013 10987 3027
rect 10953 2972 10967 2986
rect 10933 2913 10947 2927
rect 10913 2733 10927 2747
rect 10953 2813 10967 2827
rect 10993 2893 11007 2907
rect 11073 3293 11087 3307
rect 11093 3253 11107 3267
rect 11073 3193 11087 3207
rect 11053 3133 11067 3147
rect 11033 2873 11047 2887
rect 11013 2813 11027 2827
rect 10973 2773 10987 2787
rect 11093 3053 11107 3067
rect 11073 2972 11087 2986
rect 11053 2774 11067 2788
rect 10933 2713 10947 2727
rect 11033 2713 11047 2727
rect 10993 2673 11007 2687
rect 11053 2673 11067 2687
rect 10953 2653 10967 2667
rect 10993 2633 11007 2647
rect 11013 2613 11027 2627
rect 10953 2413 10967 2427
rect 10933 2373 10947 2387
rect 10913 2313 10927 2327
rect 11013 2413 11027 2427
rect 11033 2373 11047 2387
rect 10973 2333 10987 2347
rect 10973 2254 10987 2268
rect 11073 2413 11087 2427
rect 11133 3333 11147 3347
rect 11192 3492 11206 3506
rect 11213 3493 11227 3507
rect 11193 3453 11207 3467
rect 11193 3393 11207 3407
rect 11333 4193 11347 4207
rect 11292 3493 11306 3507
rect 11313 3493 11327 3507
rect 11273 3447 11287 3461
rect 11213 3333 11227 3347
rect 11173 3313 11187 3327
rect 11213 3294 11227 3308
rect 11253 3253 11267 3267
rect 11193 3233 11207 3247
rect 11153 3213 11167 3227
rect 11173 3013 11187 3027
rect 11153 2613 11167 2627
rect 11253 3013 11267 3027
rect 11193 2913 11207 2927
rect 11193 2873 11207 2887
rect 11173 2533 11187 2547
rect 11293 3413 11307 3427
rect 11273 2873 11287 2887
rect 11273 2813 11287 2827
rect 11213 2793 11227 2807
rect 11253 2793 11267 2807
rect 11233 2732 11247 2746
rect 11253 2533 11267 2547
rect 11193 2513 11207 2527
rect 11173 2474 11187 2488
rect 11213 2474 11227 2488
rect 11093 2313 11107 2327
rect 11093 2254 11107 2268
rect 10993 2212 11007 2226
rect 11033 2212 11047 2226
rect 10953 2153 10967 2167
rect 11093 2193 11107 2207
rect 11073 2173 11087 2187
rect 11073 1993 11087 2007
rect 10993 1954 11007 1968
rect 10953 1912 10967 1926
rect 11013 1912 11027 1926
rect 10933 1853 10947 1867
rect 10913 1793 10927 1807
rect 10913 1734 10927 1748
rect 10953 1773 10967 1787
rect 10993 1734 11007 1748
rect 11053 1734 11067 1748
rect 10753 1393 10767 1407
rect 10713 1353 10727 1367
rect 10733 1293 10747 1307
rect 10713 1172 10727 1186
rect 10733 1133 10747 1147
rect 10713 773 10727 787
rect 10693 613 10707 627
rect 10753 753 10767 767
rect 10813 1392 10827 1406
rect 10813 1353 10827 1367
rect 10873 1373 10887 1387
rect 10853 1333 10867 1347
rect 10813 1173 10827 1187
rect 10793 1133 10807 1147
rect 10853 973 10867 987
rect 10833 913 10847 927
rect 10853 833 10867 847
rect 10833 793 10847 807
rect 10893 1333 10907 1347
rect 10893 1153 10907 1167
rect 11013 1673 11027 1687
rect 10933 1373 10947 1387
rect 10953 1333 10967 1347
rect 10973 1214 10987 1228
rect 10933 1172 10947 1186
rect 10993 1172 11007 1186
rect 10913 993 10927 1007
rect 10933 914 10947 928
rect 10913 833 10927 847
rect 10953 793 10967 807
rect 10953 694 10967 708
rect 11033 1633 11047 1647
rect 11073 1692 11087 1706
rect 11113 1893 11127 1907
rect 11173 2413 11187 2427
rect 11233 2433 11247 2447
rect 11153 2353 11167 2367
rect 11153 2313 11167 2327
rect 11193 2393 11207 2407
rect 11173 2254 11187 2268
rect 11153 2193 11167 2207
rect 11213 2353 11227 2367
rect 11213 2273 11227 2287
rect 11193 2153 11207 2167
rect 11273 2513 11287 2527
rect 11293 2393 11307 2407
rect 11273 2293 11287 2307
rect 11253 2273 11267 2287
rect 11293 2254 11307 2268
rect 11233 2213 11247 2227
rect 11293 2153 11307 2167
rect 11253 1993 11267 2007
rect 11173 1954 11187 1968
rect 11213 1954 11227 1968
rect 11153 1913 11167 1927
rect 11133 1873 11147 1887
rect 11113 1853 11127 1867
rect 11113 1773 11127 1787
rect 11093 1573 11107 1587
rect 11073 1553 11087 1567
rect 11073 1293 11087 1307
rect 11032 1214 11046 1228
rect 11053 1213 11067 1227
rect 11053 1173 11067 1187
rect 11053 1152 11067 1166
rect 11013 853 11027 867
rect 11053 733 11067 747
rect 11053 694 11067 708
rect 10873 673 10887 687
rect 10773 652 10787 666
rect 10973 652 10987 666
rect 10713 533 10727 547
rect 10693 373 10707 387
rect 10773 453 10787 467
rect 10753 394 10767 408
rect 10813 413 10827 427
rect 11013 493 11027 507
rect 11133 1693 11147 1707
rect 11193 1873 11207 1887
rect 11233 1853 11247 1867
rect 11213 1793 11227 1807
rect 11253 1734 11267 1748
rect 11193 1692 11207 1706
rect 11153 1653 11167 1667
rect 11233 1653 11247 1667
rect 11213 1613 11227 1627
rect 11293 1613 11307 1627
rect 11253 1573 11267 1587
rect 11213 1373 11227 1387
rect 11273 1373 11287 1387
rect 11193 1293 11207 1307
rect 11233 1214 11247 1228
rect 11173 1172 11187 1186
rect 11213 1113 11227 1127
rect 11273 1113 11287 1127
rect 11073 652 11087 666
rect 11053 453 11067 467
rect 11153 914 11167 928
rect 11113 733 11127 747
rect 11093 413 11107 427
rect 10853 394 10867 408
rect 10973 394 10987 408
rect 11053 394 11067 408
rect 11153 853 11167 867
rect 11133 613 11147 627
rect 11133 413 11147 427
rect 10752 353 10766 367
rect 10773 353 10787 367
rect 10833 352 10847 366
rect 10873 352 10887 366
rect 10973 352 10987 366
rect 11073 313 11087 327
rect 11053 233 11067 247
rect 11293 973 11307 987
rect 11253 694 11267 708
rect 11193 652 11207 666
rect 11233 613 11247 627
rect 11153 313 11167 327
rect 10733 132 10747 146
rect 10533 112 10547 126
rect 10673 112 10687 126
rect 10873 132 10887 146
rect 9933 93 9947 107
rect 10753 93 10767 107
rect 11133 132 11147 146
rect 11333 2353 11347 2367
rect 11333 2293 11347 2307
rect 11333 132 11347 146
rect 11313 93 11327 107
rect 9733 33 9747 47
rect 9773 33 9787 47
rect 11093 33 11107 47
rect 7033 13 7047 27
rect 7513 13 7527 27
rect 7673 13 7687 27
rect 8593 13 8607 27
rect 8973 13 8987 27
rect 9633 13 9647 27
<< metal3 >>
rect 6507 11176 10253 11184
rect 10267 11176 10453 11184
rect 2907 11156 3793 11164
rect 1807 11136 1913 11144
rect 2287 11136 2573 11144
rect 3227 11136 3373 11144
rect 3487 11136 3853 11144
rect 4787 11136 4833 11144
rect 5087 11136 5613 11144
rect 5747 11136 6033 11144
rect 6607 11136 6853 11144
rect 6867 11136 6933 11144
rect 6947 11136 7073 11144
rect 7387 11136 7813 11144
rect 8967 11136 9073 11144
rect 1367 11116 1833 11124
rect 1847 11116 1873 11124
rect 1887 11116 2204 11124
rect 2196 11108 2204 11116
rect 8007 11116 8273 11124
rect 8287 11116 9093 11124
rect 9187 11116 9633 11124
rect -63 11097 13 11105
rect 27 11097 193 11105
rect 867 11096 1073 11104
rect 1227 11096 1313 11104
rect 1527 11096 1553 11104
rect 2067 11097 2093 11105
rect 2207 11097 2233 11105
rect 2367 11096 2493 11104
rect 3267 11097 3313 11105
rect 3407 11097 3433 11105
rect 3547 11096 3693 11104
rect 4887 11097 5013 11105
rect 5056 11097 5213 11105
rect 347 11076 493 11084
rect 807 11077 913 11085
rect 2587 11075 2713 11083
rect 167 11056 413 11064
rect 1127 11056 1293 11064
rect 1347 11056 1393 11064
rect 1607 11056 1773 11064
rect 2307 11055 2353 11063
rect 2956 11064 2964 11074
rect 2527 11056 2964 11064
rect 3007 11056 3393 11064
rect 3407 11056 3513 11064
rect 3527 11055 3673 11063
rect 3756 11064 3764 11074
rect 3867 11075 3993 11083
rect 3727 11056 3764 11064
rect 5056 11064 5064 11097
rect 5293 11097 5393 11105
rect 5007 11056 5064 11064
rect 413 11044 426 11052
rect 413 11036 1053 11044
rect 1067 11036 1533 11044
rect 2207 11036 2484 11044
rect 2476 11027 2484 11036
rect 3507 11036 3533 11044
rect 2267 11016 2313 11024
rect 2487 11016 2993 11024
rect 3487 11016 3713 11024
rect 5293 11024 5301 11097
rect 5867 11097 5933 11105
rect 6427 11097 6453 11105
rect 6567 11096 6713 11104
rect 7147 11096 7193 11104
rect 7307 11097 7333 11105
rect 7487 11097 7593 11105
rect 7867 11096 7904 11104
rect 7896 11084 7904 11096
rect 7927 11096 8073 11104
rect 8327 11096 8513 11104
rect 8747 11096 8873 11104
rect 9007 11097 9033 11105
rect 9407 11096 9472 11104
rect 9507 11096 9593 11104
rect 9787 11097 9833 11105
rect 9887 11096 10053 11104
rect 10307 11096 10344 11104
rect 10336 11087 10344 11096
rect 10387 11096 10513 11104
rect 10527 11096 10633 11104
rect 10687 11097 10713 11105
rect 10767 11096 10804 11104
rect 7896 11076 7933 11084
rect 10336 11076 10353 11087
rect 10340 11073 10353 11076
rect 10796 11084 10804 11096
rect 10827 11096 10973 11104
rect 11147 11097 11173 11105
rect 10796 11076 10864 11084
rect 7167 11056 7353 11064
rect 7367 11056 7573 11064
rect 7887 11055 7913 11063
rect 7967 11055 8053 11063
rect 8887 11055 8933 11063
rect 9387 11055 9493 11063
rect 9667 11055 9693 11063
rect 10087 11056 10273 11064
rect 10327 11055 10373 11063
rect 10856 11064 10864 11076
rect 10856 11056 10953 11064
rect 11007 11056 11193 11064
rect 6327 11036 6473 11044
rect 7087 11036 7393 11044
rect 7407 11036 7513 11044
rect 8347 11036 8713 11044
rect 8727 11036 9113 11044
rect 9367 11036 9853 11044
rect 10467 11036 10533 11044
rect 10647 11036 10773 11044
rect 4987 11016 5301 11024
rect 7127 11016 7153 11024
rect 7167 11016 7293 11024
rect 8547 11016 8973 11024
rect 627 10996 793 11004
rect 807 10996 1093 11004
rect 1747 10996 1813 11004
rect 7447 10996 8093 11004
rect 9087 10996 9893 11004
rect 9907 10996 10344 11004
rect 2567 10976 2573 10984
rect 2587 10976 3013 10984
rect 3027 10976 3453 10984
rect 3467 10976 4153 10984
rect 7047 10976 7833 10984
rect 10336 10984 10344 10996
rect 10336 10976 10493 10984
rect 10507 10976 10653 10984
rect 10707 10976 10733 10984
rect 1747 10956 5913 10964
rect 7927 10956 8753 10964
rect 8767 10956 9033 10964
rect 9047 10956 9153 10964
rect 2767 10936 3133 10944
rect 6707 10936 7113 10944
rect 7187 10936 7473 10944
rect 9627 10936 10293 10944
rect 10307 10936 10813 10944
rect 4107 10916 4173 10924
rect 4187 10916 4473 10924
rect 4487 10916 4553 10924
rect 8047 10916 8293 10924
rect 10367 10916 10673 10924
rect 27 10896 1733 10904
rect 7947 10896 9653 10904
rect 9667 10896 9793 10904
rect 1227 10876 4113 10884
rect 4127 10876 5493 10884
rect 6107 10876 6453 10884
rect 7487 10876 8393 10884
rect 9207 10876 9273 10884
rect 9287 10876 9393 10884
rect 10547 10876 10733 10884
rect 1547 10856 1933 10864
rect 1947 10856 1973 10864
rect 2687 10856 2753 10864
rect 3727 10856 5353 10864
rect 5567 10856 6493 10864
rect 8467 10856 8513 10864
rect 10107 10856 10513 10864
rect 10527 10856 10753 10864
rect 6067 10836 6553 10844
rect 7307 10836 7333 10844
rect 7507 10836 7553 10844
rect 8227 10836 8253 10844
rect 8607 10836 8733 10844
rect 9247 10836 9433 10844
rect 9447 10836 9933 10844
rect 10567 10836 11133 10844
rect 447 10816 453 10824
rect 467 10816 493 10824
rect 507 10816 1033 10824
rect 1047 10817 1153 10825
rect 1807 10816 2713 10824
rect 2727 10816 2833 10824
rect 2967 10816 3373 10824
rect 4087 10816 4153 10824
rect 4167 10816 4533 10824
rect 4547 10817 4813 10825
rect 6827 10816 6913 10824
rect 6927 10816 7373 10824
rect 7527 10816 7573 10824
rect 8367 10816 8493 10824
rect 9767 10816 9853 10824
rect 2027 10797 2173 10805
rect 2507 10796 2553 10804
rect 2927 10797 3073 10805
rect 3447 10796 3613 10804
rect 5887 10796 6053 10804
rect 6167 10797 6273 10805
rect 6367 10797 6633 10805
rect 6747 10797 6773 10805
rect 6947 10796 6993 10804
rect 7007 10797 7113 10805
rect 7127 10796 7253 10804
rect 7607 10797 7773 10805
rect 7827 10797 7893 10805
rect 7947 10796 7993 10804
rect 8167 10797 8213 10805
rect 8267 10796 8333 10804
rect 8527 10797 8693 10805
rect 8707 10796 8933 10804
rect 9047 10796 9193 10804
rect 287 10777 413 10785
rect 567 10777 653 10785
rect 1067 10776 1193 10784
rect 107 10756 833 10764
rect 1316 10764 1324 10774
rect 1527 10775 1553 10783
rect 3927 10777 4013 10785
rect 7796 10776 7913 10784
rect 1316 10756 1673 10764
rect 1127 10736 1213 10744
rect 2316 10724 2324 10773
rect 2567 10755 2653 10763
rect 2707 10756 2893 10764
rect 3176 10764 3184 10774
rect 2947 10756 3184 10764
rect 3387 10756 3633 10764
rect 3647 10756 3713 10764
rect 4047 10756 4173 10764
rect 3747 10736 3773 10744
rect 3787 10736 4193 10744
rect 4376 10744 4384 10774
rect 5607 10755 5713 10763
rect 6087 10756 6153 10764
rect 6207 10755 6333 10763
rect 6507 10755 7013 10763
rect 7027 10756 7173 10764
rect 7367 10755 7433 10763
rect 7796 10766 7804 10776
rect 7447 10755 7513 10763
rect 7567 10756 7753 10764
rect 8027 10756 8153 10764
rect 8247 10756 8313 10764
rect 8407 10755 8433 10763
rect 8667 10755 8913 10763
rect 8967 10756 9073 10764
rect 9416 10766 9424 10813
rect 9587 10797 9613 10805
rect 9856 10796 9893 10804
rect 9636 10776 9693 10784
rect 9636 10766 9644 10776
rect 9856 10784 9864 10796
rect 9907 10796 10053 10804
rect 10347 10797 10373 10805
rect 10827 10797 10893 10805
rect 10556 10784 10564 10794
rect 10967 10796 11013 10804
rect 11087 10796 11213 10804
rect 9707 10776 9864 10784
rect 9916 10776 10564 10784
rect 9127 10755 9173 10763
rect 9227 10755 9273 10763
rect 9916 10764 9924 10776
rect 9887 10756 9924 10764
rect 10116 10766 10124 10776
rect 9947 10756 10073 10764
rect 10387 10756 10533 10764
rect 10667 10755 10753 10763
rect 11007 10755 11073 10763
rect 4376 10736 4673 10744
rect 6427 10736 6573 10744
rect 6647 10736 6933 10744
rect 7067 10736 7313 10744
rect 10907 10736 11033 10744
rect 2267 10716 2324 10724
rect 3736 10724 3744 10733
rect 3367 10716 3744 10724
rect 5807 10716 6113 10724
rect 7316 10724 7324 10733
rect 7316 10716 7793 10724
rect 8147 10716 8333 10724
rect 8847 10716 9013 10724
rect 9807 10716 9833 10724
rect 1047 10696 1213 10704
rect 2187 10696 2713 10704
rect 2847 10696 2973 10704
rect 4207 10696 4233 10704
rect 5707 10696 6293 10704
rect 6307 10696 6993 10704
rect 7007 10696 8673 10704
rect 10847 10696 11233 10704
rect 47 10676 173 10684
rect 387 10676 473 10684
rect 567 10676 633 10684
rect 3087 10676 3153 10684
rect 5867 10676 6193 10684
rect 6387 10676 6453 10684
rect 6467 10676 6533 10684
rect 6547 10676 6733 10684
rect 7147 10676 8653 10684
rect 847 10656 913 10664
rect 927 10656 1273 10664
rect 1287 10656 1493 10664
rect 1507 10656 1713 10664
rect 7467 10656 7493 10664
rect 8107 10656 8173 10664
rect 8727 10656 10073 10664
rect 287 10636 413 10644
rect 2007 10636 2073 10644
rect 6487 10636 7273 10644
rect 7287 10636 7653 10644
rect 7667 10636 8033 10644
rect 8047 10636 8193 10644
rect 8487 10636 9573 10644
rect 587 10616 853 10624
rect 1707 10616 1993 10624
rect 2047 10616 2413 10624
rect 3307 10616 3373 10624
rect 4147 10616 4233 10624
rect 4247 10616 4293 10624
rect 4627 10616 4933 10624
rect 5367 10616 5393 10624
rect 5407 10616 5593 10624
rect 5827 10616 6173 10624
rect 6747 10616 7193 10624
rect 7247 10616 8073 10624
rect 9247 10616 9373 10624
rect 9427 10616 9473 10624
rect 10067 10616 10413 10624
rect 10427 10616 10533 10624
rect 10687 10616 10833 10624
rect 10947 10616 11033 10624
rect 347 10596 393 10604
rect 8107 10596 8313 10604
rect 8327 10596 8553 10604
rect 147 10577 373 10585
rect 1967 10576 2153 10584
rect 2176 10576 2233 10584
rect 207 10536 393 10544
rect 447 10535 473 10543
rect 587 10535 613 10543
rect 727 10536 833 10544
rect 896 10544 904 10573
rect 1547 10555 1693 10563
rect 2176 10564 2184 10576
rect 2247 10576 2373 10584
rect 2567 10577 2673 10585
rect 2767 10576 2893 10584
rect 2907 10577 2953 10585
rect 3127 10577 3213 10585
rect 3227 10576 3313 10584
rect 1976 10556 2184 10564
rect 1976 10546 1984 10556
rect 887 10536 904 10544
rect 2027 10535 2073 10543
rect 2507 10536 2533 10544
rect 2607 10536 2653 10544
rect 2707 10536 2913 10544
rect 2927 10536 3093 10544
rect 3356 10527 3364 10574
rect 3447 10576 3573 10584
rect 3807 10576 3933 10584
rect 4067 10577 4093 10585
rect 4467 10576 4573 10584
rect 4636 10576 4713 10584
rect 4636 10564 4644 10576
rect 4807 10577 5133 10585
rect 5287 10577 5333 10585
rect 5687 10577 5853 10585
rect 5967 10576 6053 10584
rect 6187 10576 6473 10584
rect 6527 10576 6633 10584
rect 6907 10577 6953 10585
rect 6967 10576 7053 10584
rect 7607 10576 7933 10584
rect 8187 10576 8544 10584
rect 4607 10556 4644 10564
rect 8536 10564 8544 10576
rect 8567 10576 8753 10584
rect 8767 10577 8793 10585
rect 8907 10576 9053 10584
rect 9107 10577 9273 10585
rect 9287 10576 9453 10584
rect 9507 10576 9693 10584
rect 9867 10577 9893 10585
rect 10047 10577 10133 10585
rect 10367 10576 10493 10584
rect 10807 10576 10913 10584
rect 6807 10556 7264 10564
rect 8536 10556 8733 10564
rect 3387 10535 3473 10543
rect 3487 10535 3533 10543
rect 3687 10536 3813 10544
rect 3947 10535 3993 10543
rect 4047 10535 4193 10543
rect 4307 10535 4433 10543
rect 4587 10535 4653 10543
rect 4867 10536 4893 10544
rect 5327 10536 5373 10544
rect 5587 10536 5793 10544
rect 6007 10535 6033 10543
rect 6327 10536 6493 10544
rect 6507 10536 6713 10544
rect 7027 10536 7113 10544
rect 7256 10546 7264 10556
rect 10576 10564 10584 10574
rect 10967 10577 10993 10585
rect 11167 10576 11233 10584
rect 10576 10556 10633 10564
rect 7367 10536 7393 10544
rect 7467 10536 7493 10544
rect 7507 10536 7633 10544
rect 7887 10536 7953 10544
rect 8047 10535 8113 10543
rect 8347 10535 8433 10543
rect 8787 10536 8853 10544
rect 8867 10535 8893 10543
rect 9387 10535 9473 10543
rect 9727 10536 9753 10544
rect 9927 10536 10033 10544
rect 10107 10536 10333 10544
rect 10507 10535 10593 10543
rect 10707 10535 10813 10543
rect 10927 10535 11013 10543
rect 11067 10535 11133 10543
rect 11227 10535 11333 10543
rect 4967 10516 5113 10524
rect 5987 10516 6073 10524
rect 6987 10516 7213 10524
rect 8587 10516 8673 10524
rect 10387 10516 10413 10524
rect 1807 10496 2213 10504
rect 3327 10496 3593 10504
rect 6587 10496 7333 10504
rect 7347 10496 7613 10504
rect 7627 10496 7693 10504
rect 7707 10496 8213 10504
rect 8747 10496 10053 10504
rect 10167 10496 10553 10504
rect 10747 10496 11253 10504
rect 927 10476 1213 10484
rect 1227 10476 1373 10484
rect 4827 10476 5173 10484
rect 5227 10476 5673 10484
rect 5907 10476 6113 10484
rect 6127 10476 6253 10484
rect 6576 10484 6584 10493
rect 6267 10476 6584 10484
rect 6647 10476 6724 10484
rect 2447 10456 2553 10464
rect 2567 10456 2593 10464
rect 4667 10456 4833 10464
rect 6716 10464 6724 10476
rect 6747 10476 6893 10484
rect 8667 10476 8813 10484
rect 9267 10476 9853 10484
rect 6716 10456 6933 10464
rect 7667 10456 8732 10464
rect 8767 10456 9053 10464
rect 887 10436 1213 10444
rect 1347 10436 1773 10444
rect 6547 10436 6633 10444
rect 7547 10436 9333 10444
rect 10607 10436 10953 10444
rect 1247 10416 2753 10424
rect 4687 10416 5533 10424
rect 5547 10416 5653 10424
rect 5807 10416 6073 10424
rect 6207 10416 7133 10424
rect 7447 10416 9084 10424
rect 547 10396 633 10404
rect 2367 10396 3773 10404
rect 3787 10396 4093 10404
rect 5207 10396 5773 10404
rect 6827 10396 7253 10404
rect 7316 10396 7673 10404
rect 2427 10376 2653 10384
rect 2667 10376 3393 10384
rect 3467 10376 3673 10384
rect 4096 10384 4104 10393
rect 4096 10376 4313 10384
rect 4467 10376 4853 10384
rect 5836 10376 6113 10384
rect 5836 10367 5844 10376
rect 6867 10376 6973 10384
rect 6987 10376 7053 10384
rect 7316 10384 7324 10396
rect 9076 10404 9084 10416
rect 9507 10416 10293 10424
rect 9076 10396 10653 10404
rect 10667 10396 10813 10404
rect 10827 10396 10853 10404
rect 7127 10376 7324 10384
rect 7887 10376 8153 10384
rect 8167 10376 8373 10384
rect 8387 10376 8613 10384
rect 1087 10356 1533 10364
rect 2967 10356 3052 10364
rect 3087 10356 3133 10364
rect 5307 10356 5393 10364
rect 5527 10356 5833 10364
rect 6487 10356 7533 10364
rect 9847 10356 10513 10364
rect 10527 10356 10593 10364
rect 10607 10356 10773 10364
rect 847 10336 1873 10344
rect 3987 10336 4113 10344
rect 4167 10336 4513 10344
rect 4527 10336 4793 10344
rect 4867 10336 5973 10344
rect 6947 10336 7013 10344
rect 7567 10336 7853 10344
rect 407 10316 633 10324
rect 647 10316 1073 10324
rect 2507 10316 2813 10324
rect 3127 10316 3233 10324
rect 4047 10316 4253 10324
rect 5507 10316 5653 10324
rect 5807 10316 5933 10324
rect 6547 10316 6853 10324
rect 6867 10316 7113 10324
rect 7127 10316 7313 10324
rect 7387 10316 7513 10324
rect 7527 10316 7893 10324
rect 8127 10316 8273 10324
rect 8287 10316 8453 10324
rect 8467 10316 8593 10324
rect 8607 10316 9033 10324
rect 9047 10316 9313 10324
rect 9327 10316 9373 10324
rect 9427 10316 9473 10324
rect 9787 10316 10553 10324
rect 1787 10296 1813 10304
rect 3627 10296 4453 10304
rect 5127 10296 5393 10304
rect 7427 10296 7473 10304
rect 8707 10296 9073 10304
rect 9447 10296 9593 10304
rect 187 10276 253 10284
rect 507 10277 593 10285
rect 727 10277 793 10285
rect 1207 10277 1293 10285
rect 896 10256 944 10264
rect 267 10235 373 10243
rect 627 10236 713 10244
rect 896 10246 904 10256
rect 936 10244 944 10256
rect 936 10236 1093 10244
rect 1116 10227 1124 10274
rect 1147 10236 1193 10244
rect 1636 10244 1644 10274
rect 1687 10276 2033 10284
rect 2287 10277 2333 10285
rect 2347 10276 2453 10284
rect 2647 10277 2673 10285
rect 2716 10264 2724 10274
rect 2787 10276 2913 10284
rect 4107 10277 4273 10285
rect 4367 10277 4473 10285
rect 5447 10277 5473 10285
rect 5587 10277 5613 10285
rect 2716 10256 2793 10264
rect 3156 10264 3164 10274
rect 5727 10276 6013 10284
rect 6467 10277 6533 10285
rect 6707 10277 6773 10285
rect 6907 10277 7013 10285
rect 2807 10256 3164 10264
rect 3587 10256 3713 10264
rect 3756 10256 3812 10264
rect 1636 10236 1833 10244
rect 1927 10235 2053 10243
rect 2747 10235 2773 10243
rect 2827 10236 2933 10244
rect 3087 10236 3133 10244
rect 3247 10236 3333 10244
rect 3347 10235 3413 10243
rect 3547 10236 3633 10244
rect 1527 10216 1573 10224
rect 2327 10216 2693 10224
rect 3187 10216 3293 10224
rect 3756 10224 3764 10256
rect 3847 10257 3993 10265
rect 4307 10236 4353 10244
rect 4707 10236 4833 10244
rect 3727 10216 3764 10224
rect 4376 10216 4493 10224
rect 687 10196 853 10204
rect 1367 10196 1473 10204
rect 1547 10196 1613 10204
rect 3227 10196 3433 10204
rect 4376 10204 4384 10216
rect 5016 10224 5024 10254
rect 5147 10256 5313 10264
rect 5167 10236 5233 10244
rect 5387 10236 5493 10244
rect 5607 10236 5733 10244
rect 5987 10235 6053 10243
rect 6107 10236 6193 10244
rect 6407 10235 6553 10243
rect 6607 10236 6693 10244
rect 7296 10244 7304 10274
rect 7327 10276 7653 10284
rect 7676 10276 7713 10284
rect 7676 10264 7684 10276
rect 7767 10277 7813 10285
rect 7867 10277 7913 10285
rect 7927 10277 7933 10285
rect 8507 10277 8653 10285
rect 8767 10276 8873 10284
rect 8887 10277 8993 10285
rect 9807 10276 9893 10284
rect 10067 10277 10113 10285
rect 7656 10260 7684 10264
rect 7653 10256 7684 10260
rect 7653 10247 7667 10256
rect 7296 10236 7493 10244
rect 7827 10236 7953 10244
rect 8607 10235 8633 10243
rect 8727 10235 8973 10243
rect 9067 10235 9153 10243
rect 9416 10244 9424 10273
rect 9396 10236 9424 10244
rect 5016 10216 5233 10224
rect 6747 10216 6793 10224
rect 7047 10216 7233 10224
rect 7287 10216 7433 10224
rect 8207 10216 8393 10224
rect 4007 10196 4384 10204
rect 4427 10196 4613 10204
rect 4847 10196 4873 10204
rect 5347 10196 6133 10204
rect 6767 10196 6833 10204
rect 6847 10196 6933 10204
rect 7527 10196 7733 10204
rect 8187 10196 8433 10204
rect 8447 10196 8493 10204
rect 8547 10196 8673 10204
rect 8747 10196 9193 10204
rect 9396 10206 9404 10236
rect 9867 10235 10093 10243
rect 10356 10227 10364 10274
rect 10927 10276 11013 10284
rect 10587 10236 10993 10244
rect 9687 10196 9833 10204
rect 10647 10196 11033 10204
rect 1227 10176 1353 10184
rect 1567 10176 1773 10184
rect 2387 10176 2753 10184
rect 2947 10176 2973 10184
rect 2987 10176 3133 10184
rect 6647 10176 6813 10184
rect 7627 10176 8133 10184
rect 9447 10176 9913 10184
rect 9927 10176 10013 10184
rect 10027 10176 10053 10184
rect 10067 10176 10333 10184
rect 2067 10156 3533 10164
rect 3727 10156 3873 10164
rect 4187 10156 4773 10164
rect 5107 10156 5213 10164
rect 5447 10156 7693 10164
rect 7707 10156 8173 10164
rect 8327 10156 9233 10164
rect 1427 10136 1793 10144
rect 2787 10136 3153 10144
rect 4267 10136 4373 10144
rect 4387 10136 4533 10144
rect 4547 10136 4753 10144
rect 6727 10136 7393 10144
rect 7687 10136 8113 10144
rect 8307 10136 9253 10144
rect 9307 10136 9733 10144
rect 9787 10136 9893 10144
rect 10047 10136 10133 10144
rect 11007 10136 11253 10144
rect 327 10116 453 10124
rect 827 10116 1093 10124
rect 1107 10116 1233 10124
rect 2267 10116 2373 10124
rect 2487 10116 2533 10124
rect 2767 10116 3993 10124
rect 4007 10116 4673 10124
rect 4727 10116 4873 10124
rect 5327 10116 5473 10124
rect 6167 10116 6213 10124
rect 6227 10116 6493 10124
rect 6647 10116 8313 10124
rect 8487 10116 8713 10124
rect 227 10096 493 10104
rect 507 10096 1033 10104
rect 1047 10096 1113 10104
rect 1207 10096 1853 10104
rect 2067 10096 2233 10104
rect 2407 10096 2493 10104
rect 2507 10096 2633 10104
rect 2927 10096 3284 10104
rect 2007 10076 2853 10084
rect 3276 10084 3284 10096
rect 4787 10096 5573 10104
rect 8947 10096 8973 10104
rect 9247 10096 9573 10104
rect 9587 10096 10133 10104
rect 10147 10096 10193 10104
rect 10207 10096 10373 10104
rect 10527 10096 10593 10104
rect 11047 10096 11293 10104
rect 3276 10076 3633 10084
rect 4027 10076 4693 10084
rect 6287 10076 6393 10084
rect 9087 10076 9173 10084
rect 9627 10076 9793 10084
rect 10767 10076 10813 10084
rect 187 10057 253 10065
rect 427 10057 513 10065
rect 587 10057 653 10065
rect 867 10057 1173 10065
rect 1727 10057 1753 10065
rect 1927 10056 1993 10064
rect 2216 10056 2413 10064
rect 1867 10036 2053 10044
rect 447 10015 493 10023
rect 1487 10016 1573 10024
rect 1587 10016 1713 10024
rect 2216 10026 2224 10056
rect 2467 10057 2553 10065
rect 2607 10056 2713 10064
rect 2907 10056 2973 10064
rect 3027 10056 3213 10064
rect 3307 10056 3473 10064
rect 3707 10057 3933 10065
rect 4147 10057 4273 10065
rect 4967 10056 5033 10064
rect 5087 10057 5153 10065
rect 5207 10056 5253 10064
rect 5367 10057 5393 10065
rect 5587 10057 5653 10065
rect 6207 10057 6473 10065
rect 6567 10057 6593 10065
rect 4727 10037 4753 10045
rect 4807 10036 5093 10044
rect 5736 10044 5744 10054
rect 6676 10044 6684 10054
rect 6747 10056 6913 10064
rect 6927 10057 6973 10065
rect 7187 10057 7553 10065
rect 7813 10064 7827 10073
rect 7787 10060 7827 10064
rect 7787 10056 7824 10060
rect 7867 10056 7993 10064
rect 8247 10056 8313 10064
rect 8367 10057 8433 10065
rect 8627 10056 8673 10064
rect 8847 10057 8893 10065
rect 9107 10056 9133 10064
rect 9367 10056 9513 10064
rect 9687 10056 9853 10064
rect 9967 10056 10093 10064
rect 10327 10056 10433 10064
rect 10507 10057 10553 10065
rect 10787 10064 10800 10067
rect 10787 10053 10804 10064
rect 10987 10056 11073 10064
rect 5547 10036 5744 10044
rect 6636 10036 6864 10044
rect 2387 10015 2433 10023
rect 3527 10016 3653 10024
rect 3727 10016 3733 10024
rect 3747 10016 4013 10024
rect 4027 10016 4053 10024
rect 4267 10016 4313 10024
rect 4867 10015 4973 10023
rect 4987 10016 5073 10024
rect 5247 10016 5353 10024
rect 5967 10016 5993 10024
rect 6067 10015 6133 10023
rect 6636 10024 6644 10036
rect 6856 10026 6864 10036
rect 10616 10036 10653 10044
rect 6427 10016 6644 10024
rect 6987 10016 7293 10024
rect 7547 10015 7613 10023
rect 7667 10015 7753 10023
rect 7807 10015 7853 10023
rect 8227 10015 8293 10023
rect 8387 10015 8453 10023
rect 8707 10015 8753 10023
rect 8867 10015 9153 10023
rect 9167 10016 9293 10024
rect 10616 10026 10624 10036
rect 10796 10026 10804 10053
rect 9807 10015 9833 10023
rect 10027 10015 10113 10023
rect 10447 10015 10533 10023
rect 10847 10015 10913 10023
rect 10967 10015 11093 10023
rect 527 9996 633 10004
rect 1227 9996 1773 10004
rect 1827 9996 1973 10004
rect 4367 9995 4813 10003
rect 4827 9995 4853 10003
rect 5427 9996 5513 10004
rect 5527 9996 5713 10004
rect 6207 9996 6313 10004
rect 6367 9996 6393 10004
rect 6667 9996 7053 10004
rect 7067 9996 7193 10004
rect 7207 9996 7493 10004
rect 9327 9996 9373 10004
rect 3067 9976 3233 9984
rect 3247 9976 3573 9984
rect 3647 9976 4133 9984
rect 4847 9976 4893 9984
rect 5047 9976 5213 9984
rect 5787 9976 5953 9984
rect 6187 9976 6553 9984
rect 7947 9976 8253 9984
rect 8267 9976 8353 9984
rect 9527 9976 9873 9984
rect 10087 9976 10293 9984
rect 10587 9976 11053 9984
rect 11067 9976 11193 9984
rect 2347 9956 3213 9964
rect 3267 9956 3373 9964
rect 3387 9956 3413 9964
rect 4167 9956 4393 9964
rect 4476 9956 4793 9964
rect 1887 9936 2273 9944
rect 2287 9936 3173 9944
rect 3216 9944 3224 9953
rect 3216 9936 3313 9944
rect 3547 9936 4233 9944
rect 4476 9944 4484 9956
rect 5447 9956 5553 9964
rect 5567 9956 5673 9964
rect 6827 9956 6853 9964
rect 6867 9956 7413 9964
rect 8447 9956 8493 9964
rect 8507 9956 8653 9964
rect 10827 9956 10893 9964
rect 11067 9956 11133 9964
rect 4247 9936 4484 9944
rect 4527 9936 5253 9944
rect 6627 9936 6873 9944
rect 8007 9936 8373 9944
rect 9087 9936 9413 9944
rect 9427 9936 9773 9944
rect 10087 9936 10713 9944
rect 2387 9916 4493 9924
rect 4507 9916 5233 9924
rect 7627 9916 8013 9924
rect 10107 9916 10493 9924
rect 10507 9916 10653 9924
rect 2887 9896 3453 9904
rect 3767 9896 4033 9904
rect 5187 9896 5273 9904
rect 5287 9896 5393 9904
rect 567 9876 833 9884
rect 2467 9876 2553 9884
rect 2567 9876 2693 9884
rect 2967 9876 3053 9884
rect 3567 9876 4113 9884
rect 4127 9876 4633 9884
rect 4747 9876 5013 9884
rect 6147 9876 6533 9884
rect 6547 9876 7273 9884
rect 7327 9876 7633 9884
rect 8027 9876 9113 9884
rect 207 9856 293 9864
rect 1727 9856 3113 9864
rect 3187 9856 4033 9864
rect 4047 9856 4333 9864
rect 4347 9856 4613 9864
rect 4696 9856 5093 9864
rect 4696 9847 4704 9856
rect 5107 9856 5313 9864
rect 5367 9856 5753 9864
rect 6627 9856 6793 9864
rect 7927 9856 7973 9864
rect 147 9836 413 9844
rect 427 9836 513 9844
rect 3167 9836 4693 9844
rect 4787 9836 5553 9844
rect 7976 9844 7984 9853
rect 7976 9836 8833 9844
rect 9536 9836 10333 9844
rect 9536 9827 9544 9836
rect 787 9816 1113 9824
rect 2547 9816 2633 9824
rect 3127 9816 5664 9824
rect 247 9796 573 9804
rect 2047 9796 2193 9804
rect 2747 9796 2893 9804
rect 3787 9796 3893 9804
rect 4007 9796 4253 9804
rect 4607 9796 5313 9804
rect 5367 9796 5433 9804
rect 5656 9804 5664 9816
rect 7247 9816 7593 9824
rect 7767 9816 9533 9824
rect 9947 9816 10213 9824
rect 10627 9816 10913 9824
rect 11167 9816 11213 9824
rect 5656 9796 5733 9804
rect 5927 9796 6473 9804
rect 6587 9796 6693 9804
rect 8467 9796 8893 9804
rect 9587 9796 9953 9804
rect 607 9777 753 9785
rect 767 9776 913 9784
rect 2407 9776 2493 9784
rect 2587 9776 2933 9784
rect 3667 9776 3733 9784
rect 3947 9776 4433 9784
rect 6367 9776 6733 9784
rect 7447 9776 7473 9784
rect 7847 9776 8713 9784
rect 8727 9776 8913 9784
rect 10487 9776 10753 9784
rect 147 9757 193 9765
rect 216 9756 253 9764
rect 216 9744 224 9756
rect 727 9756 893 9764
rect 1227 9756 1373 9764
rect 1427 9757 1453 9765
rect 1627 9757 1753 9765
rect 1847 9756 1933 9764
rect 2047 9756 2233 9764
rect 3127 9757 3173 9765
rect 3447 9757 3473 9765
rect 3627 9756 3813 9764
rect 3827 9757 3853 9765
rect 176 9736 224 9744
rect 176 9726 184 9736
rect 2447 9736 2613 9744
rect 3116 9744 3124 9754
rect 2987 9736 3124 9744
rect 227 9716 353 9724
rect 487 9716 633 9724
rect 1107 9716 1273 9724
rect 1327 9715 1353 9723
rect 1467 9716 1593 9724
rect 1787 9715 1813 9723
rect 1947 9715 2013 9723
rect 2107 9716 2253 9724
rect 3347 9716 3373 9724
rect 3507 9716 3633 9724
rect 3747 9716 3833 9724
rect 3896 9724 3904 9754
rect 3987 9756 4073 9764
rect 4487 9757 4553 9765
rect 4296 9727 4304 9754
rect 4827 9757 4913 9765
rect 5067 9757 5113 9765
rect 5267 9756 5433 9764
rect 5487 9756 5673 9764
rect 5693 9764 5707 9773
rect 5687 9760 5707 9764
rect 5687 9756 5704 9760
rect 5887 9756 6093 9764
rect 6227 9756 6313 9764
rect 6427 9757 6493 9765
rect 3847 9716 3904 9724
rect 4107 9716 4173 9724
rect 4287 9716 4304 9727
rect 4287 9713 4300 9716
rect 4327 9716 4473 9724
rect 4736 9724 4744 9753
rect 5836 9727 5844 9753
rect 6316 9744 6324 9754
rect 6507 9757 6613 9765
rect 6827 9757 6913 9765
rect 6967 9757 7013 9765
rect 7287 9757 7333 9765
rect 7427 9757 7513 9765
rect 7527 9756 7673 9764
rect 7807 9757 8053 9765
rect 8167 9757 8193 9765
rect 8247 9757 8513 9765
rect 8687 9756 8792 9764
rect 8827 9757 8853 9765
rect 9047 9757 9313 9765
rect 9367 9757 9653 9765
rect 9707 9757 9753 9765
rect 9807 9756 9993 9764
rect 10447 9756 10513 9764
rect 6316 9736 6444 9744
rect 4736 9716 4793 9724
rect 5007 9716 5133 9724
rect 5187 9715 5233 9723
rect 5507 9715 5713 9723
rect 6167 9716 6273 9724
rect 6347 9716 6413 9724
rect 6436 9724 6444 9736
rect 9796 9744 9804 9754
rect 6887 9736 7024 9744
rect 6436 9716 6753 9724
rect 6767 9716 6793 9724
rect 6887 9715 6993 9723
rect 7016 9724 7024 9736
rect 9536 9736 9804 9744
rect 10016 9736 10093 9744
rect 7016 9716 7033 9724
rect 7987 9716 8253 9724
rect 8267 9715 8293 9723
rect 8447 9715 8493 9723
rect 8887 9716 9033 9724
rect 9536 9724 9544 9736
rect 9347 9716 9544 9724
rect 9567 9716 9693 9724
rect 10016 9726 10024 9736
rect 9947 9716 9973 9724
rect 10256 9724 10264 9754
rect 10887 9757 10973 9765
rect 11076 9736 11273 9744
rect 11076 9726 11084 9736
rect 10256 9716 10453 9724
rect 10687 9715 10753 9723
rect 10907 9715 10993 9723
rect 327 9696 433 9704
rect 667 9696 693 9704
rect 2427 9696 2473 9704
rect 2927 9696 3213 9704
rect 3927 9696 3973 9704
rect 4267 9696 4353 9704
rect 4667 9696 4773 9704
rect 5867 9696 6053 9704
rect 6627 9696 6713 9704
rect 7307 9696 7413 9704
rect 7547 9696 7593 9704
rect 8667 9696 8713 9704
rect 8807 9696 8913 9704
rect 8927 9696 9013 9704
rect 9067 9696 9093 9704
rect 9107 9696 9153 9704
rect 1247 9676 1393 9684
rect 2067 9676 2373 9684
rect 3216 9684 3224 9693
rect 3216 9676 3713 9684
rect 4407 9676 4533 9684
rect 4707 9676 4753 9684
rect 5467 9676 5593 9684
rect 5847 9676 5872 9684
rect 5907 9676 6373 9684
rect 6927 9676 6993 9684
rect 7507 9676 7733 9684
rect 8947 9676 8973 9684
rect 9787 9676 10233 9684
rect 1307 9656 1633 9664
rect 2927 9656 3133 9664
rect 4587 9656 5033 9664
rect 5667 9656 6173 9664
rect 7147 9656 7573 9664
rect 7587 9656 8153 9664
rect 8167 9656 8473 9664
rect 8487 9656 8973 9664
rect 967 9636 1513 9644
rect 1527 9636 2293 9644
rect 2447 9636 2513 9644
rect 2527 9636 3413 9644
rect 3436 9636 3873 9644
rect 587 9616 873 9624
rect 1367 9616 2273 9624
rect 3436 9624 3444 9636
rect 3967 9636 4133 9644
rect 4207 9636 4313 9644
rect 4427 9636 4533 9644
rect 4907 9636 5053 9644
rect 5656 9644 5664 9653
rect 5327 9636 5664 9644
rect 6127 9636 6593 9644
rect 6807 9636 7153 9644
rect 7267 9636 8113 9644
rect 8507 9636 8913 9644
rect 10267 9636 10713 9644
rect 10727 9636 10853 9644
rect 2407 9616 3444 9624
rect 3696 9616 5213 9624
rect 1767 9596 2133 9604
rect 2276 9604 2284 9613
rect 3696 9604 3704 9616
rect 5827 9616 6433 9624
rect 7327 9616 7613 9624
rect 2276 9596 3704 9604
rect 4707 9596 4793 9604
rect 6607 9596 7773 9604
rect 8067 9596 8773 9604
rect 10467 9596 10733 9604
rect 10987 9596 11273 9604
rect 1467 9576 1553 9584
rect 1567 9576 1733 9584
rect 2967 9576 2993 9584
rect 3307 9576 3353 9584
rect 3767 9576 3913 9584
rect 3987 9576 4173 9584
rect 4227 9576 4373 9584
rect 4447 9576 5092 9584
rect 5127 9576 5653 9584
rect 5836 9576 6333 9584
rect 5836 9567 5844 9576
rect 6707 9576 7173 9584
rect 7447 9576 7693 9584
rect 8267 9576 8533 9584
rect 9027 9576 9273 9584
rect 9587 9576 9953 9584
rect 307 9556 393 9564
rect 3067 9556 3133 9564
rect 3387 9556 3733 9564
rect 4287 9556 4413 9564
rect 4627 9556 4713 9564
rect 4967 9556 5013 9564
rect 5727 9556 5833 9564
rect 8127 9556 8313 9564
rect 8327 9556 8453 9564
rect 9087 9556 9233 9564
rect 9427 9556 9473 9564
rect 9727 9556 9773 9564
rect 10600 9564 10613 9567
rect 10596 9556 10613 9564
rect 10600 9553 10613 9556
rect 10627 9556 10853 9564
rect 147 9537 173 9545
rect 227 9537 253 9545
rect 267 9536 373 9544
rect 447 9536 493 9544
rect 787 9537 833 9545
rect 1056 9524 1064 9534
rect 1147 9536 1253 9544
rect 1276 9536 1513 9544
rect 1276 9524 1284 9536
rect 1647 9536 2013 9544
rect 2027 9537 2093 9545
rect 2207 9536 2353 9544
rect 2873 9544 2887 9553
rect 2687 9536 2973 9544
rect 3407 9536 3513 9544
rect 3787 9536 3853 9544
rect 1056 9516 1284 9524
rect 347 9496 453 9504
rect 467 9495 513 9503
rect 907 9495 1133 9503
rect 1196 9496 1313 9504
rect 1196 9484 1204 9496
rect 1707 9495 1793 9503
rect 2347 9496 2653 9504
rect 3087 9496 3113 9504
rect 3287 9495 3373 9503
rect 3727 9496 3813 9504
rect 3976 9487 3984 9534
rect 4087 9536 4253 9544
rect 4507 9537 4733 9545
rect 5127 9537 5433 9545
rect 5667 9537 5693 9545
rect 6107 9537 6133 9545
rect 6487 9537 6513 9545
rect 6607 9537 6693 9545
rect 6947 9536 7053 9544
rect 4496 9524 4504 9534
rect 7247 9536 7373 9544
rect 7447 9536 7593 9544
rect 7647 9537 7672 9545
rect 7707 9536 7833 9544
rect 7847 9536 8093 9544
rect 8687 9536 8733 9544
rect 9027 9536 9264 9544
rect 4307 9516 4504 9524
rect 6387 9516 6873 9524
rect 6887 9516 6924 9524
rect 4247 9495 4273 9503
rect 4387 9495 4433 9503
rect 4807 9495 4933 9503
rect 5647 9496 5853 9504
rect 6127 9496 6193 9504
rect 6247 9495 6273 9503
rect 6547 9496 6593 9504
rect 6727 9496 6833 9504
rect 6916 9506 6924 9516
rect 7056 9516 8124 9524
rect 7056 9506 7064 9516
rect 8116 9506 8124 9516
rect 8227 9516 8433 9524
rect 9256 9506 9264 9536
rect 9507 9536 9853 9544
rect 9927 9537 10033 9545
rect 10127 9537 10173 9545
rect 10247 9537 10473 9545
rect 10487 9537 10573 9545
rect 7067 9495 7113 9503
rect 7227 9495 7353 9503
rect 7407 9495 7433 9503
rect 7547 9495 7613 9503
rect 7627 9496 7853 9504
rect 8467 9495 8513 9503
rect 8567 9495 8593 9503
rect 8667 9495 8753 9503
rect 8927 9495 8993 9503
rect 9427 9495 9512 9503
rect 9547 9496 9753 9504
rect 9867 9495 9933 9503
rect 10107 9496 10153 9504
rect 10167 9496 10593 9504
rect 10847 9495 11113 9503
rect 11127 9496 11153 9504
rect 1127 9476 1204 9484
rect 1367 9476 1873 9484
rect 3007 9476 3313 9484
rect 3427 9476 3513 9484
rect 4107 9476 4193 9484
rect 4987 9476 5053 9484
rect 5067 9476 5293 9484
rect 5347 9476 5393 9484
rect 5907 9476 6013 9484
rect 6347 9476 6473 9484
rect 9227 9476 10073 9484
rect 10527 9476 10553 9484
rect 867 9456 973 9464
rect 987 9456 1213 9464
rect 1547 9456 1753 9464
rect 1767 9456 2073 9464
rect 2467 9456 3393 9464
rect 3547 9456 3753 9464
rect 4487 9456 4513 9464
rect 4676 9456 4833 9464
rect 4676 9447 4684 9456
rect 4887 9456 4953 9464
rect 5467 9456 6133 9464
rect 6147 9456 7213 9464
rect 7527 9456 8253 9464
rect 8447 9456 8793 9464
rect 8807 9456 8833 9464
rect 8847 9456 9033 9464
rect 9807 9456 9993 9464
rect 10807 9456 11253 9464
rect 107 9436 633 9444
rect 647 9436 953 9444
rect 3467 9436 3533 9444
rect 4207 9436 4673 9444
rect 5167 9436 5193 9444
rect 5367 9436 5653 9444
rect 5807 9436 5913 9444
rect 6287 9436 6393 9444
rect 6567 9436 7173 9444
rect 9127 9436 9693 9444
rect 1247 9416 1273 9424
rect 4707 9416 4753 9424
rect 4987 9416 5273 9424
rect 5576 9416 6073 9424
rect 5576 9407 5584 9416
rect 6467 9416 6593 9424
rect 7827 9416 8293 9424
rect 10727 9416 11033 9424
rect 687 9396 773 9404
rect 787 9396 1013 9404
rect 1167 9396 1473 9404
rect 2936 9396 3144 9404
rect 2936 9384 2944 9396
rect 2307 9376 2944 9384
rect 3136 9384 3144 9396
rect 3507 9396 3553 9404
rect 3567 9396 3713 9404
rect 3767 9396 3833 9404
rect 4287 9396 4713 9404
rect 4727 9396 4813 9404
rect 4907 9396 5453 9404
rect 5467 9396 5573 9404
rect 5767 9396 5933 9404
rect 6967 9396 7913 9404
rect 9647 9396 10113 9404
rect 10127 9396 10393 9404
rect 3136 9376 3733 9384
rect 3927 9376 4253 9384
rect 5227 9376 5493 9384
rect 5707 9376 5904 9384
rect 587 9356 813 9364
rect 3147 9356 4693 9364
rect 4807 9356 5053 9364
rect 5107 9356 5873 9364
rect 5896 9364 5904 9376
rect 6107 9376 6313 9384
rect 6327 9376 6673 9384
rect 5896 9356 6293 9364
rect 7007 9356 8193 9364
rect 10927 9356 10953 9364
rect 1027 9336 1553 9344
rect 2007 9336 2313 9344
rect 2787 9336 2933 9344
rect 3847 9336 4173 9344
rect 4887 9336 4953 9344
rect 5227 9336 5533 9344
rect 5707 9336 5773 9344
rect 6387 9336 6713 9344
rect 7467 9336 8273 9344
rect 8287 9336 8453 9344
rect 11027 9336 11073 9344
rect 11087 9336 11273 9344
rect -63 9307 619 9315
rect 1007 9316 1913 9324
rect 3667 9316 3793 9324
rect 4027 9316 4293 9324
rect 4847 9316 5053 9324
rect 5867 9316 6913 9324
rect 8087 9316 8113 9324
rect 9747 9316 9913 9324
rect 9927 9316 10033 9324
rect 10047 9316 10313 9324
rect -63 9256 173 9264
rect 316 9236 413 9244
rect 316 9224 324 9236
rect 467 9237 493 9245
rect 611 9242 619 9307
rect 3207 9296 3593 9304
rect 4967 9296 5033 9304
rect 5087 9296 5153 9304
rect 5287 9296 5553 9304
rect 6187 9296 6513 9304
rect 6587 9296 7493 9304
rect 8647 9296 9193 9304
rect 9427 9296 9453 9304
rect 867 9276 1113 9284
rect 1927 9276 2033 9284
rect 2227 9276 2493 9284
rect 3627 9276 3913 9284
rect 4067 9276 4293 9284
rect 4507 9276 4693 9284
rect 4707 9276 4793 9284
rect 4847 9276 5253 9284
rect 5607 9276 5633 9284
rect 6007 9276 6553 9284
rect 7847 9276 7913 9284
rect 7927 9276 8413 9284
rect 8547 9276 8933 9284
rect 8947 9276 9013 9284
rect 9547 9276 9873 9284
rect 1447 9257 1613 9265
rect 2987 9256 3093 9264
rect 3107 9256 3173 9264
rect 4347 9256 4453 9264
rect 4827 9256 5093 9264
rect 5447 9256 5593 9264
rect 7907 9256 8073 9264
rect 9067 9256 9313 9264
rect 10787 9257 11073 9265
rect 611 9234 633 9242
rect 787 9236 893 9244
rect 907 9236 1353 9244
rect 2167 9237 2193 9245
rect 2236 9236 2253 9244
rect 127 9216 324 9224
rect 1527 9216 1653 9224
rect 1787 9217 1913 9225
rect 2236 9207 2244 9236
rect 2427 9237 2453 9245
rect 2727 9236 2873 9244
rect 2967 9237 3013 9245
rect 3327 9237 3373 9245
rect 3707 9237 3753 9245
rect 3216 9224 3224 9234
rect 3827 9236 4133 9244
rect 5247 9237 5333 9245
rect 5507 9237 5793 9245
rect 6187 9237 6473 9245
rect 6847 9237 6953 9245
rect 7107 9237 7133 9245
rect 7187 9236 7293 9244
rect 3216 9216 3664 9224
rect 347 9195 393 9203
rect 927 9195 1013 9203
rect 1067 9195 1093 9203
rect 1167 9196 1273 9204
rect 1387 9195 1413 9203
rect 2367 9195 2473 9203
rect 3027 9196 3193 9204
rect 3287 9195 3473 9203
rect 3547 9196 3633 9204
rect 3656 9204 3664 9216
rect 4307 9216 4484 9224
rect 4476 9207 4484 9216
rect 3656 9196 3713 9204
rect 3767 9196 4153 9204
rect 4207 9195 4233 9203
rect 4347 9196 4373 9204
rect 4476 9196 4493 9207
rect 4480 9193 4493 9196
rect 4676 9204 4684 9214
rect 4547 9196 4684 9204
rect 1487 9176 1573 9184
rect 1687 9176 1953 9184
rect 2127 9176 2272 9184
rect 2307 9176 2733 9184
rect 3127 9176 3153 9184
rect 3807 9176 3913 9184
rect 227 9156 873 9164
rect 2947 9156 3273 9164
rect 3447 9156 3613 9164
rect 3687 9156 3713 9164
rect 4367 9156 4433 9164
rect 607 9136 653 9144
rect 1587 9136 2053 9144
rect 2427 9136 2693 9144
rect 2707 9136 3433 9144
rect 3487 9136 3553 9144
rect 3947 9136 4533 9144
rect 687 9116 1333 9124
rect 2027 9116 2213 9124
rect 2627 9116 2693 9124
rect 3107 9116 3413 9124
rect 3587 9116 3653 9124
rect 3787 9116 3893 9124
rect 4696 9124 4704 9213
rect 4807 9196 4913 9204
rect 5087 9196 5233 9204
rect 5367 9196 5432 9204
rect 5467 9195 5533 9203
rect 5747 9195 5773 9203
rect 5836 9204 5844 9234
rect 7407 9236 7613 9244
rect 7967 9237 8033 9245
rect 8207 9237 8233 9245
rect 8427 9237 8493 9245
rect 8627 9237 8773 9245
rect 8927 9237 8973 9245
rect 9387 9237 9413 9245
rect 5816 9196 5844 9204
rect 5096 9176 5173 9184
rect 5096 9167 5104 9176
rect 5316 9184 5324 9192
rect 5316 9176 5424 9184
rect 4867 9156 5033 9164
rect 5087 9156 5104 9167
rect 5087 9153 5100 9156
rect 5307 9156 5393 9164
rect 5416 9164 5424 9176
rect 5487 9176 5573 9184
rect 5816 9167 5824 9196
rect 5887 9196 5993 9204
rect 6467 9196 6613 9204
rect 6707 9196 6853 9204
rect 6947 9196 7093 9204
rect 7356 9204 7364 9234
rect 8996 9216 9053 9224
rect 7167 9196 7364 9204
rect 7567 9195 7813 9203
rect 7867 9196 7953 9204
rect 8996 9206 9004 9216
rect 8627 9195 8673 9203
rect 9236 9204 9244 9234
rect 9567 9236 9653 9244
rect 10007 9237 10073 9245
rect 10127 9237 10253 9245
rect 10507 9237 10533 9245
rect 9016 9196 9473 9204
rect 5847 9176 6013 9184
rect 6247 9176 6333 9184
rect 7287 9176 7313 9184
rect 7587 9176 7673 9184
rect 8067 9176 8113 9184
rect 8527 9176 8913 9184
rect 9016 9184 9024 9196
rect 9487 9195 9553 9203
rect 9907 9196 9993 9204
rect 10047 9195 10133 9203
rect 11047 9196 11253 9204
rect 8927 9176 9024 9184
rect 9227 9176 9373 9184
rect 9420 9184 9433 9187
rect 9416 9173 9433 9184
rect 10336 9176 10733 9184
rect 5416 9156 5453 9164
rect 6027 9156 6113 9164
rect 6427 9156 6653 9164
rect 6667 9156 6753 9164
rect 6767 9156 6893 9164
rect 8447 9160 8684 9164
rect 8447 9156 8687 9160
rect 8673 9147 8687 9156
rect 9416 9164 9424 9173
rect 9007 9156 9424 9164
rect 10336 9164 10344 9176
rect 10067 9156 10344 9164
rect 10447 9156 10513 9164
rect 10527 9156 10593 9164
rect 5067 9136 5224 9144
rect 4696 9116 4753 9124
rect 4967 9116 5133 9124
rect 5216 9124 5224 9136
rect 7307 9136 7413 9144
rect 7427 9136 8013 9144
rect 8727 9136 9093 9144
rect 9727 9136 9893 9144
rect 10367 9136 11313 9144
rect 5216 9116 6833 9124
rect 8016 9124 8024 9133
rect 8016 9116 9133 9124
rect 9147 9116 9413 9124
rect 10047 9116 10673 9124
rect 10687 9116 10713 9124
rect 327 9096 433 9104
rect 1147 9096 1313 9104
rect 2367 9096 2393 9104
rect 2407 9096 3253 9104
rect 3347 9096 3393 9104
rect 3967 9096 4012 9104
rect 4047 9096 4173 9104
rect 4487 9096 4573 9104
rect 4807 9096 4933 9104
rect 5207 9096 5353 9104
rect 5527 9096 6373 9104
rect 7367 9096 8093 9104
rect 8567 9096 8733 9104
rect 9447 9096 9513 9104
rect 9587 9096 9693 9104
rect 9707 9096 10353 9104
rect 1787 9076 2333 9084
rect 2587 9076 3673 9084
rect 4247 9076 4673 9084
rect 5267 9076 6473 9084
rect 6527 9076 7273 9084
rect 7407 9076 7533 9084
rect 8667 9076 8693 9084
rect 767 9056 1093 9064
rect 1347 9056 1553 9064
rect 2807 9056 3293 9064
rect 4447 9056 4553 9064
rect 4993 9064 5007 9073
rect 4847 9056 5113 9064
rect 5607 9056 5633 9064
rect 5947 9056 6213 9064
rect 6307 9056 6393 9064
rect 7296 9056 7373 9064
rect 1147 9036 1273 9044
rect 1887 9036 1993 9044
rect 2067 9036 2533 9044
rect 3367 9036 3453 9044
rect 3707 9036 3773 9044
rect 3847 9036 4213 9044
rect 5407 9036 5853 9044
rect 7296 9044 7304 9056
rect 7987 9056 8313 9064
rect 9087 9056 9173 9064
rect 10347 9056 10633 9064
rect 7016 9036 7304 9044
rect 167 9016 213 9024
rect 747 9017 813 9025
rect 827 9016 1053 9024
rect 1067 9016 1413 9024
rect 1467 9016 1853 9024
rect 1867 9017 2033 9025
rect 2567 9016 2653 9024
rect 2707 9017 2753 9025
rect 2827 9016 2893 9024
rect 3387 9016 3513 9024
rect 3527 9016 3573 9024
rect 3747 9017 3813 9025
rect 3907 9016 4013 9024
rect 4067 9016 4244 9024
rect 127 8976 173 8984
rect 236 8967 244 8993
rect 276 8967 284 8994
rect 327 8995 453 9003
rect 4236 9004 4244 9016
rect 4267 9017 4393 9025
rect 4236 8996 4313 9004
rect 4476 9004 4484 9014
rect 4627 9016 4653 9024
rect 4927 9016 5073 9024
rect 4327 8996 4484 9004
rect 4696 9004 4704 9014
rect 5127 9017 5173 9025
rect 5247 9017 5393 9025
rect 5416 9016 5633 9024
rect 4696 8996 4813 9004
rect 5416 9004 5424 9016
rect 5947 9016 6313 9024
rect 6327 9017 6613 9025
rect 5376 8996 5424 9004
rect 847 8976 1073 8984
rect 1547 8976 1753 8984
rect 2027 8976 2073 8984
rect 2487 8975 2553 8983
rect 2747 8976 2793 8984
rect 3273 8984 3287 8993
rect 3273 8980 3373 8984
rect 3276 8976 3373 8980
rect 3447 8976 3553 8984
rect 3627 8975 3833 8983
rect 4007 8975 4113 8983
rect 4127 8975 4153 8983
rect 4167 8976 4353 8984
rect 5376 8986 5384 8996
rect 5896 8987 5904 9013
rect 7016 9006 7024 9036
rect 7667 9036 7813 9044
rect 8167 9036 8533 9044
rect 8667 9036 8973 9044
rect 10707 9036 10853 9044
rect 7387 9017 7453 9025
rect 7507 9016 7713 9024
rect 7727 9016 8253 9024
rect 9067 9016 9133 9024
rect 10607 9016 11013 9024
rect 11027 9017 11053 9025
rect 11107 9016 11173 9024
rect 7167 8997 7193 9005
rect 7267 8997 7293 9005
rect 8467 8997 8613 9005
rect 8707 9000 8864 9004
rect 8707 8996 8867 9000
rect 8853 8987 8867 8996
rect 8887 8996 8993 9004
rect 9087 8997 9113 9005
rect 9327 8995 9553 9003
rect 9607 8996 10053 9004
rect 4567 8975 4673 8983
rect 4947 8975 4993 8983
rect 5087 8975 5153 8983
rect 5207 8975 5273 8983
rect 5487 8975 5613 8983
rect 5627 8976 5764 8984
rect 276 8956 293 8967
rect 280 8953 293 8956
rect 627 8956 653 8964
rect 2787 8955 2953 8963
rect 3687 8956 4033 8964
rect 4107 8956 4413 8964
rect 4727 8956 4793 8964
rect 4807 8956 4913 8964
rect 5307 8956 5353 8964
rect 5756 8964 5764 8976
rect 6056 8976 6073 8984
rect 6056 8964 6064 8976
rect 6147 8976 6253 8984
rect 6487 8975 6813 8983
rect 7487 8976 7553 8984
rect 7827 8975 7893 8983
rect 8027 8975 8073 8983
rect 8127 8975 8153 8983
rect 8307 8976 8493 8984
rect 9596 8984 9604 8994
rect 10247 8995 10333 9003
rect 9456 8976 9604 8984
rect 5756 8956 6064 8964
rect 9456 8964 9464 8976
rect 10487 8975 10613 8983
rect 10667 8975 10693 8983
rect 10887 8975 10953 8983
rect 10967 8975 11013 8983
rect 9067 8956 9464 8964
rect 9487 8956 9933 8964
rect 11087 8956 11153 8964
rect 1047 8936 1073 8944
rect 1087 8936 1133 8944
rect 1347 8936 1833 8944
rect 1927 8936 1973 8944
rect 1987 8936 2213 8944
rect 2567 8936 2713 8944
rect 3307 8936 3393 8944
rect 3567 8936 3693 8944
rect 3767 8936 3893 8944
rect 4347 8936 4433 8944
rect 4627 8936 4893 8944
rect 4967 8936 5513 8944
rect 5647 8936 5833 8944
rect 5967 8936 6113 8944
rect 7307 8936 7593 8944
rect 8287 8936 8413 8944
rect 8587 8936 8953 8944
rect 227 8916 733 8924
rect 2527 8916 3113 8924
rect 4287 8916 4473 8924
rect 4867 8916 4993 8924
rect 5107 8916 5133 8924
rect 5267 8916 5493 8924
rect 6007 8916 6053 8924
rect 6067 8916 6513 8924
rect 6867 8916 7013 8924
rect 7027 8916 7513 8924
rect 7647 8916 7853 8924
rect 8627 8916 8713 8924
rect 9027 8916 9473 8924
rect 9787 8916 10093 8924
rect 2147 8896 2773 8904
rect 2867 8896 2973 8904
rect 3407 8896 3793 8904
rect 4547 8896 4733 8904
rect 5747 8896 5813 8904
rect 5887 8896 6373 8904
rect 7687 8896 8193 8904
rect 9976 8896 10833 8904
rect 9976 8887 9984 8896
rect 1387 8876 2433 8884
rect 2456 8876 2853 8884
rect 1327 8856 1433 8864
rect 1807 8856 1913 8864
rect 2456 8864 2464 8876
rect 2867 8876 3633 8884
rect 3647 8876 3733 8884
rect 3787 8876 3913 8884
rect 3927 8876 4213 8884
rect 4787 8876 5013 8884
rect 5227 8876 5724 8884
rect 2227 8856 2464 8864
rect 2547 8856 2713 8864
rect 2787 8856 3033 8864
rect 3147 8856 3493 8864
rect 3687 8856 4233 8864
rect 4887 8856 5033 8864
rect 5716 8864 5724 8876
rect 5987 8876 6193 8884
rect 6407 8876 7433 8884
rect 8327 8876 8533 8884
rect 9347 8876 9973 8884
rect 10847 8876 11113 8884
rect 5716 8856 6233 8864
rect 7467 8856 8693 8864
rect 8947 8856 9053 8864
rect 9407 8856 9633 8864
rect 527 8836 553 8844
rect 1247 8836 2493 8844
rect 2767 8836 3593 8844
rect 5287 8836 5933 8844
rect 6207 8836 6493 8844
rect 7287 8836 7773 8844
rect 8047 8836 8673 8844
rect 8727 8836 9113 8844
rect 10147 8836 10453 8844
rect 10647 8836 11173 8844
rect 2927 8816 3133 8824
rect 3227 8816 3573 8824
rect 3827 8816 3873 8824
rect 4507 8816 4953 8824
rect 5127 8816 5873 8824
rect 6007 8816 6293 8824
rect 6307 8816 6773 8824
rect 7027 8816 7053 8824
rect 7267 8816 8453 8824
rect 9933 8824 9947 8833
rect 9933 8820 10373 8824
rect 9936 8816 10373 8820
rect 2187 8796 2533 8804
rect 2547 8796 3173 8804
rect 3267 8796 4193 8804
rect 4827 8796 4893 8804
rect 4987 8796 6173 8804
rect 6227 8796 6293 8804
rect 7227 8796 8473 8804
rect 8707 8796 10033 8804
rect 1307 8776 1373 8784
rect 2287 8776 2473 8784
rect 3007 8776 3164 8784
rect 187 8756 333 8764
rect 467 8756 613 8764
rect 627 8756 1244 8764
rect 1236 8748 1244 8756
rect 2516 8756 2933 8764
rect 787 8736 813 8744
rect 1247 8737 1313 8745
rect 2516 8747 2524 8756
rect 3156 8764 3164 8776
rect 3287 8776 3413 8784
rect 3507 8776 3853 8784
rect 4287 8776 4933 8784
rect 5016 8776 5413 8784
rect 3156 8756 3213 8764
rect 3267 8756 3433 8764
rect 3607 8756 4393 8764
rect 4407 8756 4573 8764
rect 5016 8764 5024 8776
rect 5427 8776 6313 8784
rect 6927 8776 6984 8784
rect 4587 8756 5024 8764
rect 5436 8756 5584 8764
rect 1487 8736 1693 8744
rect 1787 8736 2353 8744
rect 2447 8736 2513 8744
rect 3387 8736 3493 8744
rect 3547 8736 3653 8744
rect 3807 8736 4593 8744
rect 4947 8736 5073 8744
rect 5436 8744 5444 8756
rect 5167 8736 5444 8744
rect 5576 8744 5584 8756
rect 5607 8756 6013 8764
rect 6976 8764 6984 8776
rect 7047 8776 7153 8784
rect 7167 8776 7713 8784
rect 7887 8776 7993 8784
rect 9027 8776 10433 8784
rect 6976 8756 7353 8764
rect 7527 8756 8333 8764
rect 8387 8756 8733 8764
rect 5576 8736 6073 8744
rect 6347 8736 6573 8744
rect 6587 8736 6873 8744
rect 6967 8736 7373 8744
rect 8187 8736 8312 8744
rect 8347 8737 8393 8745
rect 8787 8736 9173 8744
rect 9607 8736 9633 8744
rect 9647 8737 9713 8745
rect 10387 8737 10793 8745
rect 11267 8737 11293 8745
rect -63 8716 153 8724
rect 227 8716 373 8724
rect 2087 8717 2133 8725
rect 2147 8716 2273 8724
rect 2296 8716 2393 8724
rect 627 8697 753 8705
rect 1033 8704 1047 8713
rect 1033 8700 1353 8704
rect 1036 8696 1353 8700
rect 2296 8704 2304 8716
rect 2547 8717 2613 8725
rect 2667 8716 2893 8724
rect 3227 8717 3353 8725
rect 3447 8716 3633 8724
rect 3907 8717 3953 8725
rect 2156 8696 2304 8704
rect 2156 8686 2164 8696
rect 3956 8704 3964 8714
rect 4007 8716 4073 8724
rect 4116 8704 4124 8714
rect 4267 8716 4313 8724
rect 4356 8704 4364 8714
rect 4567 8716 4693 8724
rect 4707 8717 4793 8725
rect 4847 8717 4893 8725
rect 5447 8717 5553 8725
rect 5887 8716 6193 8724
rect 6707 8716 6753 8724
rect 2827 8696 3624 8704
rect 3956 8696 4364 8704
rect 867 8676 1073 8684
rect 2507 8676 2673 8684
rect 3047 8676 3113 8684
rect 3167 8675 3253 8683
rect 3427 8676 3533 8684
rect 3616 8686 3624 8696
rect 3807 8676 3873 8684
rect 4147 8675 4233 8683
rect 4396 8684 4404 8713
rect 4667 8696 4713 8704
rect 4727 8696 4804 8704
rect 4396 8676 4573 8684
rect 4747 8676 4773 8684
rect 4796 8684 4804 8696
rect 5016 8704 5024 8713
rect 4947 8696 5024 8704
rect 4796 8676 4813 8684
rect 4867 8676 4913 8684
rect 5016 8684 5024 8696
rect 5516 8696 5744 8704
rect 5016 8676 5053 8684
rect 5516 8684 5524 8696
rect 5156 8676 5524 8684
rect 1287 8656 1633 8664
rect 1727 8656 1933 8664
rect 1947 8656 2413 8664
rect 2707 8656 2913 8664
rect 3307 8656 3353 8664
rect 3527 8656 3653 8664
rect 3907 8656 3953 8664
rect 4107 8656 4273 8664
rect 4847 8656 4973 8664
rect 5156 8664 5164 8676
rect 5547 8676 5633 8684
rect 5736 8686 5744 8696
rect 5907 8676 5973 8684
rect 6147 8676 6213 8684
rect 6347 8675 6433 8683
rect 6456 8667 6464 8714
rect 7207 8716 7293 8724
rect 7407 8716 7533 8724
rect 7707 8717 7833 8725
rect 7916 8716 8453 8724
rect 7916 8704 7924 8716
rect 8467 8716 8513 8724
rect 8567 8717 8593 8725
rect 8927 8717 8973 8725
rect 9787 8716 9873 8724
rect 10287 8717 10313 8725
rect 6987 8696 7924 8704
rect 7947 8696 7973 8704
rect 8307 8696 8413 8704
rect 9627 8696 9753 8704
rect 10416 8696 10753 8704
rect 6527 8675 6673 8683
rect 6767 8675 6853 8683
rect 7007 8675 7093 8683
rect 7396 8676 7453 8684
rect 5127 8656 5164 8664
rect 5187 8656 5393 8664
rect 5747 8656 5773 8664
rect 7396 8664 7404 8676
rect 7547 8675 7593 8683
rect 7727 8676 7813 8684
rect 7827 8676 7993 8684
rect 8007 8676 8433 8684
rect 8447 8676 8493 8684
rect 8547 8676 8913 8684
rect 9047 8675 9193 8683
rect 9267 8676 9453 8684
rect 9467 8675 9573 8683
rect 10416 8684 10424 8696
rect 10947 8697 11093 8705
rect 11227 8696 11313 8704
rect 10307 8676 10424 8684
rect 11247 8676 11293 8684
rect 6947 8656 7404 8664
rect 7447 8656 7573 8664
rect 8607 8656 9033 8664
rect 9467 8656 9513 8664
rect 9767 8656 10393 8664
rect 11307 8656 11333 8664
rect 307 8636 793 8644
rect 807 8636 1173 8644
rect 1187 8636 1653 8644
rect 1676 8636 1873 8644
rect 1676 8624 1684 8636
rect 2127 8636 2313 8644
rect 3647 8636 3713 8644
rect 4147 8636 4352 8644
rect 4387 8636 4564 8644
rect 887 8616 1684 8624
rect 2207 8616 2673 8624
rect 2767 8616 3224 8624
rect 367 8596 413 8604
rect 427 8596 993 8604
rect 1007 8596 1893 8604
rect 1947 8596 2313 8604
rect 2327 8596 2693 8604
rect 2847 8596 3193 8604
rect 3216 8604 3224 8616
rect 3247 8616 3373 8624
rect 3747 8616 3873 8624
rect 3927 8616 4013 8624
rect 4087 8616 4413 8624
rect 4556 8624 4564 8636
rect 4596 8636 4893 8644
rect 4596 8624 4604 8636
rect 5067 8636 5413 8644
rect 5727 8636 6013 8644
rect 6387 8636 6513 8644
rect 6627 8636 8293 8644
rect 8807 8636 8853 8644
rect 10067 8636 10453 8644
rect 10467 8636 10913 8644
rect 4556 8616 4604 8624
rect 4707 8616 4813 8624
rect 4827 8616 4873 8624
rect 5087 8616 5213 8624
rect 5327 8616 5353 8624
rect 5447 8616 5533 8624
rect 6247 8616 6973 8624
rect 6996 8616 7073 8624
rect 3216 8596 3973 8604
rect 4107 8596 4173 8604
rect 4227 8596 4293 8604
rect 4367 8596 4393 8604
rect 4687 8596 5113 8604
rect 5407 8596 5873 8604
rect 6107 8596 6253 8604
rect 6996 8604 7004 8616
rect 7147 8616 7233 8624
rect 7627 8616 8033 8624
rect 8527 8616 8613 8624
rect 6427 8596 7004 8604
rect 7107 8596 7373 8604
rect 7387 8596 7493 8604
rect 7747 8596 7893 8604
rect 7907 8596 8324 8604
rect 207 8576 673 8584
rect 1367 8576 1533 8584
rect 1547 8576 1793 8584
rect 2287 8576 2753 8584
rect 2807 8576 3993 8584
rect 4207 8576 4653 8584
rect 4807 8576 4933 8584
rect 5367 8576 5833 8584
rect 6027 8576 6113 8584
rect 6256 8584 6264 8593
rect 8316 8587 8324 8596
rect 8347 8596 8804 8604
rect 6256 8576 6393 8584
rect 7187 8576 7353 8584
rect 7607 8576 7933 8584
rect 8327 8576 8593 8584
rect 8616 8576 8753 8584
rect 1087 8556 1933 8564
rect 2116 8556 2193 8564
rect 347 8536 453 8544
rect 467 8536 633 8544
rect 647 8536 773 8544
rect 2116 8544 2124 8556
rect 2387 8556 2493 8564
rect 2687 8556 4953 8564
rect 5027 8556 5273 8564
rect 5427 8556 5844 8564
rect 1447 8536 2124 8544
rect 2927 8536 3073 8544
rect 3087 8536 3292 8544
rect 3327 8536 3833 8544
rect 3987 8536 4253 8544
rect 4527 8536 4913 8544
rect 5047 8536 5133 8544
rect 5247 8536 5393 8544
rect 5836 8544 5844 8556
rect 5867 8556 6353 8564
rect 7287 8556 7453 8564
rect 8616 8564 8624 8576
rect 8796 8584 8804 8596
rect 8887 8596 9752 8604
rect 9787 8596 9953 8604
rect 10247 8596 11133 8604
rect 8796 8576 9673 8584
rect 10467 8576 10533 8584
rect 10867 8576 11053 8584
rect 8547 8556 8624 8564
rect 5836 8536 5953 8544
rect 6007 8536 6052 8544
rect 6087 8536 6293 8544
rect 6487 8536 6973 8544
rect 7547 8536 8333 8544
rect 10007 8536 10233 8544
rect 2647 8516 2793 8524
rect 3287 8516 3413 8524
rect 3467 8516 3553 8524
rect 3747 8516 4493 8524
rect 4567 8516 5013 8524
rect 5227 8516 5373 8524
rect 7307 8516 8433 8524
rect 9547 8516 9573 8524
rect 9587 8516 9753 8524
rect 9767 8516 10344 8524
rect 10336 8508 10344 8516
rect 10467 8516 10573 8524
rect 247 8496 413 8504
rect 1007 8497 1073 8505
rect 1127 8496 1313 8504
rect 1467 8497 1573 8505
rect 1627 8496 1733 8504
rect 1927 8497 1953 8505
rect 2407 8497 2453 8505
rect 2867 8496 3153 8504
rect 787 8476 1433 8484
rect 2176 8484 2184 8494
rect 3756 8496 3773 8504
rect 2176 8476 2373 8484
rect 3756 8484 3764 8496
rect 3827 8496 3853 8504
rect 3927 8497 3973 8505
rect 3996 8496 4013 8504
rect 3607 8476 3764 8484
rect 3996 8484 4004 8496
rect 4027 8496 4132 8504
rect 4167 8496 4233 8504
rect 3887 8476 4004 8484
rect 4456 8484 4464 8494
rect 4547 8496 4973 8504
rect 5067 8496 5133 8504
rect 5147 8496 5204 8504
rect 4456 8476 4773 8484
rect 4867 8476 5033 8484
rect 5196 8484 5204 8496
rect 5647 8497 5713 8505
rect 5767 8497 5813 8505
rect 5827 8496 6093 8504
rect 6207 8497 6233 8505
rect 6487 8496 6504 8504
rect 5196 8476 5293 8484
rect 907 8456 993 8464
rect 1107 8456 1153 8464
rect 1567 8456 1753 8464
rect 1767 8456 1913 8464
rect 1987 8456 2073 8464
rect 2167 8455 2313 8463
rect 2447 8456 2533 8464
rect 2667 8456 2693 8464
rect 2887 8455 2913 8463
rect 3467 8455 3493 8463
rect 4047 8455 4113 8463
rect 4487 8455 4533 8463
rect 4647 8456 4753 8464
rect 5427 8456 5453 8464
rect 6436 8464 6444 8493
rect 6496 8467 6504 8496
rect 6587 8496 7033 8504
rect 7227 8497 7273 8505
rect 7720 8504 7733 8507
rect 7716 8493 7733 8504
rect 7787 8496 8232 8504
rect 8267 8496 8413 8504
rect 8467 8496 8893 8504
rect 9447 8497 9493 8505
rect 9627 8496 9713 8504
rect 9907 8497 9993 8505
rect 10127 8497 10193 8505
rect 10347 8497 10413 8505
rect 10607 8496 10853 8504
rect 11067 8497 11093 8505
rect 6767 8475 6893 8483
rect 6947 8476 7033 8484
rect 6436 8456 6453 8464
rect 6916 8456 7053 8464
rect 127 8436 433 8444
rect 447 8436 973 8444
rect 1227 8436 1373 8444
rect 2847 8436 2973 8444
rect 2987 8436 3093 8444
rect 3387 8436 3413 8444
rect 3427 8436 3533 8444
rect 4207 8436 4453 8444
rect 5327 8436 5353 8444
rect 5727 8436 5853 8444
rect 6916 8446 6924 8456
rect 7127 8455 7233 8463
rect 7716 8466 7724 8493
rect 7527 8455 7673 8463
rect 667 8416 813 8424
rect 1407 8416 1633 8424
rect 1647 8416 2393 8424
rect 2587 8416 2693 8424
rect 3927 8416 4153 8424
rect 4207 8416 4553 8424
rect 4927 8416 5153 8424
rect 5607 8416 5873 8424
rect 7756 8424 7764 8474
rect 7867 8475 7993 8483
rect 8396 8476 8433 8484
rect 8396 8466 8404 8476
rect 8526 8473 8527 8480
rect 8547 8475 8673 8483
rect 8513 8467 8527 8473
rect 9007 8475 9133 8483
rect 10496 8467 10504 8474
rect 8513 8466 8540 8467
rect 8327 8455 8353 8463
rect 8513 8460 8533 8466
rect 8515 8456 8533 8460
rect 8520 8453 8533 8456
rect 9527 8456 9733 8464
rect 9787 8455 9873 8463
rect 9987 8456 10213 8464
rect 10487 8456 10504 8467
rect 10573 8464 10587 8473
rect 10573 8460 10733 8464
rect 10576 8456 10733 8460
rect 10487 8453 10500 8456
rect 8167 8436 8253 8444
rect 8267 8436 8833 8444
rect 8847 8436 9293 8444
rect 9307 8435 9353 8443
rect 7687 8416 7764 8424
rect 8867 8416 9573 8424
rect 1307 8396 1613 8404
rect 1847 8396 2193 8404
rect 3067 8396 3133 8404
rect 3147 8396 3233 8404
rect 4247 8396 4653 8404
rect 4947 8396 5253 8404
rect 5327 8396 5573 8404
rect 6047 8396 6193 8404
rect 6527 8396 6613 8404
rect 7207 8396 7313 8404
rect 7407 8396 7553 8404
rect 8147 8396 9332 8404
rect 9367 8396 9493 8404
rect 10187 8396 10473 8404
rect 2387 8376 2613 8384
rect 3627 8376 4024 8384
rect 1307 8356 1333 8364
rect 1467 8356 2293 8364
rect 2507 8356 2773 8364
rect 3347 8356 3753 8364
rect 4016 8364 4024 8376
rect 4047 8376 4353 8384
rect 4467 8376 4793 8384
rect 5287 8376 5453 8384
rect 5587 8376 5693 8384
rect 5887 8376 5993 8384
rect 6487 8376 7133 8384
rect 7647 8376 7833 8384
rect 8507 8376 8873 8384
rect 9527 8376 9893 8384
rect 4016 8356 4433 8364
rect 4887 8356 5113 8364
rect 5827 8356 5913 8364
rect 6387 8356 7373 8364
rect 7587 8356 8273 8364
rect 10707 8356 10833 8364
rect 247 8336 953 8344
rect 2467 8336 3253 8344
rect 3847 8336 4373 8344
rect 4387 8336 4733 8344
rect 4907 8336 4993 8344
rect 5167 8336 5713 8344
rect 5727 8336 5773 8344
rect 6756 8336 7033 8344
rect 327 8316 353 8324
rect 707 8316 1093 8324
rect 3287 8316 3404 8324
rect 376 8300 493 8304
rect 373 8296 493 8300
rect 373 8287 387 8296
rect 507 8296 533 8304
rect 2247 8296 2553 8304
rect 3207 8296 3333 8304
rect 3396 8304 3404 8316
rect 3807 8316 4313 8324
rect 4327 8316 4813 8324
rect 4827 8316 4873 8324
rect 5387 8316 6113 8324
rect 6756 8324 6764 8336
rect 7087 8336 7933 8344
rect 8487 8336 8713 8344
rect 6347 8316 6764 8324
rect 7147 8316 7533 8324
rect 7807 8316 7893 8324
rect 9207 8316 9464 8324
rect 3396 8296 3813 8304
rect 3947 8296 4193 8304
rect 4356 8296 5013 8304
rect 427 8276 1653 8284
rect 1807 8276 1933 8284
rect 2236 8284 2244 8293
rect 1947 8276 2244 8284
rect 2407 8276 3273 8284
rect 3907 8276 4253 8284
rect 4356 8284 4364 8296
rect 5107 8296 5413 8304
rect 5527 8296 5613 8304
rect 5896 8296 5973 8304
rect 4307 8276 4364 8284
rect 4407 8276 5053 8284
rect 5307 8276 5633 8284
rect 5896 8284 5904 8296
rect 6407 8296 6813 8304
rect 6947 8296 7293 8304
rect 7507 8296 8193 8304
rect 8207 8296 8333 8304
rect 8687 8296 8993 8304
rect 9007 8296 9433 8304
rect 9456 8304 9464 8316
rect 9507 8316 9593 8324
rect 9607 8316 9813 8324
rect 9827 8316 9853 8324
rect 10647 8316 11113 8324
rect 9456 8296 9613 8304
rect 9987 8296 10013 8304
rect 10027 8296 10393 8304
rect 5647 8276 5904 8284
rect 5967 8276 6273 8284
rect 6367 8276 8133 8284
rect 8547 8276 8853 8284
rect 10667 8276 10753 8284
rect 3707 8256 4213 8264
rect 4227 8256 5084 8264
rect 827 8236 1433 8244
rect 1487 8236 1853 8244
rect 2767 8236 3253 8244
rect 3407 8236 3833 8244
rect 4187 8236 4573 8244
rect 4707 8236 4833 8244
rect 4847 8236 4973 8244
rect 5076 8244 5084 8256
rect 5627 8256 5733 8264
rect 6807 8256 7013 8264
rect 7427 8256 7593 8264
rect 8467 8256 9393 8264
rect 10016 8256 10793 8264
rect 10016 8247 10024 8256
rect 5076 8236 5373 8244
rect 6187 8236 6253 8244
rect 6647 8236 7033 8244
rect 7126 8233 7127 8240
rect 7147 8236 7513 8244
rect 8807 8236 8913 8244
rect 9616 8236 10013 8244
rect 2207 8216 2313 8224
rect 3067 8217 3093 8225
rect 447 8196 653 8204
rect 707 8196 893 8204
rect 907 8196 933 8204
rect 1307 8197 1413 8205
rect 1487 8196 1513 8204
rect 1767 8197 1793 8205
rect 1987 8197 2073 8205
rect 2167 8196 2333 8204
rect 2347 8197 2373 8205
rect 2427 8196 2444 8204
rect 2436 8167 2444 8196
rect 2627 8196 2664 8204
rect 2656 8186 2664 8196
rect 2736 8187 2744 8213
rect 3307 8216 3892 8224
rect 3927 8216 4093 8224
rect 5116 8216 5153 8224
rect 3527 8196 3753 8204
rect 3767 8196 3884 8204
rect 3876 8184 3884 8196
rect 4187 8196 4213 8204
rect 4467 8196 4493 8204
rect 4887 8197 4933 8205
rect 5116 8204 5124 8216
rect 5196 8220 5573 8224
rect 5193 8216 5573 8220
rect 5067 8196 5124 8204
rect 5193 8207 5207 8216
rect 5727 8216 5893 8224
rect 5987 8216 6253 8224
rect 6267 8216 6333 8224
rect 7113 8224 7127 8233
rect 7027 8220 7127 8224
rect 7027 8216 7123 8220
rect 7187 8216 7253 8224
rect 7547 8217 7593 8225
rect 8607 8216 8753 8224
rect 9616 8224 9624 8236
rect 10247 8236 10444 8244
rect 9307 8216 9624 8224
rect 9636 8216 9893 8224
rect 5707 8197 5833 8205
rect 5967 8197 6053 8205
rect 6667 8197 6713 8205
rect 6867 8196 6904 8204
rect 2907 8176 2924 8184
rect 3876 8176 3913 8184
rect 227 8155 293 8163
rect 467 8155 553 8163
rect 1087 8156 1313 8164
rect 1867 8156 1953 8164
rect 2916 8164 2924 8176
rect 2916 8156 3033 8164
rect 3207 8156 3273 8164
rect 3327 8155 3393 8163
rect 3447 8155 3493 8163
rect 3547 8156 3613 8164
rect 3707 8155 3733 8163
rect 3996 8164 4004 8193
rect 6896 8187 6904 8196
rect 8167 8196 8393 8204
rect 8647 8196 8873 8204
rect 6656 8176 6793 8184
rect 3967 8156 4004 8164
rect 4027 8155 4133 8163
rect 4287 8155 4493 8163
rect 4867 8156 5044 8164
rect 296 8144 304 8152
rect 5036 8147 5044 8156
rect 5087 8156 5153 8164
rect 5267 8156 5333 8164
rect 6656 8164 6664 8176
rect 6896 8176 6913 8187
rect 6900 8173 6913 8176
rect 6647 8156 6664 8164
rect 6687 8156 6833 8164
rect 7067 8155 7113 8163
rect 7276 8164 7284 8194
rect 8947 8196 9024 8204
rect 7447 8176 7573 8184
rect 9016 8186 9024 8196
rect 9636 8204 9644 8216
rect 10436 8224 10444 8236
rect 10527 8236 10633 8244
rect 10887 8236 11233 8244
rect 10436 8216 10533 8224
rect 10547 8216 10673 8224
rect 10900 8224 10913 8227
rect 10896 8213 10913 8224
rect 11060 8224 11073 8227
rect 11056 8213 11073 8224
rect 9407 8196 9644 8204
rect 10067 8196 10084 8204
rect 7276 8156 7313 8164
rect 7696 8164 7704 8174
rect 7947 8175 8093 8183
rect 8967 8175 8992 8183
rect 9667 8177 9753 8185
rect 7696 8156 8133 8164
rect 8387 8156 8613 8164
rect 8667 8155 8833 8163
rect 9027 8156 9473 8164
rect 9787 8156 9953 8164
rect 9996 8164 10004 8193
rect 10076 8184 10084 8196
rect 10107 8196 10173 8204
rect 10727 8196 10844 8204
rect 10076 8176 10213 8184
rect 10836 8186 10844 8196
rect 10896 8184 10904 8213
rect 11056 8204 11064 8213
rect 10916 8200 11064 8204
rect 10867 8176 10904 8184
rect 10913 8196 11064 8200
rect 10913 8187 10927 8196
rect 9996 8156 10033 8164
rect 10056 8160 10073 8164
rect 10053 8156 10073 8160
rect 10053 8147 10067 8156
rect 10087 8156 10193 8164
rect 10547 8155 10573 8163
rect 10707 8155 10733 8163
rect 296 8136 413 8144
rect 427 8136 673 8144
rect 1767 8136 1793 8144
rect 2327 8140 2424 8144
rect 2327 8136 2427 8140
rect 2413 8127 2427 8136
rect 3947 8136 3973 8144
rect 5036 8136 5053 8147
rect 5040 8133 5053 8136
rect 5267 8136 5593 8144
rect 5747 8136 5873 8144
rect 6627 8136 6953 8144
rect 7067 8136 7353 8144
rect 7947 8136 7973 8144
rect 8307 8136 8853 8144
rect 8907 8136 9913 8144
rect 10527 8136 10933 8144
rect 11076 8144 11084 8174
rect 11207 8176 11313 8184
rect 11076 8136 11104 8144
rect 967 8116 1273 8124
rect 1287 8116 1473 8124
rect 1667 8116 1733 8124
rect 1827 8116 2273 8124
rect 2527 8116 2633 8124
rect 2707 8116 3013 8124
rect 3107 8116 3413 8124
rect 3507 8116 3873 8124
rect 3967 8116 4204 8124
rect 4196 8107 4204 8116
rect 4247 8116 4913 8124
rect 4987 8116 5193 8124
rect 5427 8116 5713 8124
rect 5727 8116 5753 8124
rect 5907 8116 5953 8124
rect 6067 8116 6153 8124
rect 6287 8116 6433 8124
rect 6556 8116 6933 8124
rect 887 8096 893 8104
rect 907 8096 2433 8104
rect 4196 8096 4213 8107
rect 4200 8093 4213 8096
rect 4507 8096 5313 8104
rect 5327 8096 5353 8104
rect 5547 8096 6033 8104
rect 6556 8104 6564 8116
rect 7007 8116 7413 8124
rect 7427 8116 7513 8124
rect 8847 8116 8913 8124
rect 8927 8116 9393 8124
rect 10687 8116 10893 8124
rect 11096 8124 11104 8136
rect 11207 8136 11293 8144
rect 11096 8116 11253 8124
rect 6187 8096 6564 8104
rect 6607 8096 6673 8104
rect 6847 8096 6873 8104
rect 6887 8096 7133 8104
rect 7287 8096 7393 8104
rect 8187 8096 8413 8104
rect 8767 8096 8804 8104
rect 147 8076 393 8084
rect 616 8076 853 8084
rect 616 8064 624 8076
rect 1367 8076 1533 8084
rect 1547 8076 2312 8084
rect 2347 8076 2413 8084
rect 3027 8076 3112 8084
rect 3147 8076 3193 8084
rect 3207 8076 3293 8084
rect 3727 8076 4173 8084
rect 4847 8076 4933 8084
rect 5067 8076 5293 8084
rect 5527 8076 5552 8084
rect 5587 8076 5973 8084
rect 6087 8076 6513 8084
rect 6827 8076 7013 8084
rect 7267 8076 7353 8084
rect 7407 8076 7753 8084
rect 7807 8076 7873 8084
rect 8107 8076 8373 8084
rect 8796 8084 8804 8096
rect 9387 8096 9413 8104
rect 10027 8096 10073 8104
rect 10207 8096 10693 8104
rect 10787 8096 10913 8104
rect 8796 8076 8873 8084
rect 9707 8076 9753 8084
rect 9807 8076 9872 8084
rect 9907 8076 10053 8084
rect 10387 8076 10713 8084
rect 10867 8076 10893 8084
rect 187 8056 624 8064
rect 1707 8056 1853 8064
rect 1927 8056 2013 8064
rect 2607 8056 2924 8064
rect 227 8036 553 8044
rect 636 8024 644 8053
rect 2916 8047 2924 8056
rect 2967 8056 3493 8064
rect 3507 8056 3633 8064
rect 3867 8056 4033 8064
rect 4207 8056 4613 8064
rect 4967 8056 5133 8064
rect 5367 8056 5393 8064
rect 5847 8056 5933 8064
rect 6247 8056 6473 8064
rect 6927 8056 7373 8064
rect 7387 8056 7593 8064
rect 7747 8056 7833 8064
rect 8807 8056 8893 8064
rect 9487 8056 9753 8064
rect 1527 8036 2093 8044
rect 2147 8036 2833 8044
rect 2916 8036 2933 8047
rect 2920 8033 2933 8036
rect 2987 8036 3713 8044
rect 3767 8036 3813 8044
rect 3876 8036 3993 8044
rect 3876 8027 3884 8036
rect 4267 8036 4553 8044
rect 4787 8036 5173 8044
rect 5936 8044 5944 8053
rect 5936 8036 6173 8044
rect 6713 8044 6727 8053
rect 9927 8056 10073 8064
rect 10327 8056 10353 8064
rect 10367 8056 10493 8064
rect 10507 8056 11293 8064
rect 6713 8040 7033 8044
rect 6716 8036 7033 8040
rect 7267 8036 7573 8044
rect 7967 8036 8193 8044
rect 8267 8036 9453 8044
rect 10556 8036 10873 8044
rect 10556 8027 10564 8036
rect 10887 8036 10933 8044
rect 10947 8036 11213 8044
rect 636 8016 664 8024
rect 367 7977 433 7985
rect 416 7956 513 7964
rect 416 7946 424 7956
rect 656 7966 664 8016
rect 2407 8016 2753 8024
rect 2767 8016 2793 8024
rect 3467 8016 3533 8024
rect 3867 8016 3884 8027
rect 3867 8013 3880 8016
rect 3947 8016 4764 8024
rect 1267 7996 1593 8004
rect 1667 7996 1993 8004
rect 2007 7996 2044 8004
rect 867 7976 1124 7984
rect 1116 7966 1124 7976
rect 1487 7977 1553 7985
rect 1687 7976 1813 7984
rect 2036 7984 2044 7996
rect 2087 7996 2344 8004
rect 2036 7976 2053 7984
rect 2187 7977 2233 7985
rect 2247 7977 2313 7985
rect 2336 7984 2344 7996
rect 3347 7996 3713 8004
rect 3787 7996 3833 8004
rect 3927 7996 4053 8004
rect 4307 7996 4393 8004
rect 4756 8004 4764 8016
rect 4816 8016 4973 8024
rect 4816 8007 4824 8016
rect 4987 8016 5033 8024
rect 5647 8016 5713 8024
rect 6107 8016 6173 8024
rect 6507 8016 6573 8024
rect 7127 8016 7633 8024
rect 7727 8016 7893 8024
rect 7907 8016 8233 8024
rect 8307 8016 8493 8024
rect 8507 8016 8812 8024
rect 8847 8016 9193 8024
rect 9607 8016 9853 8024
rect 9867 8016 10553 8024
rect 10607 8016 10693 8024
rect 4756 7996 4813 8004
rect 5427 7996 5613 8004
rect 2336 7976 2393 7984
rect 2507 7976 2533 7984
rect 2547 7976 2733 7984
rect 3087 7977 3133 7985
rect 3227 7977 3253 7985
rect 3967 7977 4033 7985
rect 4107 7977 4253 7985
rect 4407 7977 4473 7985
rect 4993 7984 5007 7993
rect 6047 7996 6473 8004
rect 6687 7996 7173 8004
rect 9427 7996 9824 8004
rect 9816 7988 9824 7996
rect 9947 7996 10773 8004
rect 10887 7996 11053 8004
rect 4947 7980 5007 7984
rect 4947 7976 5004 7980
rect 3736 7956 3853 7964
rect -63 7936 173 7944
rect 1627 7935 1673 7943
rect 2087 7935 2133 7943
rect 2407 7936 2513 7944
rect 2527 7936 2544 7944
rect 807 7916 853 7924
rect 867 7916 1313 7924
rect 1467 7916 1573 7924
rect 2347 7916 2373 7924
rect 2536 7924 2544 7936
rect 2947 7935 3013 7943
rect 3736 7946 3744 7956
rect 4716 7964 4724 7974
rect 5047 7976 5133 7984
rect 5187 7977 5273 7985
rect 5667 7976 5693 7984
rect 5867 7977 5913 7985
rect 6307 7976 6453 7984
rect 6567 7976 6633 7984
rect 6816 7976 6973 7984
rect 4087 7956 5053 7964
rect 5356 7947 5364 7973
rect 6816 7966 6824 7976
rect 7416 7964 7424 7974
rect 7467 7976 7773 7984
rect 7787 7977 7853 7985
rect 8287 7976 8373 7984
rect 8547 7976 8573 7984
rect 8767 7977 8833 7985
rect 8927 7977 8973 7985
rect 9027 7976 9093 7984
rect 9247 7977 9333 7985
rect 9387 7977 9453 7985
rect 9587 7977 9653 7985
rect 9827 7977 9853 7985
rect 10896 7976 11013 7984
rect 7416 7956 7684 7964
rect 3147 7936 3273 7944
rect 3527 7935 3693 7943
rect 3927 7935 3973 7943
rect 4027 7935 4053 7943
rect 4107 7935 4193 7943
rect 4567 7936 4813 7944
rect 4907 7936 5013 7944
rect 5087 7935 5153 7943
rect 5647 7936 5793 7944
rect 6207 7936 6313 7944
rect 7047 7936 7453 7944
rect 7616 7946 7624 7956
rect 7676 7944 7684 7956
rect 7676 7936 7833 7944
rect 8347 7936 8633 7944
rect 8827 7936 8953 7944
rect 9267 7936 9373 7944
rect 10116 7944 10124 7974
rect 10187 7956 10204 7964
rect 9536 7936 10153 7944
rect 2536 7916 2792 7924
rect 2827 7916 2853 7924
rect 4247 7916 4513 7924
rect 4527 7916 4853 7924
rect 5187 7916 5873 7924
rect 5987 7916 6053 7924
rect 6067 7916 6113 7924
rect 6547 7916 6813 7924
rect 7507 7916 7653 7924
rect 8227 7916 8313 7924
rect 8747 7916 8804 7924
rect 507 7896 953 7904
rect 1767 7896 1793 7904
rect 1807 7896 1833 7904
rect 1847 7896 2193 7904
rect 2267 7896 2893 7904
rect 3316 7896 3593 7904
rect 1427 7876 2073 7884
rect 3316 7884 3324 7896
rect 3827 7896 4033 7904
rect 4367 7896 4433 7904
rect 4447 7900 4524 7904
rect 4447 7896 4527 7900
rect 4513 7887 4527 7896
rect 4667 7896 4733 7904
rect 5367 7896 5413 7904
rect 5807 7896 5833 7904
rect 5967 7896 6093 7904
rect 6827 7896 7333 7904
rect 7787 7896 7873 7904
rect 8796 7904 8804 7916
rect 9067 7916 9293 7924
rect 9536 7924 9544 7936
rect 9347 7916 9544 7924
rect 9967 7916 10133 7924
rect 8796 7896 8993 7904
rect 9447 7896 9673 7904
rect 10136 7904 10144 7913
rect 10196 7904 10204 7956
rect 10287 7956 10532 7964
rect 10567 7964 10580 7967
rect 10567 7953 10584 7964
rect 10816 7964 10824 7974
rect 10896 7964 10904 7976
rect 10667 7956 10804 7964
rect 10816 7956 10904 7964
rect 10576 7926 10584 7953
rect 10796 7946 10804 7956
rect 10667 7916 10833 7924
rect 10136 7896 10204 7904
rect 11207 7896 11273 7904
rect 2907 7876 3324 7884
rect 3987 7876 4013 7884
rect 4187 7884 4200 7887
rect 4187 7873 4204 7884
rect 2387 7856 2753 7864
rect 2807 7856 3353 7864
rect 3367 7856 3753 7864
rect 3847 7856 4033 7864
rect 4196 7864 4204 7873
rect 4647 7876 4693 7884
rect 4827 7876 5172 7884
rect 5207 7876 5484 7884
rect 5476 7867 5484 7876
rect 7567 7876 7893 7884
rect 8367 7876 8773 7884
rect 9067 7876 9513 7884
rect 9707 7876 10013 7884
rect 10207 7876 11033 7884
rect 4196 7856 4293 7864
rect 4587 7856 5213 7864
rect 5487 7856 6393 7864
rect 6587 7856 6973 7864
rect 6987 7856 7253 7864
rect 8887 7856 9033 7864
rect 10647 7856 11253 7864
rect 1327 7836 2233 7844
rect 2487 7836 2653 7844
rect 3027 7836 3333 7844
rect 3487 7836 4133 7844
rect 4187 7836 4713 7844
rect 4827 7836 5273 7844
rect 5567 7836 6073 7844
rect 6487 7836 7433 7844
rect 7507 7836 8333 7844
rect 8347 7836 8433 7844
rect 8487 7836 9933 7844
rect 10007 7836 10413 7844
rect 10827 7836 11073 7844
rect 127 7816 893 7824
rect 2467 7816 2673 7824
rect 3807 7816 4184 7824
rect 4176 7807 4184 7816
rect 4347 7816 4553 7824
rect 4627 7816 4953 7824
rect 4967 7816 5033 7824
rect 5907 7816 6173 7824
rect 6487 7816 7313 7824
rect 7327 7816 7473 7824
rect 8087 7816 8453 7824
rect 10607 7816 10693 7824
rect 927 7796 1933 7804
rect 2607 7796 2633 7804
rect 2647 7796 2813 7804
rect 2947 7796 3473 7804
rect 3867 7796 4073 7804
rect 4187 7796 4493 7804
rect 5147 7796 6353 7804
rect 6407 7796 8473 7804
rect 9047 7796 9313 7804
rect 10027 7796 10093 7804
rect 10107 7796 10193 7804
rect 10207 7796 10313 7804
rect 10487 7796 10873 7804
rect 287 7776 1853 7784
rect 1867 7776 2033 7784
rect 2107 7776 2593 7784
rect 427 7756 493 7764
rect 507 7756 633 7764
rect 907 7756 1553 7764
rect 1567 7756 1713 7764
rect 2036 7764 2044 7773
rect 2667 7776 2873 7784
rect 2927 7776 3753 7784
rect 3916 7776 4353 7784
rect 3916 7764 3924 7776
rect 4667 7776 5073 7784
rect 5127 7776 5633 7784
rect 5647 7776 6093 7784
rect 6407 7776 7092 7784
rect 7127 7776 8293 7784
rect 8367 7776 8533 7784
rect 8547 7776 9573 7784
rect 9976 7776 10464 7784
rect 9976 7767 9984 7776
rect 2036 7756 3924 7764
rect 4027 7756 4053 7764
rect 4387 7756 4873 7764
rect 5067 7756 6213 7764
rect 6227 7756 6313 7764
rect 6327 7756 6373 7764
rect 6467 7756 6633 7764
rect 6647 7756 6673 7764
rect 8067 7756 8133 7764
rect 8327 7756 9973 7764
rect 10456 7764 10464 7776
rect 10456 7756 10693 7764
rect 207 7736 453 7744
rect 467 7736 673 7744
rect 2207 7736 2913 7744
rect 3947 7736 4133 7744
rect 4447 7736 4793 7744
rect 5767 7736 6173 7744
rect 6447 7736 6533 7744
rect 6887 7736 6933 7744
rect 6947 7736 7393 7744
rect 7807 7736 8113 7744
rect 8287 7736 9253 7744
rect 1287 7716 1773 7724
rect 2007 7716 2313 7724
rect 2556 7716 2773 7724
rect 2556 7707 2564 7716
rect 2827 7716 2973 7724
rect 4367 7716 5133 7724
rect 5367 7716 5473 7724
rect 5667 7716 5833 7724
rect 6367 7716 6593 7724
rect 6807 7716 7113 7724
rect 7707 7716 8253 7724
rect 8307 7716 8993 7724
rect 9827 7716 10193 7724
rect 1587 7696 1613 7704
rect 2047 7696 2093 7704
rect 2447 7696 2553 7704
rect 3207 7696 3353 7704
rect 3407 7697 3453 7705
rect 4287 7696 4313 7704
rect 6087 7696 6133 7704
rect 6147 7696 6233 7704
rect 6907 7696 7073 7704
rect 8487 7696 8513 7704
rect 9247 7696 9313 7704
rect 9627 7696 9733 7704
rect 267 7676 433 7684
rect 447 7676 873 7684
rect 987 7677 1033 7685
rect 1327 7677 1433 7685
rect 2007 7677 2073 7685
rect 2227 7676 2633 7684
rect 2707 7676 2893 7684
rect 3127 7676 3153 7684
rect 4087 7676 4433 7684
rect 4507 7677 4573 7685
rect 4767 7677 5113 7685
rect 5287 7676 5313 7684
rect 5407 7677 5433 7685
rect 5607 7676 5793 7684
rect 5987 7676 6013 7684
rect 6267 7677 6352 7685
rect 6387 7677 6433 7685
rect 6847 7677 6973 7685
rect 7047 7677 7133 7685
rect 7187 7677 7233 7685
rect 7407 7676 7433 7684
rect 3267 7656 3433 7664
rect 227 7635 253 7643
rect 347 7635 413 7643
rect 867 7636 973 7644
rect 1347 7636 1573 7644
rect 1947 7635 1973 7643
rect 2327 7636 2533 7644
rect 2627 7635 2693 7643
rect 2787 7635 2833 7643
rect 3247 7636 3333 7644
rect 3556 7644 3564 7654
rect 3807 7655 3933 7663
rect 6476 7664 6484 7674
rect 7487 7676 7593 7684
rect 7687 7677 7793 7685
rect 7847 7677 7913 7685
rect 8027 7677 8093 7685
rect 8567 7676 8693 7684
rect 8967 7676 9033 7684
rect 9087 7676 9153 7684
rect 10407 7676 10612 7684
rect 10647 7677 10733 7685
rect 10827 7684 10840 7687
rect 10827 7673 10844 7684
rect 6456 7656 6484 7664
rect 3556 7636 3693 7644
rect 4307 7635 4513 7643
rect 4747 7635 4813 7643
rect 4887 7636 5153 7644
rect 5167 7636 5193 7644
rect 5387 7636 5413 7644
rect 5587 7635 5633 7643
rect 5707 7636 5773 7644
rect 5827 7636 5893 7644
rect 6287 7636 6373 7644
rect 6456 7644 6464 7656
rect 6427 7636 6464 7644
rect 6507 7635 6533 7643
rect 6967 7636 7033 7644
rect 7227 7636 7253 7644
rect 7827 7636 7873 7644
rect 8247 7636 8373 7644
rect 8507 7635 8573 7643
rect 8727 7636 8793 7644
rect 8896 7644 8904 7673
rect 9307 7657 9453 7665
rect 9587 7656 9673 7664
rect 9896 7656 10013 7664
rect 8896 7636 8933 7644
rect 9067 7636 9133 7644
rect 9147 7635 9193 7643
rect 9896 7644 9904 7656
rect 10836 7666 10844 7673
rect 10927 7657 11073 7665
rect 11207 7656 11293 7664
rect 9716 7636 9904 7644
rect 1707 7616 1773 7624
rect 2747 7616 2873 7624
rect 3087 7616 3173 7624
rect 3447 7616 3993 7624
rect 4267 7616 4353 7624
rect 4847 7616 4933 7624
rect 5367 7616 5533 7624
rect 5647 7616 5673 7624
rect 5927 7616 6013 7624
rect 6787 7616 7193 7624
rect 7207 7616 7233 7624
rect 7467 7616 7593 7624
rect 7907 7616 8053 7624
rect 8067 7616 8173 7624
rect 8256 7616 8453 7624
rect 367 7596 473 7604
rect 567 7596 1293 7604
rect 1767 7596 2013 7604
rect 2347 7596 2593 7604
rect 2767 7596 3153 7604
rect 3167 7596 3733 7604
rect 4027 7596 4473 7604
rect 4587 7596 4693 7604
rect 4987 7596 5233 7604
rect 5427 7596 5513 7604
rect 6107 7596 6793 7604
rect 7236 7604 7244 7613
rect 7236 7596 7673 7604
rect 8256 7604 8264 7616
rect 8847 7616 8913 7624
rect 9327 7616 9593 7624
rect 9716 7624 9724 7636
rect 10147 7635 10333 7643
rect 10347 7636 10473 7644
rect 10707 7635 10753 7643
rect 9607 7616 9724 7624
rect 8147 7596 8264 7604
rect 8287 7596 8333 7604
rect 9007 7596 9204 7604
rect 1107 7576 1373 7584
rect 1927 7576 1973 7584
rect 2127 7576 2253 7584
rect 2807 7576 2873 7584
rect 3027 7576 3293 7584
rect 3767 7576 3973 7584
rect 4056 7576 4453 7584
rect 667 7556 973 7564
rect 1907 7556 3493 7564
rect 4056 7564 4064 7576
rect 4527 7576 4653 7584
rect 4847 7576 4953 7584
rect 6207 7576 6493 7584
rect 7387 7576 7493 7584
rect 7567 7576 7713 7584
rect 8587 7576 8933 7584
rect 9107 7576 9173 7584
rect 9196 7584 9204 7596
rect 9747 7596 9852 7604
rect 9887 7596 9993 7604
rect 10207 7596 10484 7604
rect 9196 7576 10053 7584
rect 10107 7576 10293 7584
rect 10476 7584 10484 7596
rect 10687 7596 10893 7604
rect 10476 7576 10533 7584
rect 3807 7556 4064 7564
rect 4087 7556 4413 7564
rect 4767 7556 5093 7564
rect 5227 7556 5793 7564
rect 7167 7556 7313 7564
rect 7927 7556 8073 7564
rect 8167 7556 8373 7564
rect 8427 7556 8513 7564
rect 8607 7556 8753 7564
rect 9547 7556 9893 7564
rect 10467 7556 10573 7564
rect 10887 7556 10953 7564
rect 1367 7536 1433 7544
rect 1747 7536 2012 7544
rect 2047 7536 2073 7544
rect 2247 7536 2513 7544
rect 2607 7536 2853 7544
rect 3707 7536 4013 7544
rect 4467 7536 5333 7544
rect 5987 7536 6573 7544
rect 6727 7536 6913 7544
rect 7247 7536 7573 7544
rect 7587 7536 7693 7544
rect 7707 7536 7893 7544
rect 8067 7536 8093 7544
rect 9047 7536 9213 7544
rect 9287 7536 9393 7544
rect 9407 7536 9753 7544
rect 9767 7536 10213 7544
rect 10387 7536 10493 7544
rect 10907 7536 10944 7544
rect 787 7516 1033 7524
rect 1587 7516 2213 7524
rect 2587 7516 3173 7524
rect 3187 7516 3433 7524
rect 3787 7516 3953 7524
rect 4007 7516 4393 7524
rect 4647 7516 4713 7524
rect 4867 7516 4993 7524
rect 5087 7516 5653 7524
rect 5847 7516 5913 7524
rect 6187 7516 6564 7524
rect 407 7493 413 7507
rect 587 7496 813 7504
rect 1067 7496 1233 7504
rect 1247 7496 1533 7504
rect 2547 7496 2753 7504
rect 2767 7496 3053 7504
rect 3487 7496 3813 7504
rect 3987 7496 4033 7504
rect 4047 7496 4073 7504
rect 4167 7496 4473 7504
rect 4487 7496 4653 7504
rect 4807 7496 5973 7504
rect 6556 7504 6564 7516
rect 6607 7516 7113 7524
rect 7427 7516 7473 7524
rect 8127 7516 8293 7524
rect 8647 7516 9313 7524
rect 9327 7516 9673 7524
rect 10307 7516 10673 7524
rect 10847 7516 10893 7524
rect 10936 7524 10944 7536
rect 10936 7516 10973 7524
rect 6556 7496 7273 7504
rect 7327 7496 7533 7504
rect 7547 7496 7573 7504
rect 7587 7496 8453 7504
rect 8727 7496 8833 7504
rect 8847 7496 8973 7504
rect 9727 7496 9793 7504
rect 10156 7496 11053 7504
rect 1047 7476 1393 7484
rect 1407 7476 1484 7484
rect 187 7457 253 7465
rect 467 7457 593 7465
rect 616 7456 633 7464
rect 616 7444 624 7456
rect 867 7457 893 7465
rect 1087 7457 1113 7465
rect 1476 7464 1484 7476
rect 1727 7476 1853 7484
rect 2067 7476 2153 7484
rect 2227 7476 2633 7484
rect 2647 7476 3793 7484
rect 4047 7476 4093 7484
rect 5207 7476 5533 7484
rect 7407 7476 7433 7484
rect 7767 7476 7813 7484
rect 8387 7476 8553 7484
rect 9087 7476 9133 7484
rect 9267 7476 9493 7484
rect 10156 7484 10164 7496
rect 9507 7476 10164 7484
rect 10267 7476 10453 7484
rect 10547 7476 10633 7484
rect 10647 7476 10853 7484
rect 10867 7476 11013 7484
rect 1476 7456 1493 7464
rect 1647 7457 1693 7465
rect 1927 7457 1953 7465
rect 2987 7456 3233 7464
rect 3307 7457 3333 7465
rect 3567 7456 3604 7464
rect 596 7436 624 7444
rect 2136 7436 2213 7444
rect 207 7416 333 7424
rect 347 7416 373 7424
rect 427 7415 493 7423
rect 596 7407 604 7436
rect 627 7416 833 7424
rect 967 7416 1293 7424
rect 2136 7426 2144 7436
rect 2267 7435 2353 7443
rect 2627 7436 3284 7444
rect 1807 7416 1893 7424
rect 2647 7416 2813 7424
rect 3276 7426 3284 7436
rect 3596 7427 3604 7456
rect 3996 7427 4004 7454
rect 4427 7456 4633 7464
rect 5047 7456 5173 7464
rect 5227 7456 5253 7464
rect 5887 7457 5973 7465
rect 6227 7456 6313 7464
rect 6316 7436 6353 7444
rect 2867 7416 3013 7424
rect 3287 7415 3533 7423
rect 3987 7416 4004 7427
rect 3987 7413 4000 7416
rect 4027 7415 4093 7423
rect 4167 7415 4373 7423
rect 4387 7415 4453 7423
rect 4467 7416 4673 7424
rect 4747 7415 4833 7423
rect 5007 7415 5033 7423
rect 5407 7416 5493 7424
rect 5507 7416 5653 7424
rect 5787 7416 5813 7424
rect 6316 7424 6324 7436
rect 6516 7444 6524 7454
rect 6567 7456 6653 7464
rect 6707 7457 6753 7465
rect 6767 7456 6833 7464
rect 6887 7457 6953 7465
rect 7007 7456 7373 7464
rect 6876 7444 6884 7454
rect 6367 7436 6524 7444
rect 6776 7436 6884 7444
rect 7413 7444 7427 7453
rect 7413 7440 7444 7444
rect 7416 7436 7444 7440
rect 6307 7416 6324 7424
rect 6567 7416 6613 7424
rect 6776 7426 6784 7436
rect 7436 7426 7444 7436
rect 6927 7415 7013 7423
rect 7456 7407 7464 7454
rect 7627 7456 7653 7464
rect 7733 7444 7747 7453
rect 7916 7456 8113 7464
rect 7676 7440 7747 7444
rect 7676 7436 7744 7440
rect 7756 7436 7793 7444
rect 7676 7426 7684 7436
rect 7756 7424 7764 7436
rect 7916 7446 7924 7456
rect 8407 7456 8473 7464
rect 7736 7420 7764 7424
rect 7733 7416 7764 7420
rect 7733 7407 7747 7416
rect 8076 7407 8084 7433
rect 1127 7396 1253 7404
rect 1267 7396 1433 7404
rect 2847 7396 3213 7404
rect 3227 7396 3293 7404
rect 3487 7396 3793 7404
rect 3807 7396 3893 7404
rect 4067 7396 4133 7404
rect 5927 7396 6052 7404
rect 6087 7396 6113 7404
rect 8356 7404 8364 7454
rect 8547 7456 8613 7464
rect 8667 7457 8693 7465
rect 8907 7457 9013 7465
rect 9067 7456 9173 7464
rect 9707 7456 9753 7464
rect 10187 7456 10293 7464
rect 11067 7457 11093 7465
rect 11107 7456 11193 7464
rect 11207 7456 11313 7464
rect 8567 7415 8593 7423
rect 8856 7424 8864 7453
rect 9840 7444 9853 7447
rect 9836 7433 9853 7444
rect 9893 7444 9907 7453
rect 9893 7440 9973 7444
rect 9896 7436 9973 7440
rect 8827 7416 8864 7424
rect 9087 7415 9213 7423
rect 9307 7416 9513 7424
rect 9567 7415 9693 7423
rect 8127 7396 8324 7404
rect 8356 7396 8413 7404
rect 987 7376 1473 7384
rect 1487 7376 1513 7384
rect 2567 7376 2593 7384
rect 2687 7376 2813 7384
rect 3367 7376 3573 7384
rect 4007 7376 4173 7384
rect 4667 7376 5133 7384
rect 5147 7376 5353 7384
rect 5447 7376 5773 7384
rect 5867 7376 6253 7384
rect 6507 7376 6813 7384
rect 7107 7376 7273 7384
rect 7367 7376 7493 7384
rect 7587 7376 7753 7384
rect 8107 7376 8213 7384
rect 8316 7384 8324 7396
rect 8647 7396 8713 7404
rect 9836 7406 9844 7433
rect 11027 7415 11073 7423
rect 10887 7396 11113 7404
rect 8316 7376 8473 7384
rect 9887 7376 10133 7384
rect 10267 7376 10444 7384
rect 487 7356 1053 7364
rect 1667 7356 1773 7364
rect 1816 7356 1944 7364
rect 1816 7344 1824 7356
rect 907 7336 1824 7344
rect 1936 7344 1944 7356
rect 2067 7356 2613 7364
rect 2807 7356 2893 7364
rect 3507 7356 4213 7364
rect 4367 7356 4692 7364
rect 4727 7356 4873 7364
rect 5287 7356 5373 7364
rect 5427 7356 5453 7364
rect 6067 7356 6253 7364
rect 6347 7356 6393 7364
rect 6467 7356 8253 7364
rect 8307 7356 8813 7364
rect 9707 7356 10393 7364
rect 10436 7364 10444 7376
rect 10436 7356 10673 7364
rect 10727 7356 11313 7364
rect 1936 7336 2093 7344
rect 2647 7336 3393 7344
rect 4647 7336 5033 7344
rect 5187 7336 5553 7344
rect 5947 7336 6273 7344
rect 6827 7336 7453 7344
rect 7527 7336 8113 7344
rect 8387 7336 8433 7344
rect 8787 7336 8893 7344
rect 9867 7336 10253 7344
rect 347 7316 1833 7324
rect 2247 7316 2524 7324
rect 1387 7296 1413 7304
rect 2347 7296 2493 7304
rect 2516 7304 2524 7316
rect 2656 7316 2993 7324
rect 2656 7304 2664 7316
rect 3967 7316 4493 7324
rect 4567 7316 5053 7324
rect 5107 7316 5333 7324
rect 6207 7316 6753 7324
rect 7147 7316 7573 7324
rect 8207 7316 9793 7324
rect 10607 7316 10753 7324
rect 2516 7296 2664 7304
rect 2887 7296 3973 7304
rect 5987 7296 6733 7304
rect 7227 7296 7513 7304
rect 8707 7296 8953 7304
rect 8967 7296 9613 7304
rect 10107 7296 10193 7304
rect 10207 7296 11113 7304
rect 287 7276 653 7284
rect 667 7276 1313 7284
rect 1367 7276 1433 7284
rect 3207 7276 3913 7284
rect 4687 7276 4833 7284
rect 5067 7276 7153 7284
rect 7387 7276 7513 7284
rect 8147 7276 8173 7284
rect 9747 7276 9853 7284
rect 10767 7276 10793 7284
rect 1547 7256 1692 7264
rect 1727 7256 1833 7264
rect 2707 7256 2933 7264
rect 3407 7256 3853 7264
rect 4867 7256 4993 7264
rect 5047 7256 5633 7264
rect 6167 7256 6313 7264
rect 6427 7256 6493 7264
rect 6727 7256 6893 7264
rect 7607 7256 7773 7264
rect 8427 7256 8824 7264
rect 1327 7236 1553 7244
rect 1567 7236 1673 7244
rect 1867 7236 2153 7244
rect 2587 7236 2953 7244
rect 3907 7236 4453 7244
rect 4627 7236 4852 7244
rect 4887 7236 6053 7244
rect 6147 7236 6293 7244
rect 6487 7236 6653 7244
rect 7127 7236 7193 7244
rect 7267 7236 7473 7244
rect 7487 7236 7713 7244
rect 7727 7236 8173 7244
rect 8816 7244 8824 7256
rect 8847 7256 8973 7264
rect 9047 7256 9773 7264
rect 9927 7256 10613 7264
rect 8816 7236 9053 7244
rect -63 7216 373 7224
rect 1247 7216 1733 7224
rect 3107 7216 3493 7224
rect 4487 7216 4793 7224
rect 4847 7216 5153 7224
rect 5547 7216 6033 7224
rect 6547 7216 6573 7224
rect 6587 7216 7013 7224
rect 8447 7216 9493 7224
rect 9567 7216 9813 7224
rect 10047 7216 10293 7224
rect 607 7196 653 7204
rect 1527 7196 1893 7204
rect 3227 7196 3453 7204
rect 3527 7196 3833 7204
rect 4307 7196 4913 7204
rect 5347 7196 6193 7204
rect 6267 7196 6524 7204
rect 1307 7177 1353 7185
rect 1367 7176 2193 7184
rect 2207 7176 2273 7184
rect 3067 7176 3344 7184
rect -63 7156 153 7164
rect 207 7157 273 7165
rect 627 7157 673 7165
rect 807 7156 1133 7164
rect 1687 7157 1773 7165
rect 1827 7156 1852 7164
rect 1887 7156 1993 7164
rect 2167 7156 2193 7164
rect 1267 7136 1373 7144
rect 2107 7136 2144 7144
rect 647 7116 793 7124
rect 867 7116 893 7124
rect 1407 7115 1493 7123
rect 1807 7116 1833 7124
rect 1907 7115 1973 7123
rect 2136 7124 2144 7136
rect 2307 7136 2333 7144
rect 2596 7144 2604 7173
rect 2787 7157 2873 7165
rect 2927 7157 2973 7165
rect 3067 7156 3113 7164
rect 3336 7164 3344 7176
rect 3887 7176 3953 7184
rect 4347 7176 4413 7184
rect 4467 7176 5253 7184
rect 5327 7176 5953 7184
rect 5967 7176 6133 7184
rect 6516 7184 6524 7196
rect 6616 7196 6773 7204
rect 6616 7187 6624 7196
rect 7407 7196 7453 7204
rect 10167 7196 10453 7204
rect 6516 7176 6613 7184
rect 6907 7176 6933 7184
rect 7116 7176 7593 7184
rect 3336 7156 3353 7164
rect 3467 7157 3633 7165
rect 4107 7157 4173 7165
rect 4867 7157 5033 7165
rect 5187 7157 5213 7165
rect 5527 7157 5573 7165
rect 5727 7156 5873 7164
rect 6087 7157 6173 7165
rect 6267 7157 6393 7165
rect 6667 7156 6853 7164
rect 6867 7157 6953 7165
rect 2596 7136 2613 7144
rect 2136 7116 2213 7124
rect 2127 7096 2313 7104
rect 1267 7076 1533 7084
rect 1707 7076 1753 7084
rect 2436 7084 2444 7134
rect 3727 7136 4153 7144
rect 2767 7115 2893 7123
rect 2947 7116 2993 7124
rect 3207 7115 3333 7123
rect 3387 7116 3513 7124
rect 3787 7115 3873 7123
rect 4356 7124 4364 7153
rect 4387 7135 4413 7143
rect 4327 7116 4364 7124
rect 3547 7096 3653 7104
rect 3987 7096 4033 7104
rect 4047 7096 4273 7104
rect 4616 7104 4624 7134
rect 4747 7136 4933 7144
rect 4956 7136 5004 7144
rect 4956 7124 4964 7136
rect 4756 7116 4964 7124
rect 4996 7124 5004 7136
rect 5476 7144 5484 7154
rect 5107 7136 5484 7144
rect 4996 7116 5013 7124
rect 4756 7104 4764 7116
rect 5196 7120 5233 7124
rect 5193 7116 5233 7120
rect 5193 7107 5207 7116
rect 5287 7115 5333 7123
rect 5407 7116 5533 7124
rect 5627 7116 5753 7124
rect 4616 7096 4764 7104
rect 4927 7096 4973 7104
rect 5916 7104 5924 7154
rect 6436 7144 6444 7154
rect 7027 7156 7053 7164
rect 6067 7136 6444 7144
rect 7056 7144 7064 7154
rect 7116 7144 7124 7176
rect 9127 7176 9164 7184
rect 7447 7157 7473 7165
rect 7056 7136 7124 7144
rect 8216 7127 8224 7154
rect 9107 7157 9133 7165
rect 8373 7144 8387 7153
rect 8373 7140 8493 7144
rect 8376 7136 8493 7140
rect 8536 7136 8613 7144
rect 5947 7116 6013 7124
rect 6427 7116 6553 7124
rect 6787 7115 6833 7123
rect 6927 7115 7153 7123
rect 7347 7115 7453 7123
rect 7547 7116 7573 7124
rect 7727 7115 7793 7123
rect 8027 7116 8073 7124
rect 8087 7116 8193 7124
rect 8216 7116 8233 7127
rect 8220 7113 8233 7116
rect 5807 7096 6093 7104
rect 6167 7096 6333 7104
rect 7507 7096 7833 7104
rect 8127 7096 8173 7104
rect 8267 7096 8333 7104
rect 8536 7104 8544 7136
rect 9156 7146 9164 7176
rect 9216 7176 9393 7184
rect 9216 7146 9224 7176
rect 9787 7176 9853 7184
rect 9927 7176 9953 7184
rect 9767 7156 9933 7164
rect 9267 7137 9393 7145
rect 10036 7124 10044 7153
rect 10436 7147 10444 7173
rect 10596 7147 10604 7173
rect 11167 7157 11233 7165
rect 11247 7154 11403 7168
rect 10027 7116 10044 7124
rect 10507 7116 10533 7124
rect 8507 7096 8544 7104
rect 8927 7096 9092 7104
rect 9127 7096 9253 7104
rect 9667 7096 9713 7104
rect 9727 7096 9773 7104
rect 9787 7096 9913 7104
rect 2127 7076 2444 7084
rect 2687 7076 2873 7084
rect 2967 7076 3053 7084
rect 3147 7076 3553 7084
rect 4127 7076 4793 7084
rect 4947 7076 5033 7084
rect 5267 7076 5353 7084
rect 5507 7076 5553 7084
rect 5827 7076 5872 7084
rect 5907 7076 5993 7084
rect 6207 7076 6273 7084
rect 6920 7084 6932 7087
rect 6916 7073 6932 7084
rect 6967 7076 7113 7084
rect 7227 7076 7373 7084
rect 7447 7076 7633 7084
rect 7647 7076 7753 7084
rect 7807 7076 7933 7084
rect 8807 7076 9213 7084
rect 9936 7076 10053 7084
rect 427 7056 793 7064
rect 1327 7056 1673 7064
rect 1687 7056 1873 7064
rect 2107 7056 2893 7064
rect 2947 7056 3212 7064
rect 3247 7056 3793 7064
rect 3987 7056 4812 7064
rect 4847 7056 5053 7064
rect 5387 7056 5473 7064
rect 5527 7056 5653 7064
rect 6307 7056 6353 7064
rect 6916 7064 6924 7073
rect 6407 7056 6924 7064
rect 7047 7056 7153 7064
rect 7247 7056 8393 7064
rect 9087 7056 9173 7064
rect 9936 7064 9944 7076
rect 10427 7076 10893 7084
rect 9747 7056 9944 7064
rect 507 7036 673 7044
rect 987 7036 1233 7044
rect 1247 7036 1273 7044
rect 1927 7036 2113 7044
rect 2176 7036 2924 7044
rect 2176 7027 2184 7036
rect 767 7016 1493 7024
rect 1507 7016 2173 7024
rect 2567 7016 2773 7024
rect 2916 7024 2924 7036
rect 2947 7036 3133 7044
rect 3327 7036 5453 7044
rect 5587 7036 5613 7044
rect 6036 7036 6073 7044
rect 2916 7016 3193 7024
rect 3547 7016 3573 7024
rect 3667 7016 4153 7024
rect 4247 7016 4373 7024
rect 4667 7016 4713 7024
rect 4807 7016 5173 7024
rect 6036 7024 6044 7036
rect 7287 7036 7433 7044
rect 7487 7036 8593 7044
rect 5707 7016 6044 7024
rect 6067 7016 6273 7024
rect 6347 7016 6633 7024
rect 6907 7016 7213 7024
rect 7387 7016 7453 7024
rect 7527 7016 7893 7024
rect 8507 7016 8573 7024
rect 9467 7016 9593 7024
rect 9987 7016 10253 7024
rect 10327 7016 10493 7024
rect 307 6996 693 7004
rect 807 6996 1453 7004
rect 1787 6996 1933 7004
rect 2927 6996 2973 7004
rect 3347 6996 3424 7004
rect 2027 6976 2233 6984
rect 2407 6976 2673 6984
rect 2727 6976 2933 6984
rect 3047 6976 3373 6984
rect 3416 6984 3424 6996
rect 3567 6996 4113 7004
rect 4847 6996 4933 7004
rect 5087 6996 5193 7004
rect 5207 7004 5220 7007
rect 5207 6996 5224 7004
rect 5207 6993 5220 6996
rect 5287 6996 5433 7004
rect 6047 6996 6153 7004
rect 6307 6996 6664 7004
rect 3416 6976 3613 6984
rect 4407 6976 4513 6984
rect 4747 6976 4953 6984
rect 5487 6976 5633 6984
rect 5987 6976 6333 6984
rect 6656 6984 6664 6996
rect 6767 6996 6833 7004
rect 6887 6996 7353 7004
rect 7727 6996 7793 7004
rect 8147 6996 8213 7004
rect 8227 6996 8293 7004
rect 8607 6996 9293 7004
rect 10607 6996 10713 7004
rect 10767 6996 10853 7004
rect 6656 6976 7473 6984
rect 7967 6976 8124 6984
rect 147 6956 173 6964
rect 287 6956 593 6964
rect 607 6956 1033 6964
rect 2307 6956 2693 6964
rect 2716 6956 3013 6964
rect 207 6936 233 6944
rect 787 6937 833 6945
rect 1016 6936 1073 6944
rect 300 6924 313 6927
rect 253 6904 267 6913
rect 227 6900 267 6904
rect 296 6913 313 6924
rect 227 6896 264 6900
rect 296 6887 304 6913
rect 1016 6907 1024 6936
rect 1127 6937 1253 6945
rect 1467 6936 1533 6944
rect 1667 6937 1733 6945
rect 2167 6937 2193 6945
rect 2327 6937 2453 6945
rect 347 6896 473 6904
rect 867 6896 973 6904
rect 296 6876 313 6887
rect 300 6873 313 6876
rect 1107 6876 1293 6884
rect 1447 6876 1513 6884
rect 1807 6876 1853 6884
rect 1976 6884 1984 6934
rect 2716 6944 2724 6956
rect 3707 6956 3853 6964
rect 4207 6956 4273 6964
rect 4387 6956 4693 6964
rect 4827 6956 4984 6964
rect 2627 6936 2724 6944
rect 2767 6936 2913 6944
rect 3236 6936 3333 6944
rect 2956 6907 2964 6934
rect 3236 6926 3244 6936
rect 3387 6936 3453 6944
rect 3567 6936 3613 6944
rect 4073 6944 4087 6953
rect 4073 6940 4124 6944
rect 4076 6936 4124 6940
rect 2407 6895 2433 6903
rect 2647 6895 2693 6903
rect 2956 6896 2973 6907
rect 2960 6893 2973 6896
rect 1976 6876 2013 6884
rect 2267 6876 2473 6884
rect 2527 6876 2573 6884
rect 2996 6884 3004 6914
rect 3767 6896 4033 6904
rect 4116 6887 4124 6936
rect 4333 6944 4347 6953
rect 4307 6940 4347 6944
rect 4307 6936 4344 6940
rect 4767 6936 4853 6944
rect 4556 6924 4564 6934
rect 4976 6944 4984 6956
rect 5047 6956 5273 6964
rect 5327 6956 5393 6964
rect 5587 6956 5633 6964
rect 5856 6956 5893 6964
rect 4976 6936 4993 6944
rect 5067 6936 5513 6944
rect 5856 6944 5864 6956
rect 5907 6956 6293 6964
rect 6427 6956 6473 6964
rect 6647 6956 6693 6964
rect 7087 6956 7293 6964
rect 7667 6956 7733 6964
rect 7787 6956 7993 6964
rect 8007 6956 8033 6964
rect 8116 6964 8124 6976
rect 8187 6976 8273 6984
rect 8827 6976 9073 6984
rect 9347 6976 9773 6984
rect 9827 6976 10133 6984
rect 10347 6976 10393 6984
rect 10467 6976 10593 6984
rect 8116 6956 8393 6964
rect 10187 6956 10273 6964
rect 10407 6956 10433 6964
rect 10456 6956 10564 6964
rect 5847 6936 5864 6944
rect 6087 6937 6113 6945
rect 6487 6936 6613 6944
rect 6807 6937 6893 6945
rect 6947 6936 6993 6944
rect 7047 6937 7093 6945
rect 7147 6937 7273 6945
rect 7347 6937 7453 6945
rect 7507 6936 7553 6944
rect 8527 6936 8613 6944
rect 8627 6936 8813 6944
rect 9107 6937 9153 6945
rect 9407 6936 9533 6944
rect 9587 6937 9673 6945
rect 9687 6936 9873 6944
rect 10456 6944 10464 6956
rect 9996 6936 10464 6944
rect 10556 6944 10564 6956
rect 10556 6936 10673 6944
rect 4316 6916 4784 6924
rect 4316 6906 4324 6916
rect 4776 6906 4784 6916
rect 4427 6895 4493 6903
rect 4547 6895 4593 6903
rect 4707 6895 4733 6903
rect 4787 6895 4913 6903
rect 5147 6895 5373 6903
rect 5527 6895 5613 6903
rect 5796 6904 5804 6933
rect 6256 6916 7024 6924
rect 5796 6896 5813 6904
rect 5987 6895 6013 6903
rect 6256 6904 6264 6916
rect 6067 6896 6264 6904
rect 6287 6896 6393 6904
rect 7016 6906 7024 6916
rect 6507 6895 6573 6903
rect 6627 6895 6693 6903
rect 6847 6895 6973 6903
rect 7236 6896 7253 6904
rect 2947 6876 3004 6884
rect 3607 6876 3713 6884
rect 4116 6876 4133 6887
rect 4120 6873 4133 6876
rect 5027 6876 5053 6884
rect 7236 6884 7244 6896
rect 7267 6896 7433 6904
rect 7567 6895 7693 6903
rect 8236 6904 8244 6933
rect 9996 6926 10004 6936
rect 8207 6896 8244 6904
rect 8327 6896 8413 6904
rect 8607 6896 8833 6904
rect 9087 6896 9313 6904
rect 9387 6895 9453 6903
rect 9467 6895 9553 6903
rect 9856 6887 9864 6913
rect 10236 6904 10244 6914
rect 10307 6916 10533 6924
rect 10236 6896 10393 6904
rect 10407 6895 10433 6903
rect 10607 6895 10653 6903
rect 10747 6896 11033 6904
rect 11047 6896 11153 6904
rect 11287 6896 11403 6904
rect 6607 6876 7244 6884
rect 8007 6876 8033 6884
rect 9367 6876 9393 6884
rect 707 6856 833 6864
rect 847 6856 953 6864
rect 1007 6856 1173 6864
rect 1567 6856 1993 6864
rect 2147 6856 2213 6864
rect 2227 6856 2533 6864
rect 3947 6856 4073 6864
rect 4227 6856 4693 6864
rect 5667 6856 6333 6864
rect 7107 6856 7333 6864
rect 7447 6856 7733 6864
rect 7747 6856 7973 6864
rect 10287 6856 10573 6864
rect 10587 6856 10913 6864
rect 10927 6856 10973 6864
rect 3067 6836 3633 6844
rect 4267 6836 4873 6844
rect 5027 6836 5393 6844
rect 5887 6836 6033 6844
rect 6047 6836 6373 6844
rect 6487 6836 6912 6844
rect 6947 6836 7213 6844
rect 7267 6836 8633 6844
rect 8647 6836 8853 6844
rect 8867 6836 9573 6844
rect 9767 6836 10293 6844
rect 1507 6816 1593 6824
rect 1767 6816 2073 6824
rect 2467 6816 2553 6824
rect 2667 6816 2733 6824
rect 3407 6816 3433 6824
rect 3447 6816 3533 6824
rect 3627 6816 3733 6824
rect 3947 6816 4193 6824
rect 4567 6816 4833 6824
rect 5287 6816 5613 6824
rect 6167 6816 6313 6824
rect 6796 6816 8533 6824
rect 2747 6796 2833 6804
rect 3447 6796 3593 6804
rect 3847 6796 4233 6804
rect 4307 6796 5013 6804
rect 6796 6804 6804 6816
rect 9827 6816 10313 6824
rect 10327 6816 10993 6824
rect 5207 6796 6804 6804
rect 7587 6796 7733 6804
rect 8967 6796 9353 6804
rect 9507 6796 9544 6804
rect 227 6776 493 6784
rect 3527 6776 4833 6784
rect 4847 6776 5293 6784
rect 5307 6776 6133 6784
rect 6347 6776 6613 6784
rect 6667 6776 6713 6784
rect 7427 6776 7933 6784
rect 8347 6776 8733 6784
rect 9536 6784 9544 6796
rect 9587 6796 10033 6804
rect 10047 6796 10253 6804
rect 9536 6776 10153 6784
rect 10167 6776 10573 6784
rect 10587 6776 10693 6784
rect 987 6756 1013 6764
rect 2407 6756 2553 6764
rect 2647 6756 2753 6764
rect 2767 6756 2913 6764
rect 3107 6756 3233 6764
rect 3327 6753 3333 6767
rect 3547 6756 3753 6764
rect 3907 6756 4133 6764
rect 4327 6756 4353 6764
rect 4907 6756 5013 6764
rect 5067 6756 5893 6764
rect 5967 6756 6253 6764
rect 6327 6756 6653 6764
rect 6976 6756 7053 6764
rect 647 6736 1133 6744
rect 3287 6736 3513 6744
rect 4067 6736 4273 6744
rect 5067 6736 5913 6744
rect 6367 6736 6592 6744
rect 6976 6744 6984 6756
rect 9487 6756 9513 6764
rect 6627 6736 6984 6744
rect 7027 6736 7473 6744
rect 8107 6736 8993 6744
rect 9007 6736 9113 6744
rect 9567 6736 9833 6744
rect 9847 6736 10133 6744
rect 10147 6736 10273 6744
rect 10627 6736 10693 6744
rect 2596 6716 4293 6724
rect 1847 6696 2153 6704
rect 2167 6696 2213 6704
rect 2596 6704 2604 6716
rect 4587 6716 4933 6724
rect 5087 6716 5173 6724
rect 5427 6716 5453 6724
rect 5627 6716 5893 6724
rect 5967 6716 6113 6724
rect 7067 6716 7353 6724
rect 9556 6724 9564 6733
rect 8607 6716 9564 6724
rect 11207 6716 11293 6724
rect 2467 6696 2604 6704
rect 3087 6696 3152 6704
rect 3187 6696 3573 6704
rect 3767 6696 4453 6704
rect 4667 6696 4753 6704
rect 4907 6696 5113 6704
rect 5387 6696 6473 6704
rect 7047 6696 7593 6704
rect 9047 6696 9113 6704
rect 9487 6696 9633 6704
rect 9647 6696 9713 6704
rect 10156 6696 10473 6704
rect 1667 6676 2353 6684
rect 2847 6676 3413 6684
rect 3576 6684 3584 6693
rect 3576 6676 4524 6684
rect 1147 6657 1193 6665
rect 1207 6657 1333 6665
rect 4516 6667 4524 6676
rect 4807 6676 5093 6684
rect 5107 6676 5193 6684
rect 5407 6676 5793 6684
rect 5847 6676 5933 6684
rect 5987 6676 6133 6684
rect 6147 6676 6193 6684
rect 7647 6676 7713 6684
rect 9387 6676 9713 6684
rect 10156 6684 10164 6696
rect 9927 6676 10164 6684
rect 2627 6656 2793 6664
rect 4516 6656 4533 6667
rect 4520 6653 4533 6656
rect 4827 6656 5273 6664
rect 5927 6656 6013 6664
rect 6027 6656 6353 6664
rect 6527 6656 6573 6664
rect 6947 6656 7033 6664
rect 8287 6656 8633 6664
rect 9707 6656 9753 6664
rect 10027 6656 10193 6664
rect 10287 6657 10633 6665
rect 11087 6656 11113 6664
rect 147 6637 233 6645
rect 387 6636 433 6644
rect 547 6636 633 6644
rect 676 6636 693 6644
rect 216 6616 333 6624
rect 216 6606 224 6616
rect 676 6624 684 6636
rect 1587 6636 1793 6644
rect 2087 6637 2413 6645
rect 2887 6637 2953 6645
rect 3107 6636 3153 6644
rect 3247 6637 3353 6645
rect 3687 6637 3753 6645
rect 4707 6637 4733 6645
rect 4787 6637 4893 6645
rect 5087 6637 5133 6645
rect 5207 6637 5373 6645
rect 5427 6637 5473 6645
rect 5727 6637 5873 6645
rect 5887 6636 6053 6644
rect 416 6616 684 6624
rect 416 6606 424 6616
rect 807 6616 833 6624
rect 1107 6616 1273 6624
rect 4053 6624 4067 6633
rect 4053 6620 4073 6624
rect 4056 6616 4073 6620
rect 4447 6616 4513 6624
rect 467 6596 493 6604
rect 507 6596 653 6604
rect 1387 6595 1413 6603
rect 1467 6595 1553 6603
rect 1787 6596 1913 6604
rect 2247 6595 2273 6603
rect 2367 6595 2393 6603
rect 2567 6595 2633 6603
rect 2987 6595 3273 6603
rect 3287 6595 3373 6603
rect 3427 6595 3573 6603
rect 3747 6595 3813 6603
rect 4687 6596 4793 6604
rect 4847 6595 4873 6603
rect 4927 6596 4973 6604
rect 5027 6596 5113 6604
rect 5407 6596 5453 6604
rect 5507 6595 5593 6603
rect 5656 6604 5664 6634
rect 6067 6636 6093 6644
rect 6247 6637 6313 6645
rect 6507 6637 6773 6645
rect 6816 6624 6824 6634
rect 6707 6616 6824 6624
rect 6976 6624 6984 6634
rect 6927 6616 6984 6624
rect 7467 6644 7480 6647
rect 7467 6633 7484 6644
rect 7947 6637 7973 6645
rect 8167 6640 8224 6644
rect 8167 6636 8227 6640
rect 7213 6624 7227 6633
rect 7213 6620 7333 6624
rect 7216 6616 7333 6620
rect 7356 6616 7433 6624
rect 5656 6596 5853 6604
rect 5907 6596 5953 6604
rect 5967 6596 6073 6604
rect 6127 6596 6233 6604
rect 6487 6595 6553 6603
rect 6667 6596 6833 6604
rect 2007 6576 2073 6584
rect 2807 6576 2913 6584
rect 3736 6584 3744 6592
rect 2927 6576 3744 6584
rect 4147 6576 4413 6584
rect 5027 6576 5153 6584
rect 5367 6576 5473 6584
rect 6327 6576 6373 6584
rect 7067 6576 7093 6584
rect 7356 6584 7364 6616
rect 7287 6576 7364 6584
rect 187 6556 253 6564
rect 2127 6556 2433 6564
rect 2547 6556 2633 6564
rect 3147 6556 3312 6564
rect 3347 6556 3533 6564
rect 4447 6556 4813 6564
rect 5547 6556 6073 6564
rect 6587 6556 6673 6564
rect 6727 6556 6753 6564
rect 6827 6556 6853 6564
rect 667 6536 1093 6544
rect 1107 6536 1593 6544
rect 1607 6536 1813 6544
rect 2567 6536 2673 6544
rect 2687 6536 2773 6544
rect 3136 6544 3144 6553
rect 2827 6536 3144 6544
rect 3307 6536 4013 6544
rect 5007 6536 5233 6544
rect 5307 6536 5353 6544
rect 6187 6536 6313 6544
rect 7476 6527 7484 6633
rect 8213 6627 8227 6636
rect 8827 6636 9053 6644
rect 9287 6636 9613 6644
rect 9807 6637 9953 6645
rect 9967 6636 10224 6644
rect 7667 6615 7693 6623
rect 7607 6596 7633 6604
rect 7647 6596 8013 6604
rect 8027 6596 8253 6604
rect 8436 6604 8444 6614
rect 9676 6624 9684 6634
rect 9547 6616 10073 6624
rect 10216 6624 10224 6636
rect 10867 6636 10933 6644
rect 10987 6636 11053 6644
rect 11167 6636 11273 6644
rect 11327 6636 11403 6644
rect 10216 6616 10233 6624
rect 10287 6617 10473 6625
rect 10607 6616 10673 6624
rect 11315 6624 11323 6633
rect 11236 6620 11323 6624
rect 11233 6616 11323 6620
rect 11233 6607 11247 6616
rect 8436 6596 8793 6604
rect 9007 6595 9033 6603
rect 9187 6596 9513 6604
rect 9667 6595 9813 6603
rect 9827 6595 9893 6603
rect 9947 6596 10012 6604
rect 10047 6595 10133 6603
rect 10947 6595 11073 6603
rect 8107 6576 8193 6584
rect 8876 6576 11213 6584
rect 7807 6556 8133 6564
rect 8876 6564 8884 6576
rect 11267 6576 11333 6584
rect 8547 6556 8884 6564
rect 8907 6556 9073 6564
rect 9507 6556 9693 6564
rect 10047 6556 10304 6564
rect 10296 6547 10304 6556
rect 10607 6556 10833 6564
rect 11107 6556 11293 6564
rect 8127 6536 8173 6544
rect 8987 6536 9053 6544
rect 10187 6536 10272 6544
rect 10307 6536 10913 6544
rect 10927 6536 11013 6544
rect 747 6516 773 6524
rect 787 6516 853 6524
rect 1007 6516 1173 6524
rect 1687 6516 2093 6524
rect 2107 6516 2273 6524
rect 2487 6516 3153 6524
rect 4056 6516 4124 6524
rect 987 6496 1073 6504
rect 2067 6496 2133 6504
rect 2407 6496 2833 6504
rect 2887 6496 2973 6504
rect 2987 6496 3173 6504
rect 3787 6496 3832 6504
rect 4056 6504 4064 6516
rect 3867 6496 4064 6504
rect 4116 6504 4124 6516
rect 4147 6516 4253 6524
rect 4407 6516 4693 6524
rect 4847 6516 5693 6524
rect 5807 6516 6413 6524
rect 6427 6516 6553 6524
rect 6807 6516 6913 6524
rect 7127 6516 7192 6524
rect 7227 6516 7353 6524
rect 7527 6516 7593 6524
rect 7847 6516 8033 6524
rect 9467 6516 9653 6524
rect 10507 6516 10733 6524
rect 10967 6516 11033 6524
rect 4116 6496 4233 6504
rect 5267 6496 5313 6504
rect 5547 6496 6633 6504
rect 6847 6496 7133 6504
rect 7507 6496 7813 6504
rect 7927 6496 9253 6504
rect 10587 6496 10693 6504
rect 367 6476 413 6484
rect 1507 6476 1833 6484
rect 1847 6476 1953 6484
rect 1967 6476 2453 6484
rect 2727 6476 2893 6484
rect 3007 6476 3193 6484
rect 3247 6476 4073 6484
rect 4476 6476 5073 6484
rect 347 6456 653 6464
rect 807 6456 1473 6464
rect 1487 6456 2493 6464
rect 2507 6456 3033 6464
rect 3047 6456 4133 6464
rect 4476 6464 4484 6476
rect 5127 6476 5933 6484
rect 6767 6476 6933 6484
rect 7147 6476 7433 6484
rect 8087 6476 8133 6484
rect 8587 6476 8833 6484
rect 9047 6476 9713 6484
rect 9807 6476 9973 6484
rect 10487 6476 10553 6484
rect 4247 6456 4484 6464
rect 5307 6456 5973 6464
rect 6447 6456 6613 6464
rect 6787 6456 6924 6464
rect 227 6436 313 6444
rect 1047 6436 1304 6444
rect 387 6417 453 6425
rect 587 6417 613 6425
rect 1187 6396 1272 6404
rect 1296 6406 1304 6436
rect 2647 6436 2804 6444
rect 1547 6416 1613 6424
rect 1627 6416 1713 6424
rect 1887 6417 1913 6425
rect 2107 6416 2133 6424
rect 2187 6417 2293 6425
rect 2627 6417 2753 6425
rect 2796 6424 2804 6436
rect 3547 6436 3573 6444
rect 3796 6436 3973 6444
rect 2796 6416 3033 6424
rect 3087 6417 3113 6425
rect 3136 6416 3153 6424
rect 2656 6396 2733 6404
rect 267 6376 393 6384
rect 407 6375 513 6383
rect 647 6376 1053 6384
rect 2167 6376 2473 6384
rect 2656 6384 2664 6396
rect 2807 6396 2993 6404
rect 2647 6376 2664 6384
rect 2687 6375 2713 6383
rect 2896 6386 2904 6396
rect 3136 6404 3144 6416
rect 3796 6424 3804 6436
rect 4307 6436 4573 6444
rect 4707 6436 5113 6444
rect 5227 6436 5393 6444
rect 5607 6436 6133 6444
rect 6467 6436 6733 6444
rect 6916 6444 6924 6456
rect 7167 6456 7272 6464
rect 7307 6456 7373 6464
rect 7567 6456 8053 6464
rect 9427 6456 9573 6464
rect 9627 6456 9893 6464
rect 9907 6456 10013 6464
rect 10707 6456 10733 6464
rect 6916 6436 7013 6444
rect 7367 6436 7513 6444
rect 8567 6436 8593 6444
rect 8847 6436 8973 6444
rect 9227 6436 9453 6444
rect 9467 6436 9533 6444
rect 3407 6416 3804 6424
rect 3827 6417 3953 6425
rect 3067 6396 3144 6404
rect 3196 6384 3204 6414
rect 4007 6416 4053 6424
rect 4107 6417 4153 6425
rect 4607 6417 4633 6425
rect 4727 6416 5093 6424
rect 5167 6417 5253 6425
rect 5327 6416 5433 6424
rect 6116 6416 6173 6424
rect 4507 6396 4873 6404
rect 3107 6376 3204 6384
rect 3887 6375 3993 6383
rect 4127 6375 4393 6383
rect 4587 6375 4673 6383
rect 4876 6384 4884 6393
rect 6116 6387 6124 6416
rect 6287 6416 6393 6424
rect 6627 6417 6773 6425
rect 6907 6416 7024 6424
rect 4876 6376 5173 6384
rect 5187 6376 5293 6384
rect 5747 6376 6092 6384
rect 7016 6386 7024 6416
rect 7047 6416 7333 6424
rect 7347 6417 7533 6425
rect 8127 6416 8273 6424
rect 8487 6417 8513 6425
rect 8536 6416 8553 6424
rect 7356 6396 7513 6404
rect 7356 6386 7364 6396
rect 7706 6393 7707 6400
rect 7727 6396 7973 6404
rect 8316 6404 8324 6414
rect 8536 6404 8544 6416
rect 8787 6417 8813 6425
rect 8887 6416 9173 6424
rect 9656 6416 9693 6424
rect 8316 6396 8544 6404
rect 6387 6375 6533 6383
rect 6647 6375 6933 6383
rect 7487 6376 7573 6384
rect 7693 6384 7707 6393
rect 7693 6380 7824 6384
rect 7696 6376 7824 6380
rect 1147 6355 1193 6363
rect 1747 6356 1873 6364
rect 1967 6356 2153 6364
rect 2387 6356 2412 6364
rect 2447 6356 2753 6364
rect 2767 6356 2873 6364
rect 3407 6356 3673 6364
rect 4207 6356 4773 6364
rect 4927 6356 5104 6364
rect 2287 6336 2564 6344
rect 187 6316 333 6324
rect 587 6316 1033 6324
rect 1107 6316 1733 6324
rect 2556 6324 2564 6336
rect 2607 6336 2633 6344
rect 2907 6336 3173 6344
rect 3187 6336 3313 6344
rect 3927 6336 4653 6344
rect 5096 6344 5104 6356
rect 5427 6356 5853 6364
rect 6347 6356 7233 6364
rect 7816 6364 7824 6376
rect 7847 6376 8113 6384
rect 8227 6375 8333 6383
rect 8487 6376 8673 6384
rect 8727 6375 8753 6383
rect 8807 6375 8833 6383
rect 9207 6376 9373 6384
rect 9387 6376 9433 6384
rect 9656 6384 9664 6416
rect 9707 6416 9793 6424
rect 9947 6416 10224 6424
rect 10216 6406 10224 6416
rect 10593 6424 10607 6433
rect 10547 6420 10607 6424
rect 10547 6416 10604 6420
rect 10627 6417 10733 6425
rect 10347 6396 10433 6404
rect 9487 6376 9664 6384
rect 10693 6384 10707 6393
rect 10527 6380 10707 6384
rect 10527 6376 10704 6380
rect 7816 6356 7993 6364
rect 9507 6356 9613 6364
rect 9627 6356 9873 6364
rect 10387 6356 10673 6364
rect 5096 6336 5813 6344
rect 5987 6336 6213 6344
rect 6236 6336 6493 6344
rect 1967 6316 2384 6324
rect 2556 6316 2593 6324
rect 1007 6296 1113 6304
rect 2167 6296 2193 6304
rect 2376 6304 2384 6316
rect 4047 6316 4433 6324
rect 4547 6316 4573 6324
rect 5087 6316 6033 6324
rect 6236 6324 6244 6336
rect 6507 6336 6873 6344
rect 6927 6336 7293 6344
rect 7407 6336 7433 6344
rect 7447 6336 7673 6344
rect 8927 6336 9733 6344
rect 6167 6316 6244 6324
rect 6267 6316 6333 6324
rect 8107 6316 8473 6324
rect 8907 6316 9353 6324
rect 9427 6316 9773 6324
rect 9827 6316 9893 6324
rect 10227 6316 10513 6324
rect 10727 6316 11233 6324
rect 2376 6296 3053 6304
rect 3307 6296 3453 6304
rect 3467 6296 3773 6304
rect 4147 6296 4384 6304
rect 1287 6276 1633 6284
rect 2047 6276 2833 6284
rect 3847 6276 3933 6284
rect 3947 6276 4353 6284
rect 4376 6284 4384 6296
rect 4787 6296 5893 6304
rect 6087 6296 6712 6304
rect 6747 6296 6972 6304
rect 7007 6296 7353 6304
rect 7527 6296 8073 6304
rect 9267 6296 10533 6304
rect 4376 6276 4913 6284
rect 5027 6276 5133 6284
rect 5896 6284 5904 6293
rect 5896 6276 7053 6284
rect 8967 6276 9053 6284
rect 9067 6276 9413 6284
rect 9787 6276 10173 6284
rect 10847 6276 10873 6284
rect 247 6256 573 6264
rect 1727 6256 2513 6264
rect 2527 6256 2853 6264
rect 3167 6256 3473 6264
rect 4407 6256 5533 6264
rect 5576 6256 5713 6264
rect 1467 6236 2193 6244
rect 2207 6236 3013 6244
rect 3607 6236 3733 6244
rect 4087 6236 4753 6244
rect 4767 6236 4953 6244
rect 5576 6244 5584 6256
rect 5787 6256 5873 6264
rect 5947 6256 6753 6264
rect 6767 6256 6953 6264
rect 7047 6256 7493 6264
rect 7547 6256 7753 6264
rect 7927 6256 8033 6264
rect 9447 6256 10273 6264
rect 10627 6256 11093 6264
rect 5287 6236 5584 6244
rect 5607 6236 6004 6244
rect 327 6216 704 6224
rect 696 6204 704 6216
rect 1627 6216 1913 6224
rect 2327 6216 2673 6224
rect 3067 6216 5473 6224
rect 5827 6216 5953 6224
rect 5996 6224 6004 6236
rect 6027 6236 6413 6244
rect 6727 6236 6913 6244
rect 7067 6236 7213 6244
rect 7407 6236 7653 6244
rect 8347 6236 8813 6244
rect 9147 6236 9233 6244
rect 9487 6236 9553 6244
rect 9567 6236 10373 6244
rect 5996 6216 6633 6224
rect 6747 6216 11233 6224
rect 696 6196 733 6204
rect 847 6196 973 6204
rect 987 6196 1293 6204
rect 1367 6196 1433 6204
rect 1527 6196 2033 6204
rect 2416 6196 2533 6204
rect 1296 6184 1304 6193
rect 1296 6176 1673 6184
rect 1687 6176 1953 6184
rect 2416 6184 2424 6196
rect 2547 6196 2733 6204
rect 2847 6196 4633 6204
rect 6107 6196 6353 6204
rect 6487 6196 6713 6204
rect 7247 6196 7553 6204
rect 7747 6196 7893 6204
rect 8767 6196 9113 6204
rect 9127 6196 9253 6204
rect 10087 6196 10653 6204
rect 10947 6196 11253 6204
rect 2167 6176 2424 6184
rect 2947 6176 3233 6184
rect 3787 6176 4133 6184
rect 4607 6176 4993 6184
rect 5307 6176 6053 6184
rect 6067 6176 6733 6184
rect 6927 6176 7133 6184
rect 8867 6176 9093 6184
rect 9547 6176 9853 6184
rect 11047 6176 11093 6184
rect 447 6156 633 6164
rect 647 6156 813 6164
rect 1207 6156 2133 6164
rect 2747 6156 2853 6164
rect 3027 6156 3093 6164
rect 3107 6156 3133 6164
rect 3267 6156 3373 6164
rect 3387 6156 3453 6164
rect 3467 6156 3713 6164
rect 6127 6160 6184 6164
rect 6127 6156 6187 6160
rect 707 6136 833 6144
rect 1827 6136 1893 6144
rect 2467 6136 2893 6144
rect -63 6116 173 6124
rect 367 6117 393 6125
rect 907 6116 1013 6124
rect 1027 6117 1073 6125
rect 1547 6117 1793 6125
rect 2153 6124 2167 6133
rect 3387 6136 3433 6144
rect 4727 6136 4913 6144
rect 5827 6137 5933 6145
rect 6173 6147 6187 6156
rect 6407 6156 6532 6164
rect 6567 6156 6793 6164
rect 6887 6156 7353 6164
rect 7367 6156 7553 6164
rect 7707 6156 7853 6164
rect 7967 6156 8113 6164
rect 8247 6156 8553 6164
rect 8967 6156 9033 6164
rect 9647 6156 9713 6164
rect 9907 6156 10193 6164
rect 10296 6156 10473 6164
rect 6927 6136 6953 6144
rect 9447 6137 9473 6145
rect 9687 6136 9813 6144
rect 9987 6136 10133 6144
rect 10296 6144 10304 6156
rect 10147 6136 10304 6144
rect 10827 6136 11033 6144
rect 1967 6120 2167 6124
rect 1967 6116 2164 6120
rect 2307 6116 2433 6124
rect 2696 6116 2773 6124
rect 1047 6096 1364 6104
rect 1356 6084 1364 6096
rect 1947 6096 2173 6104
rect 1356 6076 1373 6084
rect 1747 6075 1853 6083
rect 1867 6076 2033 6084
rect 467 6056 513 6064
rect 527 6056 693 6064
rect 1307 6036 1333 6044
rect 1447 6036 1733 6044
rect 1627 6016 2073 6024
rect 87 5996 593 6004
rect 607 5996 793 6004
rect 1336 5996 1513 6004
rect 1336 5987 1344 5996
rect 1527 5996 1593 6004
rect 2087 5996 2213 6004
rect 2276 6004 2284 6093
rect 2547 6076 2653 6084
rect 2696 6086 2704 6116
rect 2816 6104 2824 6114
rect 2947 6116 2973 6124
rect 3047 6116 3213 6124
rect 3227 6117 3553 6125
rect 4107 6116 4253 6124
rect 4467 6116 4553 6124
rect 5007 6117 5213 6125
rect 5227 6117 5333 6125
rect 5993 6124 6007 6133
rect 5387 6116 5424 6124
rect 5993 6120 6113 6124
rect 5996 6116 6113 6120
rect 2816 6096 2893 6104
rect 3787 6096 4193 6104
rect 5416 6106 5424 6116
rect 6487 6117 6613 6125
rect 6707 6116 6753 6124
rect 6827 6116 6893 6124
rect 7027 6117 7093 6125
rect 7187 6116 7213 6124
rect 7787 6117 7813 6125
rect 7867 6116 8033 6124
rect 8087 6117 8333 6125
rect 9007 6116 9044 6124
rect 4807 6096 5404 6104
rect 2767 6075 2933 6083
rect 3147 6075 3193 6083
rect 3287 6075 3433 6083
rect 3607 6076 3633 6084
rect 3827 6075 3893 6083
rect 4227 6076 4433 6084
rect 4567 6075 4633 6083
rect 5067 6076 5093 6084
rect 5107 6075 5153 6083
rect 5316 6080 5353 6084
rect 5313 6076 5353 6080
rect 5313 6067 5327 6076
rect 5396 6084 5404 6096
rect 5396 6076 5473 6084
rect 2907 6056 2993 6064
rect 3327 6056 3433 6064
rect 3547 6056 4013 6064
rect 4067 6056 4693 6064
rect 2687 6036 2793 6044
rect 3116 6036 3544 6044
rect 2507 6016 2533 6024
rect 2796 6024 2804 6033
rect 3116 6024 3124 6036
rect 2796 6016 3124 6024
rect 3347 6016 3453 6024
rect 3536 6024 3544 6036
rect 3567 6036 3693 6044
rect 3707 6036 3973 6044
rect 4147 6036 4173 6044
rect 4327 6036 4673 6044
rect 3536 6016 4113 6024
rect 4827 6016 5433 6024
rect 5656 6024 5664 6094
rect 5807 6096 5853 6104
rect 6987 6096 7293 6104
rect 7436 6087 7444 6114
rect 5867 6076 5933 6084
rect 6387 6076 6493 6084
rect 6767 6075 6873 6083
rect 6927 6076 7013 6084
rect 7207 6075 7333 6083
rect 7427 6076 7444 6087
rect 7496 6087 7504 6114
rect 9036 6106 9044 6116
rect 10067 6117 10093 6125
rect 10187 6116 10253 6124
rect 10267 6116 10313 6124
rect 10367 6116 10393 6124
rect 10467 6116 10633 6124
rect 10967 6117 10993 6125
rect 9127 6097 9273 6105
rect 9387 6096 9773 6104
rect 9833 6104 9847 6113
rect 9833 6100 9924 6104
rect 9836 6096 9924 6100
rect 7496 6076 7513 6087
rect 7427 6073 7440 6076
rect 7500 6073 7513 6076
rect 7627 6075 7693 6083
rect 7767 6076 8093 6084
rect 9627 6075 9653 6083
rect 9707 6076 9733 6084
rect 9916 6086 9924 6096
rect 9927 6076 10033 6084
rect 10347 6076 10453 6084
rect 10567 6076 10753 6084
rect 10767 6076 10833 6084
rect 10927 6075 11013 6083
rect 11267 6076 11403 6084
rect 5787 6056 5973 6064
rect 7747 6056 8053 6064
rect 8347 6056 8453 6064
rect 8467 6056 8533 6064
rect 9007 6056 9113 6064
rect 6247 6036 6313 6044
rect 6647 6036 7284 6044
rect 5656 6020 5744 6024
rect 5656 6016 5747 6020
rect 5733 6007 5747 6016
rect 5847 6016 6593 6024
rect 6787 6016 6873 6024
rect 6967 6016 7153 6024
rect 7276 6024 7284 6036
rect 7307 6036 7372 6044
rect 7407 6036 7513 6044
rect 8907 6036 9093 6044
rect 9107 6036 9373 6044
rect 9667 6036 9692 6044
rect 9727 6036 9973 6044
rect 10027 6036 10153 6044
rect 10687 6036 10773 6044
rect 10787 6036 10913 6044
rect 10987 6036 11193 6044
rect 7276 6016 7633 6024
rect 7707 6016 7833 6024
rect 8747 6016 8833 6024
rect 9687 6016 10553 6024
rect 10567 6016 10953 6024
rect 10967 6016 11213 6024
rect 11227 6016 11293 6024
rect 2276 5996 2353 6004
rect 2407 5996 2573 6004
rect 2667 5996 2893 6004
rect 3347 5996 3833 6004
rect 3927 5996 4033 6004
rect 4627 5996 4773 6004
rect 5467 5996 5573 6004
rect 6307 5996 6393 6004
rect 6827 5996 6933 6004
rect 7347 5996 7833 6004
rect 8227 5996 8493 6004
rect 8707 5996 8853 6004
rect 10467 5996 10593 6004
rect 327 5976 413 5984
rect 827 5976 1333 5984
rect 1907 5976 2313 5984
rect 2827 5976 2973 5984
rect 2987 5976 3073 5984
rect 3387 5976 3413 5984
rect 3587 5976 3653 5984
rect 3727 5976 3813 5984
rect 4027 5976 4573 5984
rect 4947 5976 5453 5984
rect 5727 5976 5753 5984
rect 6567 5976 7093 5984
rect 7767 5976 8153 5984
rect 9147 5976 9433 5984
rect 9447 5976 9573 5984
rect 11007 5976 11073 5984
rect 11087 5976 11113 5984
rect 867 5956 913 5964
rect 927 5956 1093 5964
rect 1667 5956 1773 5964
rect 1787 5956 2533 5964
rect 2587 5956 3293 5964
rect 3527 5956 3653 5964
rect 4127 5956 4893 5964
rect 4947 5956 4993 5964
rect 5167 5956 5413 5964
rect 5487 5956 5913 5964
rect 6027 5956 6253 5964
rect 6427 5956 6533 5964
rect 6767 5956 7033 5964
rect 7187 5956 7353 5964
rect 7827 5956 7993 5964
rect 8007 5956 8033 5964
rect 8087 5956 8273 5964
rect 8647 5956 8773 5964
rect 8887 5956 8973 5964
rect 10747 5956 10973 5964
rect 227 5936 1433 5944
rect 2187 5936 2553 5944
rect 2867 5936 2913 5944
rect 3127 5936 3233 5944
rect 3487 5936 4733 5944
rect 5416 5944 5424 5953
rect 5416 5936 6073 5944
rect 6127 5936 6213 5944
rect 6287 5936 6653 5944
rect 7027 5936 7053 5944
rect 7267 5936 7493 5944
rect 7647 5936 9673 5944
rect 9956 5936 10084 5944
rect 2027 5916 2573 5924
rect 2616 5916 2753 5924
rect 307 5896 553 5904
rect 807 5897 873 5905
rect 967 5897 1113 5905
rect 1187 5896 1373 5904
rect 1427 5897 1453 5905
rect 1513 5904 1527 5913
rect 1513 5900 1633 5904
rect 1516 5896 1633 5900
rect 1647 5896 1833 5904
rect 2127 5896 2153 5904
rect 2616 5904 2624 5916
rect 5447 5916 6033 5924
rect 6147 5916 6213 5924
rect 7127 5916 7153 5924
rect 8747 5916 8913 5924
rect 9067 5916 9693 5924
rect 2487 5896 2624 5904
rect 2787 5896 2993 5904
rect 3067 5897 3153 5905
rect 3247 5897 3533 5905
rect 4027 5897 4053 5905
rect 4747 5897 4773 5905
rect 4787 5896 4973 5904
rect 4987 5896 5013 5904
rect 327 5875 413 5883
rect 667 5876 864 5884
rect 856 5866 864 5876
rect 1967 5876 2393 5884
rect 2907 5876 3473 5884
rect 3976 5867 3984 5894
rect 5127 5896 5353 5904
rect 5467 5896 5833 5904
rect 6067 5897 6173 5905
rect 6387 5896 6433 5904
rect 6707 5897 6773 5905
rect 6787 5896 6973 5904
rect 6987 5896 7053 5904
rect 7207 5897 7313 5905
rect 7387 5897 7553 5905
rect 7567 5896 7613 5904
rect 7807 5897 7853 5905
rect 7947 5896 7993 5904
rect 8047 5896 8084 5904
rect 4056 5867 4064 5874
rect 4427 5877 4513 5885
rect 6253 5884 6267 5893
rect 8076 5884 8084 5896
rect 8107 5897 8213 5905
rect 8687 5897 8733 5905
rect 8827 5897 8933 5905
rect 6253 5880 6584 5884
rect 6256 5876 6584 5880
rect 8076 5880 8204 5884
rect 8076 5876 8207 5880
rect -63 5856 173 5864
rect 1407 5855 1493 5863
rect 1627 5855 1733 5863
rect 2207 5855 2293 5863
rect 2707 5855 2753 5863
rect 3007 5855 3073 5863
rect 3147 5856 3233 5864
rect 3567 5856 3753 5864
rect 3967 5856 3984 5867
rect 3967 5853 3980 5856
rect 4047 5856 4064 5867
rect 4047 5853 4060 5856
rect 4136 5847 4144 5873
rect 4587 5855 4633 5863
rect 4647 5855 4673 5863
rect 4687 5856 4913 5864
rect 5227 5855 5513 5863
rect 5527 5855 5593 5863
rect 5607 5856 5773 5864
rect 5847 5856 5873 5864
rect 6247 5855 6273 5863
rect 6467 5855 6553 5863
rect 6576 5864 6584 5876
rect 8193 5867 8207 5876
rect 6576 5856 6673 5864
rect 6687 5855 6753 5863
rect 7007 5855 7073 5863
rect 7127 5855 7173 5863
rect 7267 5856 7293 5864
rect 7527 5856 7633 5864
rect 7707 5855 7733 5863
rect 8027 5855 8073 5863
rect 8316 5864 8324 5894
rect 8736 5876 9053 5884
rect 8287 5856 8324 5864
rect 8736 5864 8744 5876
rect 8956 5866 8964 5876
rect 9207 5875 9333 5883
rect 9547 5876 9713 5884
rect 9956 5886 9964 5936
rect 10076 5924 10084 5936
rect 11067 5936 11093 5944
rect 10076 5916 10113 5924
rect 10367 5916 10513 5924
rect 10667 5916 10833 5924
rect 10847 5916 10893 5924
rect 10067 5897 10173 5905
rect 10187 5897 10313 5905
rect 10380 5904 10393 5907
rect 10376 5893 10393 5904
rect 10607 5896 10653 5904
rect 8707 5856 8744 5864
rect 8767 5855 8793 5863
rect 9716 5864 9724 5874
rect 10376 5866 10384 5893
rect 10967 5897 11033 5905
rect 11127 5896 11253 5904
rect 9687 5856 9724 5864
rect 10207 5855 10333 5863
rect 10487 5855 10573 5863
rect 10867 5856 10913 5864
rect 10927 5856 10953 5864
rect 11067 5856 11273 5864
rect 267 5835 413 5843
rect 427 5835 1193 5843
rect 1327 5836 1553 5844
rect 1927 5836 2052 5844
rect 2087 5836 2333 5844
rect 2947 5836 3393 5844
rect 3627 5836 3993 5844
rect 4587 5836 5233 5844
rect 5307 5836 5373 5844
rect 6987 5836 7193 5844
rect 7787 5836 7833 5844
rect 8516 5836 8673 5844
rect 987 5816 2633 5824
rect 2707 5816 3013 5824
rect 3407 5816 3453 5824
rect 3947 5816 3993 5824
rect 4107 5816 4293 5824
rect 4316 5816 5293 5824
rect 27 5796 593 5804
rect 767 5796 1093 5804
rect 1507 5796 2973 5804
rect 4316 5804 4324 5816
rect 5567 5816 5613 5824
rect 5747 5816 5893 5824
rect 6207 5816 6413 5824
rect 6427 5816 6633 5824
rect 6647 5816 6713 5824
rect 6736 5816 7813 5824
rect 2987 5796 4324 5804
rect 4667 5796 5113 5804
rect 6736 5804 6744 5816
rect 7867 5816 8033 5824
rect 8516 5824 8524 5836
rect 9047 5835 9193 5843
rect 9207 5836 9473 5844
rect 10127 5835 10773 5843
rect 11007 5836 11313 5844
rect 8196 5816 8524 5824
rect 6067 5796 6744 5804
rect 8196 5804 8204 5816
rect 8887 5816 8993 5824
rect 9647 5816 10253 5824
rect 10527 5816 10613 5824
rect 11207 5816 11273 5824
rect 6787 5796 8204 5804
rect 10487 5796 10813 5804
rect 1007 5776 3373 5784
rect 3387 5776 5272 5784
rect 5307 5776 6493 5784
rect 6507 5776 7273 5784
rect 7627 5776 7952 5784
rect 7987 5776 8113 5784
rect 8207 5776 8273 5784
rect 8456 5776 8533 5784
rect 1667 5756 2693 5764
rect 3267 5756 3353 5764
rect 3367 5756 3793 5764
rect 4307 5756 4713 5764
rect 4727 5756 4953 5764
rect 5027 5756 6453 5764
rect 6507 5756 6573 5764
rect 7647 5756 7693 5764
rect 8247 5756 8333 5764
rect 8456 5764 8464 5776
rect 8867 5776 9793 5784
rect 8347 5756 8464 5764
rect 9827 5756 9973 5764
rect 10016 5756 10673 5764
rect 107 5736 373 5744
rect 1167 5736 1213 5744
rect 1227 5736 1733 5744
rect 2227 5736 2453 5744
rect 2567 5736 2793 5744
rect 2927 5736 3713 5744
rect 4247 5736 5033 5744
rect 5527 5736 5924 5744
rect 1367 5716 1533 5724
rect 2127 5716 2533 5724
rect 2547 5716 3933 5724
rect 4207 5716 4813 5724
rect 5916 5724 5924 5736
rect 5967 5736 6253 5744
rect 6347 5736 6573 5744
rect 6707 5736 6793 5744
rect 6807 5736 7133 5744
rect 7367 5736 7573 5744
rect 7587 5736 7813 5744
rect 7827 5736 8073 5744
rect 8087 5736 8473 5744
rect 9527 5736 9993 5744
rect 10016 5744 10024 5756
rect 10007 5736 10024 5744
rect 10787 5736 11073 5744
rect 11147 5736 11333 5744
rect 5916 5716 7193 5724
rect 7347 5716 7612 5724
rect 7647 5716 7853 5724
rect 7947 5716 8413 5724
rect 8507 5716 8733 5724
rect 9107 5716 9213 5724
rect 9327 5716 9593 5724
rect 10267 5716 10493 5724
rect 10627 5716 10653 5724
rect 11087 5716 11113 5724
rect 11167 5716 11193 5724
rect 1607 5696 1953 5704
rect 2347 5696 2433 5704
rect 2667 5696 3833 5704
rect 3967 5696 5344 5704
rect 5336 5687 5344 5696
rect 5907 5696 9953 5704
rect 10027 5696 10273 5704
rect 10287 5696 10473 5704
rect 1167 5676 2013 5684
rect 2467 5676 2633 5684
rect 2807 5676 3053 5684
rect 3067 5676 3313 5684
rect 3987 5676 4573 5684
rect 5036 5676 5293 5684
rect 5036 5667 5044 5676
rect 5347 5676 5733 5684
rect 6107 5676 6333 5684
rect 6387 5676 6433 5684
rect 6476 5676 7633 5684
rect 6476 5667 6484 5676
rect 7867 5676 8173 5684
rect 8187 5676 8353 5684
rect 9607 5676 9944 5684
rect 1247 5656 1773 5664
rect 2827 5656 3913 5664
rect 4807 5656 5033 5664
rect 5656 5656 5773 5664
rect 636 5636 1053 5644
rect 636 5627 644 5636
rect 2647 5636 4193 5644
rect 4216 5636 4593 5644
rect 287 5616 633 5624
rect 2107 5616 2173 5624
rect 2507 5616 2573 5624
rect 2667 5616 2804 5624
rect 787 5597 833 5605
rect 1547 5597 1573 5605
rect 1827 5604 1840 5607
rect 1827 5593 1844 5604
rect 2247 5597 2293 5605
rect 2447 5596 2593 5604
rect 2796 5604 2804 5616
rect 3167 5616 3713 5624
rect 4216 5624 4224 5636
rect 5187 5636 5313 5644
rect 5656 5644 5664 5656
rect 5827 5656 5973 5664
rect 6127 5656 6213 5664
rect 6367 5656 6473 5664
rect 6627 5656 7253 5664
rect 7407 5656 7533 5664
rect 7667 5656 8413 5664
rect 8567 5656 8724 5664
rect 5547 5636 5664 5644
rect 6047 5636 6073 5644
rect 6587 5636 6873 5644
rect 6887 5636 6933 5644
rect 7767 5636 7873 5644
rect 7887 5636 7993 5644
rect 8087 5636 8253 5644
rect 4027 5616 4224 5624
rect 5687 5617 5793 5625
rect 5807 5616 5853 5624
rect 6387 5616 6413 5624
rect 6807 5616 6853 5624
rect 7047 5616 7153 5624
rect 7307 5616 7433 5624
rect 7507 5616 7553 5624
rect 7627 5616 7653 5624
rect 8207 5616 8233 5624
rect 2796 5596 2813 5604
rect 3027 5597 3193 5605
rect 3907 5596 4173 5604
rect 4267 5597 4293 5605
rect 4567 5596 4893 5604
rect 407 5576 553 5584
rect 907 5556 953 5564
rect 1087 5556 1133 5564
rect 1836 5566 1844 5593
rect 1907 5576 2213 5584
rect 4336 5584 4344 5594
rect 4947 5597 5053 5605
rect 5147 5597 5213 5605
rect 5293 5604 5307 5613
rect 5293 5600 5344 5604
rect 5296 5596 5344 5600
rect 5253 5584 5267 5593
rect 5336 5586 5344 5596
rect 5947 5597 5993 5605
rect 6467 5596 6613 5604
rect 6687 5597 6733 5605
rect 7067 5597 7093 5605
rect 7456 5596 7513 5604
rect 4336 5576 4364 5584
rect 1687 5555 1773 5563
rect 1887 5556 2033 5564
rect 2087 5556 2273 5564
rect 2567 5555 2633 5563
rect 2807 5556 2893 5564
rect 3047 5556 3133 5564
rect 3407 5556 3453 5564
rect 3887 5556 4033 5564
rect 4356 5564 4364 5576
rect 4976 5580 5267 5584
rect 4976 5576 5264 5580
rect 4356 5556 4533 5564
rect 4976 5564 4984 5576
rect 5547 5576 5633 5584
rect 7456 5584 7464 5596
rect 7867 5597 7933 5605
rect 8047 5597 8153 5605
rect 8387 5597 8513 5605
rect 8600 5604 8612 5607
rect 8596 5593 8612 5604
rect 8647 5597 8673 5605
rect 8716 5604 8724 5656
rect 8827 5656 9353 5664
rect 9647 5656 9713 5664
rect 9936 5664 9944 5676
rect 10076 5676 10264 5684
rect 10076 5664 10084 5676
rect 9936 5656 10084 5664
rect 10256 5664 10264 5676
rect 10256 5656 10713 5664
rect 11096 5647 11104 5693
rect 11227 5656 11313 5664
rect 9887 5636 10093 5644
rect 11180 5644 11193 5647
rect 11176 5633 11193 5644
rect 8767 5616 8893 5624
rect 9207 5617 9253 5625
rect 9467 5616 9493 5624
rect 9927 5616 10133 5624
rect 10767 5616 10813 5624
rect 8716 5596 8744 5604
rect 8596 5584 8604 5593
rect 7287 5576 7344 5584
rect 7416 5580 7464 5584
rect 8536 5580 8604 5584
rect 4967 5556 4984 5564
rect 5007 5560 5224 5564
rect 5007 5556 5227 5560
rect 5213 5547 5227 5556
rect 5247 5555 5313 5563
rect 5667 5556 5733 5564
rect 5927 5556 6013 5564
rect 7336 5566 7344 5576
rect 7413 5576 7464 5580
rect 8533 5576 8604 5580
rect 8736 5584 8744 5596
rect 9427 5596 9653 5604
rect 10167 5596 10313 5604
rect 10367 5604 10380 5607
rect 10367 5593 10384 5604
rect 8736 5576 8764 5584
rect 7413 5567 7427 5576
rect 8533 5567 8547 5576
rect 6367 5555 6473 5563
rect 6807 5555 6893 5563
rect 7627 5555 7733 5563
rect 7947 5556 8013 5564
rect 8067 5556 8193 5564
rect 8587 5556 8613 5564
rect 8756 5564 8764 5576
rect 8807 5575 8833 5583
rect 9036 5564 9044 5574
rect 9167 5576 9233 5584
rect 10376 5586 10384 5593
rect 10856 5587 10864 5613
rect 10916 5587 10924 5613
rect 8756 5556 8784 5564
rect 9036 5556 9133 5564
rect 427 5536 653 5544
rect 667 5536 753 5544
rect 1067 5536 1153 5544
rect 2327 5536 2453 5544
rect 3287 5536 3313 5544
rect 3947 5536 4073 5544
rect 4087 5536 4113 5544
rect 4167 5536 4312 5544
rect 4347 5536 4393 5544
rect 4587 5536 4673 5544
rect 4787 5536 4933 5544
rect 6327 5536 6593 5544
rect 7767 5536 7793 5544
rect 8367 5536 8453 5544
rect 8776 5544 8784 5556
rect 9347 5556 9393 5564
rect 9507 5555 9633 5563
rect 10047 5555 10073 5563
rect 10127 5555 10153 5563
rect 10207 5555 10293 5563
rect 8776 5536 8813 5544
rect 8867 5536 8893 5544
rect 9907 5536 10113 5544
rect 1287 5516 1564 5524
rect 1127 5496 1473 5504
rect 1556 5504 1564 5516
rect 2547 5516 2613 5524
rect 3227 5516 3293 5524
rect 3956 5516 4033 5524
rect 1556 5496 1893 5504
rect 2567 5496 2613 5504
rect 3547 5496 3573 5504
rect 3956 5504 3964 5516
rect 4447 5516 4753 5524
rect 4847 5516 4993 5524
rect 5107 5516 5313 5524
rect 5827 5516 6093 5524
rect 6107 5516 6173 5524
rect 6347 5516 6533 5524
rect 6667 5516 6813 5524
rect 6967 5516 7153 5524
rect 7907 5516 8093 5524
rect 8167 5516 8193 5524
rect 8207 5516 8293 5524
rect 8407 5516 8553 5524
rect 9247 5516 9353 5524
rect 9367 5516 9433 5524
rect 9587 5516 9673 5524
rect 9727 5516 9913 5524
rect 10287 5516 10333 5524
rect 3587 5496 3964 5504
rect 5067 5496 5213 5504
rect 6867 5496 7053 5504
rect 7387 5496 7553 5504
rect 7867 5496 7913 5504
rect 8507 5496 8633 5504
rect 47 5476 173 5484
rect 827 5476 853 5484
rect 1367 5476 1533 5484
rect 2067 5476 2173 5484
rect 2287 5476 2393 5484
rect 2487 5476 2653 5484
rect 2767 5476 2853 5484
rect 2907 5476 3393 5484
rect 4007 5476 4413 5484
rect 4707 5476 4733 5484
rect 4907 5476 5813 5484
rect 5987 5476 6053 5484
rect 6547 5476 6773 5484
rect 6827 5476 7073 5484
rect 8067 5476 8113 5484
rect 8127 5476 8453 5484
rect 8467 5476 9413 5484
rect 10347 5476 10473 5484
rect 887 5456 1833 5464
rect 2227 5456 2673 5464
rect 2807 5456 3493 5464
rect 4587 5456 4633 5464
rect 5107 5456 5133 5464
rect 5147 5456 5533 5464
rect 5647 5456 5713 5464
rect 7467 5456 7653 5464
rect 7967 5456 8873 5464
rect 767 5436 1353 5444
rect 1967 5436 2233 5444
rect 2276 5436 2804 5444
rect 687 5416 1313 5424
rect 2276 5424 2284 5436
rect 1887 5416 2284 5424
rect 2367 5416 2553 5424
rect 2576 5416 2633 5424
rect 1047 5396 1093 5404
rect 1107 5396 1233 5404
rect 1447 5396 1713 5404
rect 1727 5396 1813 5404
rect 2576 5404 2584 5416
rect 2796 5424 2804 5436
rect 5227 5436 6113 5444
rect 6367 5436 6453 5444
rect 6807 5436 7692 5444
rect 7727 5436 7833 5444
rect 8407 5436 8533 5444
rect 8967 5436 9173 5444
rect 9187 5436 9513 5444
rect 10167 5436 10933 5444
rect 2796 5416 2953 5424
rect 3687 5416 4233 5424
rect 4247 5416 4313 5424
rect 4387 5416 4553 5424
rect 4567 5416 4613 5424
rect 5347 5416 5853 5424
rect 6267 5416 6973 5424
rect 8007 5416 8113 5424
rect 8267 5416 8293 5424
rect 8387 5416 8493 5424
rect 9547 5416 9853 5424
rect 10867 5416 10924 5424
rect 2307 5396 2584 5404
rect 3027 5396 3113 5404
rect 3127 5396 3233 5404
rect 4047 5396 4433 5404
rect 4476 5396 4684 5404
rect 367 5377 453 5385
rect 607 5377 673 5385
rect 1527 5377 1633 5385
rect 1847 5376 1913 5384
rect 1927 5376 2093 5384
rect 2147 5377 2193 5385
rect 2327 5376 2413 5384
rect 2467 5377 2593 5385
rect 2747 5377 2813 5385
rect 3327 5377 3353 5385
rect 3367 5376 3713 5384
rect 3767 5376 3813 5384
rect 3056 5364 3064 5374
rect 3867 5376 3973 5384
rect 4107 5377 4153 5385
rect 4476 5384 4484 5396
rect 4676 5387 4684 5396
rect 4767 5396 5193 5404
rect 7007 5396 7293 5404
rect 7307 5396 7473 5404
rect 7687 5396 7833 5404
rect 10107 5396 10333 5404
rect 10727 5396 10813 5404
rect 10916 5404 10924 5416
rect 10916 5396 10944 5404
rect 4367 5376 4484 5384
rect 4687 5376 5253 5384
rect 5267 5377 5293 5385
rect 5687 5377 5713 5385
rect 5827 5376 5973 5384
rect 6127 5376 6173 5384
rect 6367 5376 6393 5384
rect 6447 5376 6473 5384
rect 6647 5376 6773 5384
rect 6867 5376 6884 5384
rect 2987 5356 3064 5364
rect 6876 5364 6884 5376
rect 6907 5377 6933 5385
rect 7527 5376 7644 5384
rect 4547 5356 5324 5364
rect 6876 5356 6953 5364
rect 227 5336 393 5344
rect 827 5336 853 5344
rect 1027 5336 1073 5344
rect 1427 5336 1573 5344
rect 1827 5335 1893 5343
rect 2067 5335 2113 5343
rect 2167 5335 2413 5343
rect 2427 5336 2472 5344
rect 2507 5335 2573 5343
rect 2627 5335 2653 5343
rect 2847 5336 2933 5344
rect 3107 5336 3173 5344
rect 3527 5336 3633 5344
rect 3787 5335 3853 5343
rect 4187 5335 4513 5343
rect 4567 5336 4653 5344
rect 4767 5336 4853 5344
rect 5316 5346 5324 5356
rect 7636 5364 7644 5376
rect 7707 5376 7873 5384
rect 7896 5376 8053 5384
rect 7896 5364 7904 5376
rect 8267 5376 8313 5384
rect 8607 5376 8713 5384
rect 8847 5377 8913 5385
rect 9807 5376 9933 5384
rect 9947 5377 10093 5385
rect 10147 5376 10193 5384
rect 10356 5376 10393 5384
rect 7487 5356 7624 5364
rect 7636 5356 7904 5364
rect 5687 5335 5953 5343
rect 6007 5335 6033 5343
rect 6107 5335 6193 5343
rect 6487 5335 6613 5343
rect 6787 5335 6833 5343
rect 7616 5346 7624 5356
rect 9527 5356 9613 5364
rect 9887 5356 9924 5364
rect 6947 5336 7093 5344
rect 7687 5335 7713 5343
rect 7907 5335 7993 5343
rect 8867 5336 9113 5344
rect 9916 5344 9924 5356
rect 10356 5347 10364 5376
rect 10447 5376 10473 5384
rect 10487 5376 10893 5384
rect 10936 5384 10944 5396
rect 10936 5376 10964 5384
rect 10387 5357 10413 5365
rect 10847 5357 10913 5365
rect 9916 5336 10033 5344
rect 10047 5336 10073 5344
rect 10287 5336 10313 5344
rect 167 5316 633 5324
rect 647 5316 693 5324
rect 3227 5316 3253 5324
rect 3327 5316 3413 5324
rect 3767 5316 4213 5324
rect 5607 5316 6713 5324
rect 6727 5316 7124 5324
rect -63 5296 433 5304
rect 1387 5296 1513 5304
rect 2147 5296 2193 5304
rect 2267 5296 2653 5304
rect 2827 5296 2973 5304
rect 3807 5296 4013 5304
rect 4087 5296 4433 5304
rect 4647 5296 4993 5304
rect 5887 5296 5973 5304
rect 6367 5296 6493 5304
rect 6747 5296 7093 5304
rect 7116 5304 7124 5316
rect 8047 5316 8333 5324
rect 8347 5316 8473 5324
rect 8947 5316 9153 5324
rect 9547 5316 9633 5324
rect 10627 5316 10753 5324
rect 10827 5316 10913 5324
rect 7116 5296 7953 5304
rect 8047 5296 8193 5304
rect 9327 5296 9413 5304
rect 9987 5296 10113 5304
rect 10156 5296 10353 5304
rect 10156 5287 10164 5296
rect 647 5276 993 5284
rect 1327 5276 2113 5284
rect 2387 5276 2533 5284
rect 3027 5276 3153 5284
rect 3207 5276 3333 5284
rect 3787 5276 4593 5284
rect 4707 5276 4853 5284
rect 4867 5276 5044 5284
rect 1147 5256 2233 5264
rect 5036 5264 5044 5276
rect 5136 5276 5244 5284
rect 5136 5264 5144 5276
rect 5236 5267 5244 5276
rect 5567 5276 5653 5284
rect 6127 5276 6193 5284
rect 6207 5276 6753 5284
rect 6867 5276 7233 5284
rect 7587 5276 7693 5284
rect 7707 5276 7733 5284
rect 8527 5276 8613 5284
rect 8627 5276 8733 5284
rect 9267 5276 9473 5284
rect 9827 5276 9933 5284
rect 10087 5276 10153 5284
rect 10956 5284 10964 5376
rect 11076 5366 11084 5593
rect 11176 5544 11184 5633
rect 11247 5617 11273 5625
rect 11207 5576 11293 5584
rect 11176 5536 11253 5544
rect 11187 5376 11224 5384
rect 11216 5327 11224 5376
rect 11256 5327 11264 5353
rect 10867 5276 10964 5284
rect 5036 5256 5144 5264
rect 5247 5256 5373 5264
rect 5707 5256 5913 5264
rect 6187 5256 6333 5264
rect 6487 5256 6773 5264
rect 6827 5256 6873 5264
rect 7027 5256 7173 5264
rect 7307 5256 8253 5264
rect 8727 5256 8773 5264
rect 10047 5256 10213 5264
rect 10307 5256 10613 5264
rect 1547 5236 2213 5244
rect 2267 5236 2573 5244
rect 2667 5236 3073 5244
rect 3087 5236 3113 5244
rect 3287 5236 3733 5244
rect 3747 5236 4393 5244
rect 4487 5236 4693 5244
rect 4847 5236 5053 5244
rect 5336 5236 5733 5244
rect 867 5216 1033 5224
rect 1367 5216 2593 5224
rect 2727 5216 3033 5224
rect 3847 5216 4373 5224
rect 5336 5224 5344 5236
rect 5867 5236 6453 5244
rect 6467 5236 6753 5244
rect 6987 5236 7313 5244
rect 7367 5236 7613 5244
rect 7667 5236 7793 5244
rect 7807 5236 7873 5244
rect 8887 5236 9373 5244
rect 9387 5236 9653 5244
rect 9867 5236 10013 5244
rect 10787 5236 11233 5244
rect 11247 5236 11273 5244
rect 4947 5216 5344 5224
rect 5387 5216 5693 5224
rect 5767 5216 6953 5224
rect 8107 5216 8433 5224
rect 10487 5216 10533 5224
rect 10767 5216 10953 5224
rect 2227 5196 2433 5204
rect 2867 5196 3953 5204
rect 4327 5196 4813 5204
rect 6347 5196 6533 5204
rect 6587 5196 6653 5204
rect 6807 5196 6913 5204
rect 7047 5196 7233 5204
rect 7367 5196 7413 5204
rect 7547 5196 7592 5204
rect 7627 5196 8393 5204
rect 8567 5196 9033 5204
rect 10207 5196 10413 5204
rect 10627 5196 10993 5204
rect 207 5176 973 5184
rect 1047 5176 1173 5184
rect 1187 5176 1633 5184
rect 1707 5176 2153 5184
rect 2456 5176 2604 5184
rect 1427 5156 1853 5164
rect 2456 5164 2464 5176
rect 2407 5156 2464 5164
rect 2596 5164 2604 5176
rect 3307 5176 3773 5184
rect 5353 5184 5367 5193
rect 4256 5180 5367 5184
rect 4256 5176 5364 5180
rect 4256 5167 4264 5176
rect 6767 5176 6993 5184
rect 7467 5176 8893 5184
rect 9927 5176 10053 5184
rect 11187 5176 11293 5184
rect 2596 5156 3013 5164
rect 3867 5156 4253 5164
rect 4387 5156 4793 5164
rect 4887 5156 5253 5164
rect 6387 5156 6573 5164
rect 7847 5156 8373 5164
rect 707 5136 733 5144
rect 2336 5136 2573 5144
rect 467 5116 913 5124
rect 927 5116 953 5124
rect 1567 5116 1873 5124
rect 1887 5116 2093 5124
rect 2336 5124 2344 5136
rect 2627 5136 3353 5144
rect 3367 5136 4093 5144
rect 5047 5136 5133 5144
rect 5407 5136 5993 5144
rect 6407 5136 6473 5144
rect 6796 5136 6953 5144
rect 2107 5116 2344 5124
rect 2376 5116 2553 5124
rect 267 5096 333 5104
rect 1227 5096 1333 5104
rect 1347 5096 2013 5104
rect 296 5076 513 5084
rect 296 5046 304 5076
rect 567 5077 613 5085
rect 627 5076 713 5084
rect 1007 5077 1073 5085
rect 1487 5077 1593 5085
rect 1727 5077 1833 5085
rect 2307 5076 2353 5084
rect 1947 5056 2213 5064
rect 2376 5064 2384 5116
rect 2607 5116 3273 5124
rect 4407 5116 4593 5124
rect 4687 5116 4993 5124
rect 5307 5116 5613 5124
rect 5807 5116 5853 5124
rect 6487 5116 6533 5124
rect 6796 5124 6804 5136
rect 7327 5136 8653 5144
rect 10447 5136 11153 5144
rect 6647 5116 6804 5124
rect 6847 5116 6933 5124
rect 7147 5116 7293 5124
rect 7607 5116 8013 5124
rect 10267 5116 10293 5124
rect 3447 5096 3533 5104
rect 5107 5096 5193 5104
rect 6067 5096 6293 5104
rect 6456 5096 6513 5104
rect 2447 5077 2533 5085
rect 2667 5076 2733 5084
rect 2787 5076 3033 5084
rect 3127 5077 3153 5085
rect 3567 5077 3633 5085
rect 3827 5076 3884 5084
rect 2316 5056 2384 5064
rect 547 5035 813 5043
rect 987 5036 1113 5044
rect 1207 5036 1393 5044
rect 1867 5035 1893 5043
rect 2007 5036 2033 5044
rect 2087 5036 2193 5044
rect 2316 5046 2324 5056
rect 3236 5047 3244 5073
rect 2527 5036 2713 5044
rect 2767 5036 2853 5044
rect 3107 5035 3173 5043
rect 3876 5046 3884 5076
rect 4207 5077 4293 5085
rect 4487 5076 4553 5084
rect 3547 5035 3613 5043
rect 4287 5036 4333 5044
rect 4507 5035 4613 5043
rect 4716 5044 4724 5074
rect 5676 5076 5813 5084
rect 5196 5064 5204 5073
rect 4807 5056 5024 5064
rect 5196 5056 5253 5064
rect 4716 5036 4913 5044
rect 5016 5044 5024 5056
rect 5676 5064 5684 5076
rect 5867 5076 5933 5084
rect 5627 5056 5684 5064
rect 6007 5056 6064 5064
rect 5016 5036 5133 5044
rect 5947 5035 6033 5043
rect 6056 5044 6064 5056
rect 6056 5036 6073 5044
rect 6096 5044 6104 5074
rect 6327 5076 6424 5084
rect 6096 5036 6273 5044
rect 1267 5016 1613 5024
rect 2447 5016 2493 5024
rect 3227 5016 3313 5024
rect 4707 5016 4773 5024
rect 5067 5016 5173 5024
rect 5587 5016 5793 5024
rect 6416 5024 6424 5076
rect 6456 5047 6464 5096
rect 7187 5104 7200 5107
rect 7187 5096 7833 5104
rect 7187 5093 7204 5096
rect 8367 5096 8553 5104
rect 9487 5097 9713 5105
rect 10027 5096 10133 5104
rect 10607 5097 10713 5105
rect 10767 5096 10793 5104
rect 11041 5096 11403 5104
rect 6747 5076 6784 5084
rect 6776 5064 6784 5076
rect 6776 5056 6813 5064
rect 6947 5056 7113 5064
rect 7196 5066 7204 5093
rect 7507 5076 7713 5084
rect 7947 5077 8073 5085
rect 7627 5056 7753 5064
rect 6507 5036 6573 5044
rect 6667 5036 6753 5044
rect 7756 5044 7764 5053
rect 7756 5036 7833 5044
rect 7856 5044 7864 5074
rect 8207 5076 8313 5084
rect 8707 5077 8773 5085
rect 8967 5077 8993 5085
rect 9047 5076 9084 5084
rect 9076 5066 9084 5076
rect 9967 5076 10093 5084
rect 10107 5076 10433 5084
rect 11047 5076 11253 5084
rect 9187 5057 9313 5065
rect 9447 5056 9513 5064
rect 9847 5056 10253 5064
rect 10567 5056 10633 5064
rect 7856 5036 7913 5044
rect 7927 5036 8033 5044
rect 8047 5036 8133 5044
rect 8347 5036 8613 5044
rect 8987 5036 9013 5044
rect 9947 5035 10013 5043
rect 10267 5036 10533 5044
rect 10667 5036 10873 5044
rect 10967 5036 11053 5044
rect 11167 5035 11273 5043
rect 6416 5016 6473 5024
rect 6807 5016 7133 5024
rect 7147 5016 7313 5024
rect 7887 5016 7933 5024
rect 8547 5016 8673 5024
rect 8727 5016 8813 5024
rect 8967 5016 9093 5024
rect 9147 5016 9833 5024
rect 787 4996 1173 5004
rect 1767 4996 1973 5004
rect 2087 4996 2893 5004
rect 3187 4996 3293 5004
rect 3467 4996 3633 5004
rect 4127 4996 4653 5004
rect 5007 4996 5164 5004
rect 147 4976 493 4984
rect 747 4976 1273 4984
rect 2227 4976 2333 4984
rect 2567 4976 2613 4984
rect 2687 4976 2753 4984
rect 3047 4976 3393 4984
rect 3696 4976 4053 4984
rect 627 4956 773 4964
rect 1187 4956 1693 4964
rect 2287 4956 2313 4964
rect 2367 4956 2433 4964
rect 2667 4956 2833 4964
rect 3207 4956 3253 4964
rect 3696 4964 3704 4976
rect 4887 4976 4953 4984
rect 5087 4976 5133 4984
rect 5156 4984 5164 4996
rect 5267 4996 6693 5004
rect 7167 4996 7253 5004
rect 7267 4996 7644 5004
rect 5156 4976 6113 4984
rect 6167 4976 7113 4984
rect 7636 4984 7644 4996
rect 7727 4996 8313 5004
rect 8807 4996 9173 5004
rect 10107 4996 10893 5004
rect 10947 4996 11093 5004
rect 7347 4976 7604 4984
rect 7636 4976 7913 4984
rect 3407 4956 3704 4964
rect 3736 4956 3833 4964
rect 187 4936 1153 4944
rect 1167 4936 1893 4944
rect 1907 4936 2793 4944
rect 3736 4944 3744 4956
rect 4747 4956 5533 4964
rect 6167 4956 6212 4964
rect 6247 4956 6513 4964
rect 6647 4956 6713 4964
rect 7596 4964 7604 4976
rect 8427 4976 8453 4984
rect 8467 4976 8713 4984
rect 7596 4956 9893 4964
rect 11027 4956 11233 4964
rect 3487 4936 3744 4944
rect 4567 4936 4673 4944
rect 4727 4936 4853 4944
rect 5027 4936 5273 4944
rect 5547 4936 5753 4944
rect 5927 4936 6033 4944
rect 6427 4936 6893 4944
rect 7147 4936 7273 4944
rect 7327 4936 7533 4944
rect 7587 4936 7693 4944
rect 7807 4936 7912 4944
rect 7947 4936 8273 4944
rect 8667 4936 9473 4944
rect 9927 4936 10293 4944
rect 10867 4936 11053 4944
rect 1607 4916 1653 4924
rect 2147 4916 2273 4924
rect 2607 4916 2733 4924
rect 2867 4916 3753 4924
rect 3767 4916 4093 4924
rect 4627 4916 5293 4924
rect 5307 4916 5413 4924
rect 5587 4916 5673 4924
rect 6147 4916 6233 4924
rect 6447 4916 6793 4924
rect 8107 4916 8133 4924
rect 8487 4916 8573 4924
rect 9047 4916 9413 4924
rect 10067 4916 10473 4924
rect 587 4896 893 4904
rect 907 4896 1133 4904
rect 2307 4896 2373 4904
rect 2927 4896 3064 4904
rect 307 4876 1353 4884
rect 2327 4876 2364 4884
rect 647 4856 713 4864
rect 927 4856 1293 4864
rect 1427 4857 1573 4865
rect 1667 4856 1773 4864
rect 1867 4857 1933 4865
rect 2107 4856 2193 4864
rect 2267 4856 2333 4864
rect 2356 4864 2364 4876
rect 2396 4876 2553 4884
rect 2396 4864 2404 4876
rect 2567 4876 2773 4884
rect 3056 4884 3064 4896
rect 4827 4896 5192 4904
rect 5227 4896 5333 4904
rect 5987 4896 6113 4904
rect 6827 4896 7013 4904
rect 7247 4896 7413 4904
rect 7527 4896 7973 4904
rect 8167 4896 8413 4904
rect 9807 4896 10233 4904
rect 3056 4876 3313 4884
rect 3367 4876 3813 4884
rect 3827 4876 3853 4884
rect 4096 4876 4213 4884
rect 2356 4856 2404 4864
rect 2527 4856 2553 4864
rect 2847 4857 2913 4865
rect 2967 4857 3033 4865
rect 3427 4857 3513 4865
rect 3727 4857 3753 4865
rect 3276 4844 3284 4854
rect 3167 4836 3284 4844
rect 3756 4827 3764 4834
rect 4096 4844 4104 4876
rect 4547 4876 5013 4884
rect 5127 4876 5173 4884
rect 5367 4876 5593 4884
rect 5947 4876 6193 4884
rect 7167 4876 7213 4884
rect 7227 4876 8073 4884
rect 8127 4876 8533 4884
rect 9447 4876 10873 4884
rect 10887 4876 10913 4884
rect 4376 4856 4853 4864
rect 4027 4836 4104 4844
rect 4376 4846 4384 4856
rect 4967 4857 5253 4865
rect 5307 4856 5364 4864
rect 207 4815 293 4823
rect 427 4815 573 4823
rect 667 4815 793 4823
rect 887 4815 1033 4823
rect 1147 4816 1453 4824
rect 1467 4816 1593 4824
rect 1687 4815 1713 4823
rect 2127 4816 2144 4824
rect 2136 4807 2144 4816
rect 2207 4815 2313 4823
rect 2367 4815 2433 4823
rect 2587 4815 2633 4823
rect 3307 4816 3333 4824
rect 3407 4816 3433 4824
rect 3567 4816 3693 4824
rect 3747 4816 3764 4827
rect 3747 4813 3760 4816
rect 1907 4796 1953 4804
rect 2147 4796 2533 4804
rect 2847 4796 2964 4804
rect 367 4776 413 4784
rect 807 4776 1553 4784
rect 1787 4776 1973 4784
rect 2387 4776 2513 4784
rect 2587 4776 2813 4784
rect 2827 4776 2933 4784
rect 2956 4784 2964 4796
rect 3087 4796 3153 4804
rect 3387 4796 3493 4804
rect 3980 4804 3993 4807
rect 3976 4793 3993 4804
rect 4196 4804 4204 4833
rect 4607 4836 4753 4844
rect 5356 4844 5364 4856
rect 5387 4856 5573 4864
rect 6236 4856 6473 4864
rect 5356 4836 5524 4844
rect 4787 4815 4813 4823
rect 5087 4815 5213 4823
rect 5327 4815 5453 4823
rect 5516 4824 5524 4836
rect 5516 4816 5553 4824
rect 4196 4796 4533 4804
rect 5596 4804 5604 4834
rect 5847 4835 5933 4843
rect 6236 4844 6244 4856
rect 6587 4857 6653 4865
rect 6947 4857 6993 4865
rect 7287 4857 7373 4865
rect 8367 4857 8493 4865
rect 8767 4856 8933 4864
rect 8947 4856 8993 4864
rect 9827 4856 10013 4864
rect 10127 4857 10173 4865
rect 10227 4857 10273 4865
rect 10287 4856 10433 4864
rect 6167 4836 6244 4844
rect 7127 4836 7253 4844
rect 7267 4837 7473 4845
rect 8696 4827 8704 4853
rect 8896 4836 9053 4844
rect 6267 4815 6413 4823
rect 6467 4816 6573 4824
rect 6887 4815 6913 4823
rect 7027 4816 7193 4824
rect 7347 4815 7393 4823
rect 7587 4816 7713 4824
rect 8267 4816 8333 4824
rect 8507 4816 8553 4824
rect 8896 4824 8904 4836
rect 9067 4837 9453 4845
rect 8867 4816 8904 4824
rect 9487 4816 9833 4824
rect 9847 4815 9913 4823
rect 10027 4816 10193 4824
rect 10247 4816 10413 4824
rect 11087 4815 11153 4823
rect 5596 4796 5933 4804
rect 6327 4796 6533 4804
rect 7567 4796 7733 4804
rect 2956 4776 3173 4784
rect 3267 4776 3453 4784
rect 3976 4784 3984 4793
rect 7887 4795 7913 4803
rect 8907 4796 8953 4804
rect 9467 4796 9953 4804
rect 10007 4796 11013 4804
rect 3667 4776 3984 4784
rect 4027 4776 4113 4784
rect 4607 4776 4633 4784
rect 4687 4776 5373 4784
rect 8427 4776 8733 4784
rect 8787 4776 9064 4784
rect 1227 4756 1493 4764
rect 2027 4756 2113 4764
rect 3527 4756 3793 4764
rect 5047 4756 5333 4764
rect 6007 4756 6033 4764
rect 6047 4756 6393 4764
rect 7007 4756 8153 4764
rect 8267 4756 8433 4764
rect 9056 4764 9064 4776
rect 9056 4756 9393 4764
rect 9407 4756 9593 4764
rect 10947 4756 11093 4764
rect 1787 4736 1933 4744
rect 2487 4736 2513 4744
rect 2527 4736 2953 4744
rect 3067 4736 3833 4744
rect 6567 4736 6693 4744
rect 7827 4736 8073 4744
rect 9947 4736 10073 4744
rect 327 4716 593 4724
rect 1107 4716 1693 4724
rect 1747 4716 2133 4724
rect 2407 4716 2493 4724
rect 2507 4716 2633 4724
rect 2987 4716 3353 4724
rect 3407 4716 3693 4724
rect 4167 4716 4213 4724
rect 4227 4716 4713 4724
rect 5247 4716 5853 4724
rect 6527 4716 7233 4724
rect 7327 4716 7453 4724
rect 7887 4716 8493 4724
rect 9627 4716 10453 4724
rect 10467 4716 10673 4724
rect 867 4696 1673 4704
rect 2147 4696 3344 4704
rect 247 4676 833 4684
rect 1087 4676 1633 4684
rect 1647 4676 1893 4684
rect 2287 4676 2593 4684
rect 3087 4676 3273 4684
rect 3336 4684 3344 4696
rect 3487 4696 3653 4704
rect 3747 4696 3913 4704
rect 4047 4696 5813 4704
rect 5927 4696 6053 4704
rect 6487 4696 7504 4704
rect 3336 4676 3673 4684
rect 3767 4676 3933 4684
rect 5527 4676 6113 4684
rect 6187 4676 6553 4684
rect 6687 4676 7013 4684
rect 7307 4676 7473 4684
rect 7496 4684 7504 4696
rect 7907 4696 8013 4704
rect 8027 4696 8293 4704
rect 8367 4696 9193 4704
rect 9247 4696 9273 4704
rect 7496 4676 8893 4684
rect 9707 4676 10133 4684
rect 10547 4676 11273 4684
rect 1056 4656 1933 4664
rect 1056 4644 1064 4656
rect 1987 4656 2233 4664
rect 2467 4656 2553 4664
rect 2967 4656 3333 4664
rect 3347 4656 3532 4664
rect 3567 4656 3733 4664
rect 3747 4656 3993 4664
rect 4667 4656 5053 4664
rect 5067 4656 5353 4664
rect 5587 4656 6313 4664
rect 7447 4656 7593 4664
rect 8987 4656 9133 4664
rect 9527 4656 10233 4664
rect 287 4636 1064 4644
rect 1707 4636 2493 4644
rect 2556 4644 2564 4653
rect 2556 4636 5133 4644
rect 5147 4636 6373 4644
rect 6387 4636 6713 4644
rect 6727 4636 6793 4644
rect 6807 4636 7133 4644
rect 7147 4636 7293 4644
rect 8847 4636 10013 4644
rect 10167 4636 10213 4644
rect 10307 4636 10993 4644
rect 1467 4616 1533 4624
rect 2047 4616 2393 4624
rect 2627 4616 3553 4624
rect 3627 4616 3953 4624
rect 5387 4616 5553 4624
rect 5567 4616 6013 4624
rect 6127 4616 6393 4624
rect 6407 4616 6544 4624
rect 427 4596 853 4604
rect 1587 4596 1693 4604
rect 1887 4596 1993 4604
rect 2107 4596 3573 4604
rect 3667 4596 4273 4604
rect 4287 4596 4433 4604
rect 4507 4596 4833 4604
rect 4847 4596 4953 4604
rect 5127 4596 5953 4604
rect 5976 4596 6333 4604
rect 207 4576 373 4584
rect 1307 4576 1433 4584
rect 1447 4576 1533 4584
rect 1547 4576 1753 4584
rect 1767 4576 1813 4584
rect 2207 4576 2253 4584
rect 2307 4576 2333 4584
rect 2507 4576 2973 4584
rect 3027 4576 3233 4584
rect 3247 4576 3373 4584
rect 3827 4576 4033 4584
rect 5307 4576 5433 4584
rect 5447 4576 5573 4584
rect 5976 4584 5984 4596
rect 6387 4596 6413 4604
rect 6427 4596 6513 4604
rect 6536 4604 6544 4616
rect 6567 4616 6733 4624
rect 7827 4616 8173 4624
rect 8227 4616 8804 4624
rect 6536 4596 6953 4604
rect 7287 4596 7413 4604
rect 7987 4596 8093 4604
rect 8796 4604 8804 4616
rect 10247 4616 10273 4624
rect 8796 4596 8993 4604
rect 9467 4596 9833 4604
rect 11167 4596 11193 4604
rect 5727 4576 5984 4584
rect 6056 4576 8113 4584
rect 547 4557 613 4565
rect 707 4556 733 4564
rect 827 4557 853 4565
rect 1347 4557 1373 4565
rect 1387 4556 1573 4564
rect 2287 4557 2433 4565
rect 2647 4557 2733 4565
rect 3167 4557 3213 4565
rect 847 4536 953 4544
rect 147 4515 173 4523
rect 447 4516 533 4524
rect 647 4515 733 4523
rect 1116 4507 1124 4554
rect 2056 4544 2064 4554
rect 3227 4557 3253 4565
rect 3607 4557 3653 4565
rect 4067 4557 4133 4565
rect 4667 4556 4884 4564
rect 2056 4536 2664 4544
rect 1247 4516 1464 4524
rect 767 4496 873 4504
rect 1307 4496 1373 4504
rect 1456 4504 1464 4516
rect 1487 4516 1553 4524
rect 1887 4516 1993 4524
rect 2227 4515 2253 4523
rect 2327 4516 2633 4524
rect 2656 4524 2664 4536
rect 2827 4536 2964 4544
rect 2956 4526 2964 4536
rect 3287 4536 3473 4544
rect 4056 4536 4193 4544
rect 2656 4516 2693 4524
rect 3587 4520 3624 4524
rect 3587 4516 3627 4520
rect 3613 4507 3627 4516
rect 3687 4515 3773 4523
rect 3967 4515 3993 4523
rect 4056 4524 4064 4536
rect 4236 4544 4244 4554
rect 4207 4536 4244 4544
rect 4876 4544 4884 4556
rect 4947 4556 5113 4564
rect 5607 4557 5633 4565
rect 5747 4557 5773 4565
rect 6056 4564 6064 4576
rect 8127 4576 8233 4584
rect 8247 4576 8333 4584
rect 8376 4576 8453 4584
rect 5967 4556 6064 4564
rect 6087 4556 6473 4564
rect 6616 4556 7033 4564
rect 4876 4536 4904 4544
rect 4007 4516 4064 4524
rect 4147 4516 4253 4524
rect 4727 4516 4853 4524
rect 4896 4524 4904 4536
rect 6616 4544 6624 4556
rect 7127 4557 7153 4565
rect 7207 4557 7233 4565
rect 7887 4556 8013 4564
rect 6007 4536 6624 4544
rect 6647 4536 6893 4544
rect 4896 4516 4913 4524
rect 5327 4516 5453 4524
rect 5507 4516 5573 4524
rect 5727 4516 5793 4524
rect 6307 4515 6373 4523
rect 6987 4516 7093 4524
rect 7187 4516 7273 4524
rect 7376 4524 7384 4554
rect 8356 4527 8364 4553
rect 8376 4546 8384 4576
rect 10607 4577 10653 4585
rect 10667 4576 10713 4584
rect 9247 4557 9293 4565
rect 9667 4557 9773 4565
rect 9867 4557 9893 4565
rect 9987 4556 10213 4564
rect 10316 4556 10873 4564
rect 8387 4536 8453 4544
rect 7376 4516 7433 4524
rect 8027 4515 8053 4523
rect 1456 4496 1593 4504
rect 1607 4496 1793 4504
rect 3167 4496 3193 4504
rect 5947 4496 6073 4504
rect 6087 4496 6253 4504
rect 6747 4496 6853 4504
rect 7347 4496 7793 4504
rect 967 4476 1093 4484
rect 1107 4476 1313 4484
rect 1336 4476 1753 4484
rect 547 4456 673 4464
rect 1336 4464 1344 4476
rect 1867 4476 2033 4484
rect 2047 4476 2133 4484
rect 2307 4476 2333 4484
rect 2487 4476 2553 4484
rect 2647 4476 3113 4484
rect 3367 4476 3513 4484
rect 3527 4476 3593 4484
rect 3647 4476 3793 4484
rect 3947 4476 4013 4484
rect 4207 4476 4893 4484
rect 6947 4476 7673 4484
rect 7727 4476 7853 4484
rect 8007 4476 8053 4484
rect 8267 4476 8313 4484
rect 907 4456 1344 4464
rect 1707 4456 2153 4464
rect 3347 4456 3413 4464
rect 3867 4456 4933 4464
rect 5107 4456 6524 4464
rect 4347 4436 5233 4444
rect 5296 4436 6333 4444
rect 5296 4427 5304 4436
rect 6516 4444 6524 4456
rect 7127 4456 7213 4464
rect 7227 4456 7353 4464
rect 7407 4456 7553 4464
rect 8616 4464 8624 4534
rect 8747 4536 8933 4544
rect 10316 4546 10324 4556
rect 10887 4556 10953 4564
rect 11127 4556 11193 4564
rect 10367 4537 10493 4545
rect 10627 4536 11053 4544
rect 10653 4527 10667 4536
rect 9147 4515 9173 4523
rect 9227 4516 9273 4524
rect 9487 4516 9613 4524
rect 9627 4516 9673 4524
rect 9787 4516 9953 4524
rect 9967 4516 10113 4524
rect 8727 4496 8773 4504
rect 8907 4496 9044 4504
rect 9036 4484 9044 4496
rect 10267 4496 11213 4504
rect 9036 4476 9433 4484
rect 8447 4456 8544 4464
rect 8616 4456 8713 4464
rect 8536 4447 8544 4456
rect 10027 4456 10273 4464
rect 10287 4456 10853 4464
rect 6516 4436 8513 4444
rect 8536 4436 8553 4447
rect 8540 4433 8553 4436
rect 9027 4436 9233 4444
rect 9567 4436 9853 4444
rect 227 4416 393 4424
rect 2547 4416 2893 4424
rect 3367 4416 3493 4424
rect 3907 4416 5293 4424
rect 5367 4416 5633 4424
rect 5647 4416 6173 4424
rect 6547 4416 8273 4424
rect 8547 4416 8833 4424
rect 9707 4416 9793 4424
rect 10487 4416 10593 4424
rect 10687 4416 10753 4424
rect 2087 4396 2353 4404
rect 2727 4396 3073 4404
rect 3187 4396 3553 4404
rect 3687 4396 3753 4404
rect 3927 4396 4233 4404
rect 4447 4396 4873 4404
rect 4887 4396 4973 4404
rect 5527 4396 5593 4404
rect 5847 4396 5973 4404
rect 6327 4396 6353 4404
rect 6527 4396 6593 4404
rect 6607 4396 7333 4404
rect 7527 4396 7613 4404
rect 7967 4396 8264 4404
rect 8256 4387 8264 4396
rect 8527 4396 8933 4404
rect 8947 4396 9093 4404
rect 9607 4396 9673 4404
rect 9807 4396 9893 4404
rect 9907 4396 10073 4404
rect 10207 4396 10313 4404
rect 227 4376 673 4384
rect 847 4376 913 4384
rect 2767 4376 2933 4384
rect 5467 4376 5733 4384
rect 6567 4376 6593 4384
rect 6607 4376 6873 4384
rect 7207 4376 7493 4384
rect 7547 4376 7833 4384
rect 8267 4376 8433 4384
rect 8567 4376 8853 4384
rect 9127 4376 9413 4384
rect 9487 4376 9593 4384
rect 10127 4376 10573 4384
rect 920 4364 933 4367
rect 916 4353 933 4364
rect 1227 4356 1353 4364
rect 2607 4356 2673 4364
rect 3707 4356 3733 4364
rect 3747 4356 3813 4364
rect 4847 4356 4913 4364
rect 5327 4356 5353 4364
rect 6047 4356 6493 4364
rect 6907 4356 7093 4364
rect 7187 4356 8193 4364
rect 8287 4356 8533 4364
rect 9747 4356 9813 4364
rect 687 4337 733 4345
rect 916 4344 924 4353
rect 896 4336 924 4344
rect 376 4307 384 4333
rect 436 4324 444 4334
rect 436 4316 513 4324
rect 707 4296 833 4304
rect 896 4306 904 4336
rect 1167 4337 1193 4345
rect 1287 4336 1393 4344
rect 1407 4337 1513 4345
rect 1707 4337 1833 4345
rect 2027 4337 2073 4345
rect 1876 4316 1993 4324
rect 947 4296 1133 4304
rect 1387 4295 1433 4303
rect 1447 4296 1493 4304
rect 1876 4306 1884 4316
rect 2096 4306 2104 4353
rect 2267 4337 2373 4345
rect 2387 4337 2533 4345
rect 2587 4336 2753 4344
rect 2807 4336 2913 4344
rect 2927 4336 2993 4344
rect 3047 4337 3073 4345
rect 3227 4337 3373 4345
rect 3507 4336 3673 4344
rect 3456 4324 3464 4334
rect 3907 4337 3953 4345
rect 4007 4337 4113 4345
rect 4127 4337 4153 4345
rect 4207 4336 4373 4344
rect 4427 4337 4453 4345
rect 4567 4337 4633 4345
rect 4807 4336 4833 4344
rect 5167 4337 5513 4345
rect 5567 4336 5653 4344
rect 5727 4337 5813 4345
rect 6027 4337 6532 4345
rect 6567 4337 6633 4345
rect 6647 4336 6753 4344
rect 7147 4336 7384 4344
rect 3456 4316 3484 4324
rect 2387 4296 2413 4304
rect 2527 4296 2713 4304
rect 3027 4295 3053 4303
rect 3476 4304 3484 4316
rect 3787 4316 4184 4324
rect 4176 4306 4184 4316
rect 5296 4316 5373 4324
rect 3476 4296 3693 4304
rect 3476 4287 3484 4296
rect 4447 4296 4473 4304
rect 4587 4295 4613 4303
rect 4667 4296 4853 4304
rect 5027 4295 5113 4303
rect 5296 4304 5304 4316
rect 5387 4316 5453 4324
rect 7376 4324 7384 4336
rect 7407 4336 7593 4344
rect 7647 4337 7693 4345
rect 8027 4337 8133 4345
rect 8647 4337 8673 4345
rect 8987 4337 9153 4345
rect 9387 4337 9473 4345
rect 9860 4344 9873 4347
rect 9856 4333 9873 4344
rect 9947 4336 10313 4344
rect 10467 4336 10533 4344
rect 5867 4316 6664 4324
rect 7376 4316 7624 4324
rect 5127 4296 5304 4304
rect 5327 4296 5353 4304
rect 5367 4296 5493 4304
rect 5547 4295 5593 4303
rect 5667 4295 5733 4303
rect 5827 4296 6153 4304
rect 6656 4306 6664 4316
rect 6347 4295 6613 4303
rect 6667 4296 6733 4304
rect 7047 4296 7352 4304
rect 7387 4296 7433 4304
rect 7616 4306 7624 4316
rect 7547 4295 7573 4303
rect 7707 4296 7813 4304
rect 7867 4296 7933 4304
rect 8507 4296 8633 4304
rect 8747 4296 8773 4304
rect 8827 4296 9133 4304
rect 9407 4296 9513 4304
rect 9856 4306 9864 4333
rect 10576 4324 10584 4334
rect 11027 4336 11233 4344
rect 10576 4316 11084 4324
rect 9627 4296 9813 4304
rect 9927 4296 10033 4304
rect 10527 4295 10973 4303
rect 11076 4304 11084 4316
rect 11076 4296 11213 4304
rect 1647 4276 1693 4284
rect 2447 4276 2613 4284
rect 2927 4276 2973 4284
rect 3167 4276 3253 4284
rect 3467 4276 3484 4287
rect 3467 4273 3480 4276
rect 3747 4276 3853 4284
rect 3947 4276 4553 4284
rect 4767 4276 5453 4284
rect 6987 4276 7073 4284
rect 7087 4276 7393 4284
rect 7467 4276 8113 4284
rect 10187 4276 11053 4284
rect 227 4256 413 4264
rect 527 4256 633 4264
rect 647 4256 833 4264
rect 1347 4256 1393 4264
rect 1787 4256 2013 4264
rect 2947 4256 3033 4264
rect 3647 4256 3973 4264
rect 4547 4256 4973 4264
rect 5067 4256 5253 4264
rect 5427 4256 5753 4264
rect 6227 4256 6633 4264
rect 7067 4256 7373 4264
rect 8427 4256 9033 4264
rect 9647 4256 9744 4264
rect 167 4236 193 4244
rect 467 4236 933 4244
rect 1327 4236 1453 4244
rect 1687 4236 2253 4244
rect 2887 4236 3293 4244
rect 3827 4236 4433 4244
rect 5107 4236 5153 4244
rect 5807 4236 6133 4244
rect 6627 4236 6993 4244
rect 7447 4236 7893 4244
rect 8207 4236 8893 4244
rect 9347 4236 9573 4244
rect 9736 4244 9744 4256
rect 9827 4256 10033 4264
rect 10047 4256 10093 4264
rect 10107 4256 10133 4264
rect 10307 4256 10553 4264
rect 10567 4256 11073 4264
rect 9736 4236 10113 4244
rect 10467 4236 10773 4244
rect 947 4216 1053 4224
rect 2247 4216 2853 4224
rect 2907 4216 3053 4224
rect 3067 4216 3473 4224
rect 3696 4216 3773 4224
rect 427 4196 813 4204
rect 1587 4196 1713 4204
rect 1727 4196 2053 4204
rect 2387 4196 3172 4204
rect 3696 4204 3704 4216
rect 3967 4216 3993 4224
rect 4727 4216 4853 4224
rect 5187 4216 5313 4224
rect 6007 4216 6353 4224
rect 6367 4216 6413 4224
rect 6647 4216 7193 4224
rect 7307 4216 7853 4224
rect 8127 4216 8293 4224
rect 8347 4216 8633 4224
rect 8707 4216 8793 4224
rect 8807 4216 8913 4224
rect 9427 4216 9633 4224
rect 9727 4216 10173 4224
rect 3207 4196 3704 4204
rect 3847 4196 4333 4204
rect 4587 4196 5424 4204
rect 1447 4176 1613 4184
rect 2267 4176 3713 4184
rect 3867 4176 4413 4184
rect 4687 4176 4873 4184
rect 5416 4184 5424 4196
rect 5447 4196 5573 4204
rect 5927 4196 6093 4204
rect 6767 4196 7153 4204
rect 8607 4196 8953 4204
rect 9987 4196 10333 4204
rect 10487 4196 10533 4204
rect 10547 4196 10613 4204
rect 10987 4196 11333 4204
rect 5416 4176 5553 4184
rect 5847 4176 6613 4184
rect 6667 4176 7993 4184
rect 8007 4176 8033 4184
rect 8047 4176 8253 4184
rect 8267 4176 8973 4184
rect 10107 4176 10233 4184
rect 1147 4156 1573 4164
rect 2127 4156 4513 4164
rect 4527 4156 5053 4164
rect 5207 4156 5593 4164
rect 6427 4156 6493 4164
rect 6727 4156 6853 4164
rect 6967 4156 7273 4164
rect 7847 4156 7973 4164
rect 8447 4156 8653 4164
rect 1207 4136 2133 4144
rect 2327 4136 2493 4144
rect 2507 4136 3173 4144
rect 3187 4136 3273 4144
rect 3287 4136 3433 4144
rect 3487 4136 3733 4144
rect 4047 4136 4113 4144
rect 4627 4136 4693 4144
rect 4947 4136 5073 4144
rect 5307 4136 6613 4144
rect 7076 4136 7173 4144
rect 747 4116 2773 4124
rect 2787 4116 3092 4124
rect 3127 4116 5953 4124
rect 7076 4124 7084 4136
rect 7367 4136 7953 4144
rect 8147 4136 10573 4144
rect 10587 4136 11113 4144
rect 6027 4116 7084 4124
rect 7127 4116 7153 4124
rect 7627 4116 7813 4124
rect 8347 4116 8493 4124
rect 10247 4116 10373 4124
rect 787 4096 1373 4104
rect 1427 4096 1513 4104
rect 1527 4096 1833 4104
rect 1907 4096 2353 4104
rect 2367 4096 2533 4104
rect 3287 4096 3413 4104
rect 3567 4096 4133 4104
rect 4207 4096 4233 4104
rect 4247 4096 4553 4104
rect 4607 4096 5493 4104
rect 5567 4096 5853 4104
rect 5907 4096 6693 4104
rect 6787 4096 6933 4104
rect 7007 4096 8373 4104
rect 8727 4096 9553 4104
rect 10547 4096 10693 4104
rect 10707 4096 10993 4104
rect 607 4076 1213 4084
rect 1987 4076 2333 4084
rect 2347 4076 2413 4084
rect 3087 4076 3453 4084
rect 3527 4076 3993 4084
rect 4107 4076 5253 4084
rect 5267 4076 5873 4084
rect 6047 4076 6213 4084
rect 7047 4076 7173 4084
rect 7567 4076 7853 4084
rect 7967 4076 8593 4084
rect 9287 4076 9393 4084
rect 11167 4076 11253 4084
rect 1367 4056 1473 4064
rect 1687 4056 1893 4064
rect 2167 4056 2333 4064
rect 2767 4056 3013 4064
rect 3087 4056 3473 4064
rect 3607 4056 3673 4064
rect 4036 4056 4473 4064
rect 567 4037 633 4045
rect 1007 4037 1033 4045
rect 1227 4036 1292 4044
rect 1527 4037 1573 4045
rect 376 4007 384 4033
rect 707 4016 864 4024
rect 667 3995 733 4003
rect 856 4004 864 4016
rect 1316 4007 1324 4034
rect 2147 4016 2433 4024
rect 856 3996 1053 4004
rect 1107 3995 1133 4003
rect 1307 3996 1324 4007
rect 1307 3993 1320 3996
rect 1347 3995 1432 4003
rect 1467 3995 1593 4003
rect 1887 3995 1993 4003
rect 2107 3996 2453 4004
rect 2476 4004 2484 4033
rect 2687 4037 2693 4045
rect 2707 4037 2713 4045
rect 2987 4036 3033 4044
rect 3216 4024 3224 4034
rect 3787 4036 3853 4044
rect 4036 4044 4044 4056
rect 7647 4056 7673 4064
rect 7687 4056 8033 4064
rect 8047 4056 8113 4064
rect 8247 4056 8513 4064
rect 8527 4056 8613 4064
rect 9627 4057 10533 4065
rect 10647 4056 10673 4064
rect 10696 4056 11033 4064
rect 3867 4036 4044 4044
rect 4067 4036 4253 4044
rect 4267 4036 4352 4044
rect 4387 4036 4493 4044
rect 4747 4037 4793 4045
rect 4887 4037 4933 4045
rect 5027 4037 5113 4045
rect 5167 4037 5213 4045
rect 3693 4024 3707 4033
rect 2887 4016 3224 4024
rect 3396 4020 3707 4024
rect 3396 4016 3704 4020
rect 2476 3996 2513 4004
rect 2947 3995 2993 4003
rect 3396 4004 3404 4016
rect 4007 4016 4653 4024
rect 4696 4024 4704 4034
rect 5347 4036 5453 4044
rect 5867 4036 5893 4044
rect 6127 4036 6152 4044
rect 6987 4037 7053 4045
rect 7527 4037 7593 4045
rect 4667 4016 4704 4024
rect 3047 3996 3404 4004
rect 3427 3996 3553 4004
rect 3667 3996 3733 4004
rect 3887 3995 3913 4003
rect 4007 3995 4073 4003
rect 4287 3995 4373 4003
rect 4427 3996 4513 4004
rect 4527 3995 4573 4003
rect 4767 3995 4893 4003
rect 4936 4000 4953 4004
rect 4933 3996 4953 4000
rect 4933 3987 4947 3996
rect 5127 3996 5233 4004
rect 5247 3996 5293 4004
rect 5767 3996 5933 4004
rect 6176 4004 6184 4033
rect 6176 3996 6193 4004
rect 6367 3995 6393 4003
rect 6656 4004 6664 4033
rect 7316 4016 7613 4024
rect 6647 3996 6664 4004
rect 6847 3996 6913 4004
rect 6967 3995 7073 4003
rect 7127 3996 7213 4004
rect 7316 4006 7324 4016
rect 7776 4024 7784 4034
rect 8407 4037 8473 4045
rect 7707 4016 7784 4024
rect 7387 3996 7533 4004
rect 7816 4004 7824 4033
rect 8736 4024 8744 4053
rect 8767 4037 8813 4045
rect 8867 4037 8933 4045
rect 8987 4036 9133 4044
rect 9187 4037 9253 4045
rect 9447 4036 9713 4044
rect 9847 4036 9993 4044
rect 8696 4016 8744 4024
rect 7807 3996 7824 4004
rect 7987 3996 8073 4004
rect 8247 3996 8313 4004
rect 8696 4006 8704 4016
rect 10387 4017 10473 4025
rect 10696 4024 10704 4056
rect 11067 4036 11173 4044
rect 10676 4016 10704 4024
rect 8747 3995 8793 4003
rect 8967 3996 9273 4004
rect 9347 3996 9373 4004
rect 9867 3995 9893 4003
rect 9907 3996 10133 4004
rect 10247 3996 10493 4004
rect 10676 4004 10684 4016
rect 10607 3996 10684 4004
rect 347 3976 433 3984
rect 2687 3976 2793 3984
rect 2927 3976 2973 3984
rect 3167 3976 3213 3984
rect 3327 3976 3393 3984
rect 3647 3976 3813 3984
rect 3827 3976 3853 3984
rect 4707 3976 4793 3984
rect 5487 3976 5713 3984
rect 7567 3976 7593 3984
rect 8336 3976 8453 3984
rect 627 3956 853 3964
rect 2107 3956 2233 3964
rect 2467 3956 2553 3964
rect 3207 3956 3953 3964
rect 4427 3956 4913 3964
rect 4967 3956 5433 3964
rect 6147 3956 6753 3964
rect 6887 3956 6913 3964
rect 7047 3956 8013 3964
rect 8336 3964 8344 3976
rect 8887 3976 9633 3984
rect 10007 3976 10053 3984
rect 10836 3984 10844 4014
rect 10967 4016 11233 4024
rect 11047 3996 11193 4004
rect 10836 3976 10953 3984
rect 8167 3956 8344 3964
rect 9207 3956 9593 3964
rect 11027 3956 11093 3964
rect 227 3936 593 3944
rect 647 3936 693 3944
rect 1647 3936 1913 3944
rect 1967 3936 2393 3944
rect 2447 3936 3073 3944
rect 3227 3936 3433 3944
rect 3627 3936 4013 3944
rect 4147 3936 4593 3944
rect 4727 3936 4813 3944
rect 4976 3936 5033 3944
rect 1067 3916 1213 3924
rect 1227 3916 3213 3924
rect 3227 3916 3533 3924
rect 3767 3916 4313 3924
rect 4367 3916 4473 3924
rect 4747 3916 4833 3924
rect 4976 3924 4984 3936
rect 5047 3936 5193 3944
rect 6447 3936 6653 3944
rect 6707 3936 6904 3944
rect 4927 3916 4984 3924
rect 5227 3916 6104 3924
rect 407 3896 513 3904
rect 1087 3896 1133 3904
rect 1147 3896 1373 3904
rect 2007 3896 2273 3904
rect 2507 3896 2953 3904
rect 3007 3896 3153 3904
rect 3247 3896 3453 3904
rect 3807 3896 3933 3904
rect 4047 3896 4413 3904
rect 4507 3896 4984 3904
rect 627 3876 713 3884
rect 1287 3876 1393 3884
rect 1407 3876 2313 3884
rect 2327 3876 3373 3884
rect 3387 3876 3953 3884
rect 4027 3876 4473 3884
rect 4976 3884 4984 3896
rect 5007 3896 5153 3904
rect 5627 3896 5793 3904
rect 5867 3896 5893 3904
rect 5907 3896 6073 3904
rect 6096 3904 6104 3916
rect 6127 3916 6273 3924
rect 6896 3924 6904 3936
rect 7096 3936 8344 3944
rect 7096 3924 7104 3936
rect 6896 3916 7104 3924
rect 7287 3916 7353 3924
rect 7576 3916 7613 3924
rect 6096 3896 6773 3904
rect 7576 3904 7584 3916
rect 7767 3916 8313 3924
rect 8336 3924 8344 3936
rect 8367 3936 8453 3944
rect 10296 3940 10513 3944
rect 10293 3936 10513 3940
rect 10293 3927 10307 3936
rect 8336 3916 8853 3924
rect 8867 3916 9153 3924
rect 9787 3916 10013 3924
rect 10027 3916 10173 3924
rect 11007 3916 11073 3924
rect 6827 3896 7084 3904
rect 4976 3876 5213 3884
rect 5267 3876 6793 3884
rect 7076 3884 7084 3896
rect 7376 3896 7584 3904
rect 7076 3876 7133 3884
rect 7376 3884 7384 3896
rect 7607 3896 8513 3904
rect 8647 3896 8973 3904
rect 10527 3896 10573 3904
rect 7347 3876 7384 3884
rect 7456 3876 8333 3884
rect 1327 3856 2493 3864
rect 2547 3856 3113 3864
rect 3407 3856 3453 3864
rect 3467 3856 3893 3864
rect 4787 3856 5024 3864
rect 487 3836 593 3844
rect 607 3836 653 3844
rect 747 3836 1853 3844
rect 2147 3836 2204 3844
rect 247 3817 553 3825
rect 707 3816 853 3824
rect 907 3817 993 3825
rect 1347 3817 1413 3825
rect 1627 3816 1693 3824
rect 1707 3816 1833 3824
rect 1847 3816 2013 3824
rect 2196 3824 2204 3836
rect 2436 3836 2513 3844
rect 2436 3824 2444 3836
rect 2747 3836 3284 3844
rect 3276 3828 3284 3836
rect 3867 3836 4053 3844
rect 5016 3844 5024 3856
rect 5527 3856 5673 3864
rect 5987 3856 6353 3864
rect 6627 3856 6773 3864
rect 6847 3856 7253 3864
rect 7456 3864 7464 3876
rect 8387 3876 8624 3884
rect 7267 3856 7464 3864
rect 7487 3856 7653 3864
rect 7827 3856 8293 3864
rect 8407 3856 8533 3864
rect 8616 3864 8624 3876
rect 8667 3876 9173 3884
rect 9187 3876 9413 3884
rect 9427 3876 9893 3884
rect 10067 3876 10813 3884
rect 8616 3856 8644 3864
rect 5016 3836 5693 3844
rect 8636 3844 8644 3856
rect 8827 3856 8933 3864
rect 9427 3856 9473 3864
rect 10967 3856 11093 3864
rect 8636 3836 8664 3844
rect 2196 3816 2444 3824
rect 2487 3816 2533 3824
rect 2707 3816 2724 3824
rect 1356 3796 1493 3804
rect 87 3775 213 3783
rect 227 3776 273 3784
rect 627 3775 673 3783
rect 727 3775 773 3783
rect 787 3775 1073 3783
rect 1167 3776 1213 3784
rect 1356 3786 1364 3796
rect 1507 3796 1713 3804
rect 1727 3796 2173 3804
rect 2427 3796 2633 3804
rect 2716 3804 2724 3816
rect 2927 3816 3033 3824
rect 3287 3817 3333 3825
rect 2716 3796 2813 3804
rect 3247 3804 3260 3807
rect 3247 3793 3264 3804
rect 1807 3776 2133 3784
rect 3256 3784 3264 3793
rect 3256 3776 3313 3784
rect 3356 3786 3364 3833
rect 3387 3816 3493 3824
rect 3667 3817 3733 3825
rect 4027 3816 4113 3824
rect 4287 3817 4353 3825
rect 4547 3817 4713 3825
rect 4927 3816 4993 3824
rect 5127 3816 5313 3824
rect 5407 3817 5473 3825
rect 5747 3817 5793 3825
rect 5947 3817 6033 3825
rect 6107 3817 6133 3825
rect 6187 3816 6233 3824
rect 5053 3804 5067 3813
rect 5016 3800 5067 3804
rect 5016 3796 5064 3800
rect 3407 3775 3453 3783
rect 3567 3775 3593 3783
rect 3647 3775 3673 3783
rect 3747 3776 3833 3784
rect 4127 3776 4193 3784
rect 4367 3776 4493 3784
rect 4667 3776 4953 3784
rect 5016 3786 5024 3796
rect 6176 3804 6184 3814
rect 6407 3816 6464 3824
rect 6087 3796 6184 3804
rect 6456 3804 6464 3816
rect 6487 3817 6653 3825
rect 7007 3817 7033 3825
rect 7087 3817 7113 3825
rect 7127 3816 7393 3824
rect 7407 3816 7473 3824
rect 7527 3817 7573 3825
rect 7627 3816 7693 3824
rect 8167 3816 8213 3824
rect 8267 3816 8373 3824
rect 8487 3816 8613 3824
rect 8656 3824 8664 3836
rect 10487 3836 10853 3844
rect 8656 3816 9113 3824
rect 9127 3816 9273 3824
rect 9347 3817 9373 3825
rect 9387 3816 9633 3824
rect 9827 3816 9933 3824
rect 10496 3816 10653 3824
rect 6456 3796 6504 3804
rect 5207 3776 5233 3784
rect 5247 3775 5333 3783
rect 5516 3776 5713 3784
rect 827 3756 913 3764
rect 1487 3756 2213 3764
rect 2287 3756 2313 3764
rect 2667 3756 2733 3764
rect 3067 3756 3193 3764
rect 3247 3756 3513 3764
rect 3987 3756 4253 3764
rect 5516 3764 5524 3776
rect 5727 3776 5833 3784
rect 6256 3776 6373 3784
rect 5487 3756 5524 3764
rect 6256 3764 6264 3776
rect 6427 3776 6473 3784
rect 6496 3784 6504 3796
rect 7147 3796 7333 3804
rect 7767 3797 7793 3805
rect 7847 3796 8013 3804
rect 10027 3796 10473 3804
rect 6496 3776 6593 3784
rect 6867 3776 7113 3784
rect 7507 3776 7553 3784
rect 8016 3776 8253 3784
rect 8016 3767 8024 3776
rect 8367 3776 8453 3784
rect 8547 3775 8653 3783
rect 8827 3775 9133 3783
rect 9147 3776 9333 3784
rect 9687 3776 9873 3784
rect 9956 3784 9964 3794
rect 10496 3804 10504 3816
rect 10487 3796 10504 3804
rect 9927 3776 9964 3784
rect 10527 3775 10553 3783
rect 10887 3775 10953 3783
rect 6167 3756 6264 3764
rect 7007 3756 7233 3764
rect 8007 3756 8024 3767
rect 8007 3753 8020 3756
rect 9287 3756 9393 3764
rect 9407 3756 9613 3764
rect 10807 3756 11153 3764
rect 816 3744 824 3753
rect 587 3736 824 3744
rect 1376 3736 1453 3744
rect 187 3716 413 3724
rect 427 3716 753 3724
rect 1376 3724 1384 3736
rect 1527 3736 1813 3744
rect 2327 3736 2453 3744
rect 2467 3736 2613 3744
rect 2847 3736 2893 3744
rect 3267 3736 3453 3744
rect 3507 3736 4133 3744
rect 4307 3736 4753 3744
rect 4867 3736 4993 3744
rect 5567 3736 5753 3744
rect 6287 3736 6633 3744
rect 6807 3736 7593 3744
rect 8167 3736 8393 3744
rect 8527 3736 8813 3744
rect 8947 3736 9133 3744
rect 9987 3736 10053 3744
rect 10507 3736 10593 3744
rect 10647 3736 10833 3744
rect 10927 3736 10953 3744
rect 887 3716 1384 3724
rect 2067 3716 2633 3724
rect 3013 3724 3027 3733
rect 2827 3720 3027 3724
rect 2827 3716 3024 3720
rect 3047 3716 5493 3724
rect 6676 3716 7133 3724
rect 1407 3696 1773 3704
rect 1787 3696 1833 3704
rect 2087 3696 2413 3704
rect 2427 3696 2593 3704
rect 2667 3696 2873 3704
rect 3067 3696 3284 3704
rect 567 3676 993 3684
rect 1007 3676 1033 3684
rect 1047 3676 1573 3684
rect 3027 3676 3253 3684
rect 3276 3684 3284 3696
rect 3307 3696 3373 3704
rect 3467 3696 3693 3704
rect 3847 3696 3913 3704
rect 4287 3696 4433 3704
rect 4487 3696 4892 3704
rect 4927 3696 5473 3704
rect 5567 3696 5693 3704
rect 5707 3696 5892 3704
rect 6676 3704 6684 3716
rect 7307 3716 7493 3724
rect 8187 3716 8313 3724
rect 8327 3716 8833 3724
rect 9447 3716 9613 3724
rect 5927 3696 6684 3704
rect 6756 3696 7324 3704
rect 3276 3676 3353 3684
rect 3407 3676 3533 3684
rect 6756 3684 6764 3696
rect 5167 3676 6764 3684
rect 6787 3676 6993 3684
rect 7316 3684 7324 3696
rect 7347 3696 7473 3704
rect 7487 3696 8093 3704
rect 8867 3696 8913 3704
rect 9087 3696 9253 3704
rect 11087 3696 11113 3704
rect 7316 3676 9013 3684
rect 9367 3676 9493 3684
rect 9507 3676 10353 3684
rect 10367 3676 10773 3684
rect 10787 3676 10813 3684
rect 10827 3676 11233 3684
rect 967 3656 993 3664
rect 1596 3656 1724 3664
rect 287 3636 513 3644
rect 1596 3644 1604 3656
rect 527 3636 1604 3644
rect 1716 3644 1724 3656
rect 1867 3656 2053 3664
rect 2227 3656 2493 3664
rect 2507 3656 2572 3664
rect 2607 3656 3673 3664
rect 3727 3656 4533 3664
rect 4967 3656 5453 3664
rect 5787 3656 6013 3664
rect 6467 3656 7073 3664
rect 7407 3656 7793 3664
rect 8287 3656 8373 3664
rect 10187 3656 10293 3664
rect 1716 3636 1933 3644
rect 2347 3636 2493 3644
rect 2947 3636 3153 3644
rect 3287 3636 3353 3644
rect 3407 3636 4853 3644
rect 5056 3636 5392 3644
rect 867 3616 973 3624
rect 1707 3616 2073 3624
rect 2207 3616 2513 3624
rect 2647 3616 2913 3624
rect 5056 3624 5064 3636
rect 5427 3636 5913 3644
rect 5987 3636 6233 3644
rect 6767 3636 6813 3644
rect 7507 3636 7893 3644
rect 8847 3636 8913 3644
rect 9067 3636 9253 3644
rect 4487 3616 5064 3624
rect 5087 3616 5933 3624
rect 5947 3616 6373 3624
rect 7187 3616 7433 3624
rect 9116 3616 10153 3624
rect 247 3596 473 3604
rect 487 3596 933 3604
rect 1587 3596 1733 3604
rect 1907 3596 2173 3604
rect 2187 3596 3473 3604
rect 3687 3596 4793 3604
rect 6733 3604 6747 3613
rect 6733 3600 7973 3604
rect 6736 3596 7973 3600
rect 8507 3596 8744 3604
rect 1347 3576 1853 3584
rect 1916 3580 2253 3584
rect 1913 3576 2253 3580
rect 1913 3567 1927 3576
rect 2587 3576 3273 3584
rect 3287 3576 3433 3584
rect 3627 3576 4713 3584
rect 4847 3576 5384 3584
rect 467 3556 573 3564
rect 587 3556 873 3564
rect 927 3556 1873 3564
rect 2407 3556 2533 3564
rect 2636 3556 3233 3564
rect 947 3536 1413 3544
rect 1607 3536 1653 3544
rect 1667 3536 1753 3544
rect 2636 3544 2644 3556
rect 3296 3556 3493 3564
rect 3296 3544 3304 3556
rect 3667 3556 3693 3564
rect 3887 3556 4473 3564
rect 4767 3556 5093 3564
rect 5376 3564 5384 3576
rect 5687 3576 5813 3584
rect 6247 3576 6273 3584
rect 6287 3576 6873 3584
rect 7027 3576 7513 3584
rect 7587 3576 7833 3584
rect 8267 3576 8473 3584
rect 8736 3584 8744 3596
rect 9116 3604 9124 3616
rect 9027 3596 9124 3604
rect 10327 3596 10413 3604
rect 8736 3576 9013 3584
rect 9367 3576 9953 3584
rect 5376 3556 5433 3564
rect 5887 3556 7253 3564
rect 7927 3556 7993 3564
rect 8447 3556 8533 3564
rect 9247 3556 9333 3564
rect 9827 3556 9893 3564
rect 10147 3556 10353 3564
rect 2587 3536 2644 3544
rect 2656 3536 3304 3544
rect 2656 3528 2664 3536
rect 3947 3536 4033 3544
rect 5527 3536 5633 3544
rect 5807 3536 6433 3544
rect 6727 3536 6933 3544
rect 7887 3536 8293 3544
rect 8307 3536 8553 3544
rect 8907 3536 8953 3544
rect 9916 3536 10073 3544
rect 9916 3528 9924 3536
rect 147 3476 173 3484
rect 196 3484 204 3514
rect 367 3516 413 3524
rect 607 3517 653 3525
rect 847 3517 873 3525
rect 967 3516 1113 3524
rect 1536 3516 1553 3524
rect 1536 3487 1544 3516
rect 1927 3517 1993 3525
rect 2247 3516 2273 3524
rect 1996 3504 2004 3514
rect 2467 3517 2493 3525
rect 2666 3514 2667 3528
rect 2687 3516 2833 3524
rect 3007 3516 3053 3524
rect 3147 3517 3313 3525
rect 2613 3504 2627 3513
rect 3316 3504 3324 3514
rect 3547 3516 3593 3524
rect 3636 3516 3904 3524
rect 3636 3504 3644 3516
rect 1996 3496 2164 3504
rect 2613 3500 2644 3504
rect 2616 3496 2644 3500
rect 3316 3496 3644 3504
rect 3896 3504 3904 3516
rect 4247 3517 4293 3525
rect 4387 3517 4433 3525
rect 4516 3516 4552 3524
rect 3896 3496 4053 3504
rect 196 3476 253 3484
rect 447 3476 673 3484
rect 767 3476 893 3484
rect 987 3475 1093 3483
rect 1587 3476 1693 3484
rect 1807 3476 1913 3484
rect 2156 3484 2164 3496
rect 2156 3476 2193 3484
rect 2447 3476 2573 3484
rect 2636 3486 2644 3496
rect 4516 3504 4524 3516
rect 4587 3516 4613 3524
rect 4667 3516 4733 3524
rect 4907 3517 4953 3525
rect 5027 3517 5073 3525
rect 5636 3516 5733 3524
rect 4476 3496 4524 3504
rect 3087 3475 3113 3483
rect 3527 3476 3613 3484
rect 3687 3476 4064 3484
rect 1247 3456 1393 3464
rect 1947 3456 1993 3464
rect 2227 3456 2313 3464
rect 2727 3456 3033 3464
rect 3167 3456 3253 3464
rect 3307 3456 3393 3464
rect 3447 3456 3564 3464
rect 1327 3436 1353 3444
rect 1867 3436 2753 3444
rect 2767 3436 3133 3444
rect 3556 3444 3564 3456
rect 3647 3456 3773 3464
rect 3887 3456 3913 3464
rect 4056 3464 4064 3476
rect 4476 3484 4484 3496
rect 4467 3476 4484 3484
rect 4547 3475 4633 3483
rect 4747 3475 4833 3483
rect 4887 3476 5013 3484
rect 5107 3476 5293 3484
rect 5636 3484 5644 3516
rect 6467 3524 6480 3527
rect 6467 3513 6484 3524
rect 7167 3517 7293 3525
rect 7567 3517 7593 3525
rect 7607 3516 7673 3524
rect 5547 3476 5644 3484
rect 6076 3484 6084 3494
rect 6207 3496 6293 3504
rect 6307 3496 6353 3504
rect 6476 3506 6484 3513
rect 5907 3476 6084 3484
rect 4056 3456 4333 3464
rect 4427 3456 4773 3464
rect 4907 3456 4973 3464
rect 6527 3456 6573 3464
rect 6716 3464 6724 3494
rect 6847 3496 7033 3504
rect 7116 3484 7124 3514
rect 7727 3517 7793 3525
rect 7947 3517 8013 3525
rect 9107 3520 9224 3524
rect 9107 3516 9227 3520
rect 7756 3496 8513 3504
rect 7116 3476 7353 3484
rect 7547 3476 7692 3484
rect 7756 3484 7764 3496
rect 7727 3476 7764 3484
rect 7787 3476 7933 3484
rect 8036 3486 8044 3496
rect 8607 3497 8753 3505
rect 9213 3507 9227 3516
rect 9627 3517 9793 3525
rect 9847 3517 9913 3525
rect 9967 3516 9993 3524
rect 10227 3517 10273 3525
rect 10367 3524 10380 3527
rect 10453 3524 10467 3533
rect 10367 3513 10384 3524
rect 8887 3496 9053 3504
rect 9347 3496 9513 3504
rect 9727 3496 10173 3504
rect 10376 3506 10384 3513
rect 10436 3520 10467 3524
rect 10436 3516 10464 3520
rect 10436 3504 10444 3516
rect 10407 3496 10444 3504
rect 10627 3497 10753 3505
rect 10796 3507 10804 3533
rect 10836 3507 10844 3553
rect 10836 3496 10853 3507
rect 10840 3493 10853 3496
rect 10896 3487 10904 3553
rect 11187 3536 11253 3544
rect 10913 3524 10927 3533
rect 10913 3520 10944 3524
rect 10916 3516 10944 3520
rect 9547 3476 9633 3484
rect 10067 3476 10212 3484
rect 10247 3476 10453 3484
rect 10467 3476 10733 3484
rect 6716 3456 7033 3464
rect 7107 3456 7153 3464
rect 7807 3456 7993 3464
rect 8107 3456 8453 3464
rect 8467 3456 8973 3464
rect 9027 3456 9253 3464
rect 9807 3456 9913 3464
rect 10267 3456 10333 3464
rect 10387 3456 10833 3464
rect 3556 3436 3933 3444
rect 4387 3436 4433 3444
rect 5287 3436 5313 3444
rect 5707 3436 5833 3444
rect 6187 3436 6313 3444
rect 7547 3436 7712 3444
rect 7747 3436 8212 3444
rect 8247 3436 9013 3444
rect 9027 3436 9093 3444
rect 9847 3436 9933 3444
rect 10207 3436 10293 3444
rect 10427 3436 10473 3444
rect 767 3416 953 3424
rect 2487 3416 2713 3424
rect 3207 3416 3253 3424
rect 5047 3416 5153 3424
rect 5236 3416 6313 3424
rect 5236 3407 5244 3416
rect 6887 3416 8513 3424
rect 9127 3416 9153 3424
rect 9687 3416 9733 3424
rect 10047 3416 10153 3424
rect 10347 3416 10393 3424
rect 10447 3416 10904 3424
rect 10896 3407 10904 3416
rect 1447 3396 1573 3404
rect 2847 3396 2893 3404
rect 2907 3396 3733 3404
rect 3887 3396 3952 3404
rect 3987 3396 4333 3404
rect 4547 3396 4853 3404
rect 4967 3396 5233 3404
rect 5767 3396 5893 3404
rect 6387 3396 6533 3404
rect 6547 3396 6593 3404
rect 6607 3396 6793 3404
rect 7047 3396 7313 3404
rect 7447 3396 7733 3404
rect 8227 3396 8493 3404
rect 8567 3396 9053 3404
rect 9476 3396 10193 3404
rect 227 3376 913 3384
rect 1367 3376 1853 3384
rect 1927 3376 2673 3384
rect 3147 3376 3964 3384
rect 1427 3356 1793 3364
rect 1967 3356 2353 3364
rect 2367 3356 2893 3364
rect 3127 3356 3233 3364
rect 3956 3364 3964 3376
rect 4367 3376 4913 3384
rect 5387 3376 5853 3384
rect 5867 3376 5913 3384
rect 6427 3376 6693 3384
rect 6927 3376 7593 3384
rect 7607 3376 7793 3384
rect 9476 3384 9484 3396
rect 10247 3396 10373 3404
rect 10467 3396 10513 3404
rect 10607 3396 10793 3404
rect 10896 3396 10913 3407
rect 10900 3393 10913 3396
rect 10936 3404 10944 3516
rect 11075 3407 11083 3494
rect 11096 3464 11104 3493
rect 11227 3496 11292 3504
rect 11196 3484 11204 3492
rect 11196 3476 11236 3484
rect 11096 3456 11193 3464
rect 11228 3425 11236 3476
rect 11315 3458 11324 3493
rect 11287 3450 11324 3458
rect 11228 3417 11293 3425
rect 10936 3396 11033 3404
rect 11127 3396 11193 3404
rect 7807 3376 9484 3384
rect 9587 3376 9733 3384
rect 9787 3376 10013 3384
rect 10027 3376 10133 3384
rect 10256 3376 10433 3384
rect 3956 3356 4453 3364
rect 4467 3356 4673 3364
rect 4696 3356 4833 3364
rect 967 3336 1253 3344
rect 1267 3336 1333 3344
rect 1927 3336 1973 3344
rect 2047 3336 2073 3344
rect 2087 3336 2173 3344
rect 2387 3336 2433 3344
rect 2576 3336 2833 3344
rect 1727 3316 1813 3324
rect 2027 3316 2053 3324
rect 2067 3316 2313 3324
rect 2407 3316 2433 3324
rect 2576 3324 2584 3336
rect 3067 3336 3513 3344
rect 3527 3336 3633 3344
rect 4107 3336 4253 3344
rect 4307 3336 4413 3344
rect 4587 3336 4612 3344
rect 4696 3344 4704 3356
rect 4847 3356 4993 3364
rect 5007 3356 5084 3364
rect 4647 3336 4704 3344
rect 5076 3347 5084 3356
rect 5127 3356 5653 3364
rect 6327 3356 6873 3364
rect 7687 3356 7773 3364
rect 7907 3356 8273 3364
rect 8507 3356 9633 3364
rect 9787 3356 9813 3364
rect 10256 3364 10264 3376
rect 10227 3356 10264 3364
rect 5076 3336 5093 3347
rect 5080 3333 5093 3336
rect 5147 3336 5273 3344
rect 5287 3336 5413 3344
rect 6567 3336 6613 3344
rect 7227 3336 7353 3344
rect 7367 3336 8293 3344
rect 8307 3336 8413 3344
rect 8427 3336 9273 3344
rect 9287 3336 9653 3344
rect 9667 3336 9853 3344
rect 9867 3336 10053 3344
rect 10067 3336 10093 3344
rect 10267 3336 10793 3344
rect 11147 3336 11213 3344
rect 2447 3316 2584 3324
rect 3327 3316 3353 3324
rect 3747 3316 3973 3324
rect 4347 3316 4393 3324
rect 4447 3316 5053 3324
rect 5347 3316 5453 3324
rect 6216 3316 6344 3324
rect 227 3297 273 3305
rect 176 3247 184 3294
rect 387 3296 413 3304
rect 467 3297 533 3305
rect 627 3297 673 3305
rect 1067 3297 1153 3305
rect 1167 3296 1373 3304
rect 207 3256 253 3264
rect 416 3247 424 3294
rect 1387 3296 1473 3304
rect 1647 3296 1873 3304
rect 1887 3296 1953 3304
rect 2367 3297 2633 3305
rect 2647 3296 2713 3304
rect 2787 3296 2933 3304
rect 3027 3297 3133 3305
rect 3427 3297 3473 3305
rect 3567 3297 3613 3305
rect 3667 3296 3713 3304
rect 4047 3297 4093 3305
rect 4227 3297 4313 3305
rect 4567 3296 4693 3304
rect 4707 3296 4793 3304
rect 4867 3297 4953 3305
rect 4967 3297 5013 3305
rect 5067 3297 5193 3305
rect 5507 3296 5553 3304
rect 5607 3297 5733 3305
rect 5967 3296 6073 3304
rect 6216 3304 6224 3316
rect 6207 3296 6224 3304
rect 6336 3304 6344 3316
rect 6827 3316 7033 3324
rect 7387 3316 7713 3324
rect 8187 3316 8253 3324
rect 8467 3316 8553 3324
rect 8867 3316 8973 3324
rect 9427 3316 9573 3324
rect 9887 3316 9913 3324
rect 10627 3316 10813 3324
rect 11187 3316 11264 3324
rect 6336 3296 6584 3304
rect 1807 3276 2813 3284
rect 3047 3276 3453 3284
rect 4527 3276 4933 3284
rect 6287 3276 6313 3284
rect 6576 3284 6584 3296
rect 6727 3296 7073 3304
rect 7147 3296 7313 3304
rect 7547 3296 7593 3304
rect 7696 3296 7753 3304
rect 6576 3276 6604 3284
rect 547 3256 653 3264
rect 727 3255 753 3263
rect 1267 3256 1293 3264
rect 1467 3256 1633 3264
rect 1847 3256 2073 3264
rect 2327 3255 2453 3263
rect 2667 3255 2733 3263
rect 2927 3255 2953 3263
rect 407 3236 424 3247
rect 407 3233 420 3236
rect 447 3236 513 3244
rect 967 3236 993 3244
rect 1387 3236 1713 3244
rect 1787 3236 2153 3244
rect 2167 3236 2573 3244
rect 2976 3244 2984 3273
rect 3127 3255 3233 3263
rect 3547 3256 3593 3264
rect 3687 3256 3853 3264
rect 3876 3256 4113 3264
rect 2976 3236 3033 3244
rect 3347 3236 3373 3244
rect 3876 3244 3884 3256
rect 4727 3255 4773 3263
rect 5107 3256 5513 3264
rect 5527 3256 5633 3264
rect 5647 3256 5693 3264
rect 5707 3256 5793 3264
rect 6427 3256 6553 3264
rect 6596 3264 6604 3276
rect 7696 3267 7704 3296
rect 7780 3304 7793 3307
rect 7776 3293 7793 3304
rect 8776 3300 9133 3304
rect 8773 3296 9133 3300
rect 6596 3256 6713 3264
rect 6887 3256 6973 3264
rect 7107 3255 7133 3263
rect 7347 3255 7553 3263
rect 7776 3266 7784 3293
rect 3627 3236 3884 3244
rect 3927 3236 4173 3244
rect 4196 3236 5033 3244
rect 587 3216 913 3224
rect 1027 3216 1153 3224
rect 1167 3216 1313 3224
rect 1427 3216 1513 3224
rect 1907 3216 2013 3224
rect 2227 3216 2313 3224
rect 2827 3216 3293 3224
rect 4196 3224 4204 3236
rect 5167 3236 5273 3244
rect 5287 3236 5473 3244
rect 6167 3236 6253 3244
rect 6267 3235 6313 3243
rect 7307 3236 7373 3244
rect 7607 3236 7733 3244
rect 7856 3244 7864 3293
rect 8056 3280 8173 3284
rect 8053 3276 8173 3280
rect 8053 3267 8067 3276
rect 8476 3276 8513 3284
rect 8476 3266 8484 3276
rect 8773 3287 8787 3296
rect 9187 3297 9213 3305
rect 9307 3296 9373 3304
rect 9627 3296 9713 3304
rect 9907 3296 9933 3304
rect 10007 3296 10093 3304
rect 10847 3297 10973 3305
rect 11087 3296 11213 3304
rect 8593 3264 8607 3273
rect 9796 3267 9804 3293
rect 11256 3267 11264 3316
rect 8593 3260 8753 3264
rect 8596 3256 8753 3260
rect 8896 3260 8953 3264
rect 8893 3256 8953 3260
rect 8893 3247 8907 3256
rect 9267 3255 9353 3263
rect 9527 3256 9593 3264
rect 10027 3255 10113 3263
rect 11007 3256 11093 3264
rect 7807 3236 7864 3244
rect 8087 3236 8193 3244
rect 8247 3236 8313 3244
rect 9007 3244 9020 3247
rect 9007 3233 9024 3244
rect 9087 3236 9173 3244
rect 9927 3236 10253 3244
rect 10887 3236 11193 3244
rect 3467 3216 4204 3224
rect 4267 3216 4413 3224
rect 4587 3216 4733 3224
rect 4747 3216 4813 3224
rect 5667 3216 5933 3224
rect 7067 3216 7513 3224
rect 8367 3216 8513 3224
rect 9016 3224 9024 3233
rect 9016 3216 9153 3224
rect 9227 3216 9613 3224
rect 10567 3216 10613 3224
rect 10907 3216 11153 3224
rect 1207 3196 1533 3204
rect 1667 3196 1873 3204
rect 2087 3196 2233 3204
rect 2627 3196 3093 3204
rect 3847 3196 4513 3204
rect 4927 3196 6213 3204
rect 7667 3196 7832 3204
rect 7867 3196 8313 3204
rect 9007 3196 9193 3204
rect 9207 3196 9633 3204
rect 9647 3196 9793 3204
rect 9807 3196 10073 3204
rect 10787 3196 10853 3204
rect 10927 3196 11073 3204
rect 547 3176 813 3184
rect 927 3176 1584 3184
rect 1576 3164 1584 3176
rect 1687 3176 1833 3184
rect 2327 3176 3113 3184
rect 3587 3176 3793 3184
rect 3887 3176 4633 3184
rect 4827 3176 4893 3184
rect 4967 3176 5013 3184
rect 5307 3176 5373 3184
rect 5567 3176 6093 3184
rect 6707 3176 7433 3184
rect 7707 3176 8433 3184
rect 8447 3176 8973 3184
rect 9047 3176 9113 3184
rect 10507 3176 10753 3184
rect 1576 3156 2213 3164
rect 2587 3156 2864 3164
rect 1147 3136 1573 3144
rect 1727 3136 1813 3144
rect 2027 3136 2193 3144
rect 2287 3136 2553 3144
rect 2856 3144 2864 3156
rect 2907 3156 3093 3164
rect 3907 3156 3993 3164
rect 4727 3156 5373 3164
rect 6947 3156 7073 3164
rect 7467 3156 7493 3164
rect 9687 3156 9973 3164
rect 10407 3156 10913 3164
rect 2856 3136 3553 3144
rect 3607 3136 3873 3144
rect 4067 3136 4093 3144
rect 4407 3136 5133 3144
rect 5887 3136 7153 3144
rect 7247 3136 7273 3144
rect 7627 3136 8953 3144
rect 9527 3136 11053 3144
rect 247 3116 633 3124
rect 647 3116 833 3124
rect 847 3116 873 3124
rect 887 3116 1953 3124
rect 1967 3116 2413 3124
rect 2427 3116 2853 3124
rect 2907 3116 3133 3124
rect 3147 3116 3472 3124
rect 3507 3116 3613 3124
rect 3947 3116 4033 3124
rect 4527 3116 5153 3124
rect 5627 3116 5713 3124
rect 8467 3116 8553 3124
rect 8627 3116 8913 3124
rect 9607 3116 9873 3124
rect 10007 3116 10733 3124
rect 487 3096 553 3104
rect 827 3096 1753 3104
rect 1827 3096 1933 3104
rect 1987 3096 2253 3104
rect 2827 3096 3013 3104
rect 3227 3096 3833 3104
rect 4007 3096 5173 3104
rect 8947 3096 9493 3104
rect 9567 3096 9673 3104
rect 1327 3076 2373 3084
rect 2467 3076 2533 3084
rect 2647 3076 2753 3084
rect 3307 3076 3713 3084
rect 4047 3076 4673 3084
rect 4687 3076 4893 3084
rect 4947 3076 5293 3084
rect 5487 3076 5593 3084
rect 6607 3076 7173 3084
rect 7487 3076 7553 3084
rect 7887 3076 8273 3084
rect 8387 3076 9513 3084
rect 347 3056 593 3064
rect 667 3056 1124 3064
rect 1116 3044 1124 3056
rect 1307 3056 1793 3064
rect 1847 3056 2012 3064
rect 2047 3056 2404 3064
rect 1116 3036 1313 3044
rect 2396 3044 2404 3056
rect 2427 3056 2552 3064
rect 2587 3056 3073 3064
rect 3127 3056 3853 3064
rect 3867 3056 3993 3064
rect 4047 3056 4073 3064
rect 4147 3056 4553 3064
rect 5416 3056 6173 3064
rect 1647 3036 1784 3044
rect 2396 3036 2893 3044
rect 1776 3024 1784 3036
rect 5416 3044 5424 3056
rect 7787 3056 8353 3064
rect 8427 3056 8813 3064
rect 9027 3056 9093 3064
rect 9707 3056 9853 3064
rect 10527 3056 11093 3064
rect 3007 3036 5424 3044
rect 5447 3036 5913 3044
rect 6327 3036 6733 3044
rect 6927 3036 6993 3044
rect 8047 3036 8344 3044
rect 1776 3016 1933 3024
rect 2167 3016 2304 3024
rect 747 2996 933 3004
rect 1347 2996 1373 3004
rect 1387 2997 1453 3005
rect 1507 2996 1713 3004
rect 2296 3007 2304 3016
rect 2407 3016 2493 3024
rect 2707 3016 2753 3024
rect 3407 3016 3553 3024
rect 3707 3016 4033 3024
rect 4087 3016 4433 3024
rect 4507 3016 4553 3024
rect 4707 3016 4773 3024
rect 5407 3016 5933 3024
rect 7487 3016 7633 3024
rect 7647 3016 7773 3024
rect 8336 3024 8344 3036
rect 9336 3036 9373 3044
rect 8336 3016 8404 3024
rect 1727 2996 1873 3004
rect 2296 2996 2313 3007
rect 2300 2993 2313 2996
rect 2367 2996 2573 3004
rect 2647 2997 2713 3005
rect 2947 2997 2993 3005
rect 3087 2997 3173 3005
rect 3200 3004 3213 3007
rect 3196 2993 3213 3004
rect 3436 3000 3573 3004
rect 3433 2996 3573 3000
rect 1496 2976 2053 2984
rect 387 2955 433 2963
rect 1327 2956 1473 2964
rect 1496 2964 1504 2976
rect 1487 2956 1504 2964
rect 1527 2956 1633 2964
rect 1647 2955 1693 2963
rect 2007 2956 2073 2964
rect 2087 2956 2173 2964
rect 2327 2955 2433 2963
rect 2487 2956 2633 2964
rect 2787 2955 2913 2963
rect 3196 2966 3204 2993
rect 3433 2987 3447 2996
rect 3647 2997 3673 3005
rect 3987 2997 4053 3005
rect 4187 2996 4313 3004
rect 4907 2997 4933 3005
rect 5067 2997 5133 3005
rect 5187 2996 5833 3004
rect 6007 2997 6113 3005
rect 6127 2996 6273 3004
rect 6547 2996 6633 3004
rect 7927 2996 7973 3004
rect 8027 2997 8093 3005
rect 4113 2984 4127 2993
rect 4113 2980 4333 2984
rect 4116 2976 4333 2980
rect 3007 2956 3153 2964
rect 3607 2955 3653 2963
rect 3947 2955 4033 2963
rect 4407 2955 4493 2963
rect 4927 2955 5013 2963
rect 5027 2956 5193 2964
rect 5587 2956 5813 2964
rect 5867 2956 5993 2964
rect 6247 2955 6293 2963
rect 6647 2955 6713 2963
rect 7327 2955 7433 2963
rect 7447 2956 7653 2964
rect 7907 2956 8033 2964
rect 8136 2964 8144 2994
rect 8307 2996 8364 3004
rect 8136 2956 8333 2964
rect 8356 2964 8364 2996
rect 8396 2984 8404 3016
rect 9147 3016 9233 3024
rect 8987 2996 9013 3004
rect 9207 3004 9220 3007
rect 9260 3004 9273 3007
rect 9207 2993 9224 3004
rect 8396 2976 8413 2984
rect 8356 2956 8373 2964
rect 8656 2964 8664 2974
rect 8787 2976 8853 2984
rect 8467 2956 8664 2964
rect 9067 2956 9133 2964
rect 9216 2966 9224 2993
rect 9256 2993 9273 3004
rect 9336 3004 9344 3036
rect 9416 3036 9533 3044
rect 9416 3024 9424 3036
rect 10087 3036 10413 3044
rect 9316 3000 9344 3004
rect 9313 2996 9344 3000
rect 9356 3016 9424 3024
rect 9256 2966 9264 2993
rect 9313 2987 9327 2996
rect 9356 2986 9364 3016
rect 9727 3016 9753 3024
rect 10787 3024 10800 3027
rect 10787 3013 10804 3024
rect 10947 3016 10973 3024
rect 11187 3016 11253 3024
rect 9847 2996 10093 3004
rect 9407 2977 9533 2985
rect 9667 2976 9813 2984
rect 10247 2977 10392 2985
rect 10596 2987 10604 3013
rect 10427 2976 10513 2984
rect 10647 2977 10773 2985
rect 907 2936 1052 2944
rect 1087 2936 1113 2944
rect 1127 2936 1273 2944
rect 1387 2936 1453 2944
rect 1847 2936 1933 2944
rect 2627 2936 2673 2944
rect 3827 2936 3913 2944
rect 4107 2936 4173 2944
rect 4247 2936 4273 2944
rect 4327 2936 4353 2944
rect 4887 2936 4973 2944
rect 5267 2936 5553 2944
rect 5787 2936 7253 2944
rect 7527 2936 7644 2944
rect 847 2916 1173 2924
rect 2107 2916 2213 2924
rect 3007 2916 3673 2924
rect 3967 2916 4113 2924
rect 4447 2916 5052 2924
rect 5087 2916 5393 2924
rect 5867 2916 5973 2924
rect 6427 2916 6713 2924
rect 6767 2916 6993 2924
rect 7287 2916 7453 2924
rect 7636 2924 7644 2936
rect 8127 2936 8193 2944
rect 9307 2936 9913 2944
rect 10107 2936 10193 2944
rect 10796 2944 10804 3013
rect 10967 2975 11073 2983
rect 10627 2936 10804 2944
rect 7636 2916 8353 2924
rect 9187 2916 9273 2924
rect 9647 2916 9833 2924
rect 10947 2916 11193 2924
rect 207 2896 653 2904
rect 876 2896 1013 2904
rect 876 2884 884 2896
rect 1027 2896 1113 2904
rect 1227 2896 1393 2904
rect 1507 2896 1613 2904
rect 1967 2896 2033 2904
rect 2107 2896 2293 2904
rect 2347 2896 2813 2904
rect 3047 2896 3153 2904
rect 3207 2896 3253 2904
rect 3747 2896 4213 2904
rect 4667 2896 4753 2904
rect 4867 2896 5373 2904
rect 5527 2896 6233 2904
rect 8087 2896 8113 2904
rect 8907 2896 9133 2904
rect 9327 2900 9584 2904
rect 9327 2896 9587 2900
rect 807 2876 884 2884
rect 1047 2876 1153 2884
rect 2816 2884 2824 2893
rect 9573 2887 9587 2896
rect 10047 2896 10113 2904
rect 10647 2896 10993 2904
rect 2816 2876 3613 2884
rect 3627 2876 4813 2884
rect 5207 2876 5313 2884
rect 5327 2876 5533 2884
rect 5627 2876 6093 2884
rect 7287 2876 7413 2884
rect 8367 2876 8533 2884
rect 8587 2876 8753 2884
rect 8927 2876 9213 2884
rect 10207 2876 10233 2884
rect 10607 2876 10633 2884
rect 10887 2876 11033 2884
rect 11207 2876 11273 2884
rect 496 2856 893 2864
rect 496 2844 504 2856
rect 907 2856 933 2864
rect 947 2856 1953 2864
rect 2087 2856 2293 2864
rect 3027 2856 3973 2864
rect 4027 2856 4153 2864
rect 4407 2856 4733 2864
rect 4827 2856 4872 2864
rect 4907 2856 5293 2864
rect 6127 2856 6564 2864
rect 147 2836 504 2844
rect 527 2836 1733 2844
rect 2067 2836 3384 2844
rect 847 2816 873 2824
rect 1987 2816 2473 2824
rect 2556 2816 3053 2824
rect 2556 2807 2564 2816
rect 3376 2824 3384 2836
rect 3427 2836 3753 2844
rect 4187 2836 4693 2844
rect 4787 2836 5313 2844
rect 6556 2844 6564 2856
rect 7247 2856 7524 2864
rect 7516 2847 7524 2856
rect 7727 2856 8193 2864
rect 8347 2856 8453 2864
rect 9067 2856 9173 2864
rect 9187 2856 9413 2864
rect 9607 2856 9733 2864
rect 10627 2856 10713 2864
rect 6556 2836 6933 2844
rect 7527 2836 7933 2844
rect 8227 2836 8253 2844
rect 8487 2836 8993 2844
rect 9007 2836 9533 2844
rect 9847 2836 10773 2844
rect 3376 2816 3693 2824
rect 4207 2816 4293 2824
rect 4447 2816 4833 2824
rect 5707 2816 6113 2824
rect 6547 2816 6833 2824
rect 8207 2816 8453 2824
rect 8627 2816 9013 2824
rect 9887 2816 9953 2824
rect 10227 2816 10373 2824
rect 10387 2816 10953 2824
rect 11027 2816 11273 2824
rect 187 2796 233 2804
rect 647 2796 973 2804
rect 987 2796 1073 2804
rect 1967 2796 2353 2804
rect 2447 2796 2553 2804
rect 2607 2796 2653 2804
rect 4007 2796 4053 2804
rect 4267 2796 4853 2804
rect 5127 2796 5153 2804
rect 5307 2796 5332 2804
rect 5367 2796 5613 2804
rect 7407 2796 7893 2804
rect 9147 2796 9633 2804
rect 9647 2796 9673 2804
rect 10467 2796 10493 2804
rect 10507 2796 10813 2804
rect 11227 2796 11253 2804
rect 227 2776 353 2784
rect 656 2776 673 2784
rect 656 2764 664 2776
rect 1087 2777 1153 2785
rect 1607 2777 1633 2785
rect 2007 2776 2233 2784
rect 2247 2777 2273 2785
rect 2667 2776 2684 2784
rect 236 2756 664 2764
rect 236 2746 244 2756
rect 1747 2756 2613 2764
rect 2676 2764 2684 2776
rect 2707 2776 2853 2784
rect 3107 2776 3133 2784
rect 2676 2756 3213 2764
rect 3296 2764 3304 2774
rect 3347 2776 3513 2784
rect 3527 2776 3853 2784
rect 4127 2777 4213 2785
rect 3296 2756 3553 2764
rect 3567 2756 3873 2764
rect 3936 2747 3944 2774
rect 3976 2764 3984 2774
rect 4347 2776 4432 2784
rect 4467 2776 4493 2784
rect 4647 2776 4793 2784
rect 4927 2777 5173 2785
rect 5187 2777 5213 2785
rect 5467 2776 5573 2784
rect 5767 2777 5793 2785
rect 5987 2776 6013 2784
rect 6027 2777 6073 2785
rect 6147 2776 6273 2784
rect 6287 2776 6413 2784
rect 6427 2777 6493 2785
rect 6647 2777 6673 2785
rect 7156 2776 7353 2784
rect 3976 2756 4033 2764
rect 7156 2764 7164 2776
rect 7027 2756 7164 2764
rect 367 2735 413 2743
rect 847 2735 873 2743
rect 1147 2736 1193 2744
rect 1207 2736 1333 2744
rect 1407 2736 1633 2744
rect 1787 2735 1873 2743
rect 1887 2736 2073 2744
rect 2207 2736 2253 2744
rect 2367 2735 2413 2743
rect 2767 2736 3013 2744
rect 3027 2736 3073 2744
rect 3127 2736 3793 2744
rect 3927 2736 3944 2747
rect 3927 2733 3940 2736
rect 4087 2736 4224 2744
rect 467 2716 513 2724
rect 567 2716 673 2724
rect 1067 2716 1113 2724
rect 1676 2716 2173 2724
rect 407 2696 533 2704
rect 1676 2704 1684 2716
rect 2547 2716 3473 2724
rect 4216 2724 4224 2736
rect 4307 2735 4373 2743
rect 4467 2736 4553 2744
rect 4767 2735 4853 2743
rect 4967 2735 5093 2743
rect 5367 2735 5453 2743
rect 5647 2735 5693 2743
rect 6087 2736 6253 2744
rect 6487 2736 6533 2744
rect 6707 2735 6853 2743
rect 6967 2735 6993 2743
rect 7187 2736 7213 2744
rect 7356 2727 7364 2774
rect 7967 2776 8073 2784
rect 8127 2777 8153 2785
rect 8287 2777 8373 2785
rect 8467 2776 9053 2784
rect 9507 2777 9553 2785
rect 9767 2777 9913 2785
rect 10067 2777 10333 2785
rect 10587 2777 10733 2785
rect 10907 2776 10973 2784
rect 7456 2744 7464 2754
rect 7847 2756 7913 2764
rect 9067 2756 9153 2764
rect 7427 2736 7464 2744
rect 7907 2735 8053 2743
rect 8107 2736 8313 2744
rect 8507 2736 8553 2744
rect 8973 2744 8987 2753
rect 8567 2740 8987 2744
rect 8567 2736 8984 2740
rect 9027 2736 9473 2744
rect 9707 2736 10033 2744
rect 10107 2736 10133 2744
rect 10567 2736 10913 2744
rect 11056 2744 11064 2774
rect 11056 2736 11233 2744
rect 4216 2716 4713 2724
rect 5127 2716 5253 2724
rect 5827 2716 6013 2724
rect 6027 2716 6053 2724
rect 7447 2716 7853 2724
rect 9047 2716 9233 2724
rect 9247 2716 9253 2724
rect 10327 2716 10513 2724
rect 10947 2716 11033 2724
rect 1187 2696 1684 2704
rect 2007 2696 2093 2704
rect 2367 2696 2593 2704
rect 2807 2696 2853 2704
rect 3107 2696 3753 2704
rect 3767 2696 3813 2704
rect 4227 2696 4793 2704
rect 4927 2696 5273 2704
rect 5407 2696 5793 2704
rect 5847 2696 5993 2704
rect 7387 2696 7413 2704
rect 7887 2696 8253 2704
rect 9767 2696 9813 2704
rect 9836 2696 10113 2704
rect 707 2676 2793 2684
rect 2887 2676 3313 2684
rect 3327 2676 3453 2684
rect 3507 2676 4273 2684
rect 4287 2676 4533 2684
rect 4827 2676 4893 2684
rect 5067 2676 5593 2684
rect 7067 2676 7213 2684
rect 7867 2676 8013 2684
rect 8187 2676 8213 2684
rect 8367 2676 8553 2684
rect 9836 2684 9844 2696
rect 10127 2696 10793 2704
rect 9307 2676 9844 2684
rect 11007 2676 11053 2684
rect 1207 2656 2333 2664
rect 2387 2656 2533 2664
rect 3087 2656 3193 2664
rect 3627 2656 4313 2664
rect 4847 2656 4993 2664
rect 5216 2656 5573 2664
rect 287 2636 313 2644
rect 447 2636 1073 2644
rect 1127 2636 1373 2644
rect 1387 2636 1933 2644
rect 1947 2636 2093 2644
rect 3687 2636 4213 2644
rect 5216 2644 5224 2656
rect 6487 2656 6873 2664
rect 8267 2656 8653 2664
rect 9567 2656 9733 2664
rect 10727 2656 10953 2664
rect 4807 2636 5224 2644
rect 5247 2636 5273 2644
rect 5696 2636 6313 2644
rect 527 2616 653 2624
rect 667 2616 813 2624
rect 1807 2616 2153 2624
rect 2496 2616 2613 2624
rect 2496 2604 2504 2616
rect 3167 2616 3273 2624
rect 3867 2616 4313 2624
rect 5696 2624 5704 2636
rect 6327 2636 6393 2644
rect 7707 2636 7953 2644
rect 8136 2636 8193 2644
rect 4367 2616 5704 2624
rect 6427 2616 7013 2624
rect 7087 2616 7333 2624
rect 8136 2624 8144 2636
rect 9427 2636 10993 2644
rect 7767 2616 8144 2624
rect 8887 2616 9133 2624
rect 9407 2616 9893 2624
rect 11027 2616 11153 2624
rect 876 2596 2504 2604
rect 876 2584 884 2596
rect 2527 2596 2993 2604
rect 3047 2596 3333 2604
rect 3807 2596 4253 2604
rect 4727 2596 5013 2604
rect 5167 2596 5233 2604
rect 5247 2596 5753 2604
rect 6747 2596 7053 2604
rect 7167 2596 7293 2604
rect 7747 2596 8153 2604
rect 8727 2593 8733 2607
rect 9987 2596 10173 2604
rect 10587 2596 10673 2604
rect 547 2576 884 2584
rect 907 2576 1233 2584
rect 1927 2576 2173 2584
rect 2347 2576 3653 2584
rect 3667 2576 3753 2584
rect 3836 2576 4213 2584
rect 467 2556 1793 2564
rect 2747 2556 2833 2564
rect 3027 2556 3433 2564
rect 3836 2564 3844 2576
rect 4327 2576 7313 2584
rect 7327 2576 7453 2584
rect 8927 2576 9193 2584
rect 9307 2576 9613 2584
rect 10087 2576 10253 2584
rect 10267 2576 10473 2584
rect 3487 2556 3844 2564
rect 3856 2556 5193 2564
rect 547 2536 893 2544
rect 1127 2536 1473 2544
rect 1787 2536 2013 2544
rect 2207 2536 2453 2544
rect 3856 2544 3864 2556
rect 6716 2556 7153 2564
rect 6716 2547 6724 2556
rect 8247 2556 8333 2564
rect 8647 2556 9173 2564
rect 9287 2556 9813 2564
rect 2667 2536 3864 2544
rect 4227 2536 4273 2544
rect 5007 2536 5213 2544
rect 5587 2536 5673 2544
rect 5687 2536 6173 2544
rect 6287 2536 6633 2544
rect 6647 2536 6713 2544
rect 7147 2536 7693 2544
rect 7947 2536 8313 2544
rect 8807 2536 9033 2544
rect 9107 2536 9973 2544
rect 11187 2536 11253 2544
rect 947 2516 1233 2524
rect 1547 2516 1633 2524
rect 2047 2516 2073 2524
rect 2087 2516 2133 2524
rect 2907 2516 3413 2524
rect 3887 2516 4073 2524
rect 4267 2516 4293 2524
rect 4307 2516 4413 2524
rect 4907 2516 4973 2524
rect 5267 2516 6233 2524
rect 6787 2516 7433 2524
rect 7927 2516 8473 2524
rect 9227 2516 9673 2524
rect 10267 2516 10353 2524
rect 11207 2516 11273 2524
rect 607 2496 773 2504
rect 1867 2496 2253 2504
rect 2647 2496 2693 2504
rect 4787 2496 4853 2504
rect 5027 2496 5173 2504
rect 6547 2496 6753 2504
rect 6927 2496 7193 2504
rect 7647 2496 8353 2504
rect 8787 2496 9033 2504
rect 9867 2496 9893 2504
rect 10547 2496 10593 2504
rect 187 2477 333 2485
rect 647 2477 753 2485
rect 867 2476 1053 2484
rect 1267 2477 1293 2485
rect 1347 2477 1393 2485
rect 1507 2476 1573 2484
rect 1600 2484 1613 2487
rect 1596 2473 1613 2484
rect 1827 2477 1973 2485
rect 2347 2477 2473 2485
rect 2587 2477 2733 2485
rect 3067 2477 3173 2485
rect 3427 2476 3613 2484
rect 3827 2476 3873 2484
rect 127 2436 193 2444
rect 387 2436 453 2444
rect 507 2436 573 2444
rect 887 2435 933 2443
rect 1107 2436 1313 2444
rect 1367 2435 1433 2443
rect 1596 2446 1604 2473
rect 2796 2456 2893 2464
rect 1487 2436 1553 2444
rect 2287 2436 2313 2444
rect 2327 2436 2633 2444
rect 2796 2444 2804 2456
rect 2727 2436 2804 2444
rect 2936 2427 2944 2474
rect 3376 2464 3384 2474
rect 3947 2477 4013 2485
rect 4080 2484 4093 2487
rect 4076 2473 4093 2484
rect 4227 2477 4253 2485
rect 4367 2476 4473 2484
rect 4687 2476 4753 2484
rect 4967 2476 5093 2484
rect 5156 2476 5193 2484
rect 3376 2456 3513 2464
rect 2967 2435 2993 2443
rect 3287 2436 3433 2444
rect 4076 2446 4084 2473
rect 5156 2446 5164 2476
rect 5327 2476 5373 2484
rect 5396 2476 5593 2484
rect 5396 2446 5404 2476
rect 5707 2477 5753 2485
rect 5807 2477 5893 2485
rect 7547 2477 7593 2485
rect 7707 2476 7813 2484
rect 8627 2477 8693 2485
rect 9427 2476 9553 2484
rect 9567 2476 9593 2484
rect 10307 2476 10433 2484
rect 10447 2477 10493 2485
rect 10827 2477 11173 2485
rect 6087 2456 6813 2464
rect 6827 2455 7093 2463
rect 7167 2455 7213 2463
rect 7853 2464 7867 2473
rect 7853 2460 7893 2464
rect 7856 2456 7893 2460
rect 7967 2457 8113 2465
rect 8247 2456 8553 2464
rect 3807 2435 3993 2443
rect 4087 2440 4304 2444
rect 4087 2436 4307 2440
rect 4293 2427 4307 2436
rect 4567 2435 4593 2443
rect 4827 2435 4933 2443
rect 4987 2435 5013 2443
rect 5336 2436 5353 2444
rect 687 2416 833 2424
rect 2767 2416 2813 2424
rect 3167 2416 3364 2424
rect 1247 2396 1753 2404
rect 3207 2396 3333 2404
rect 3356 2404 3364 2416
rect 5336 2424 5344 2436
rect 6267 2436 6593 2444
rect 7267 2435 7313 2443
rect 7327 2435 7393 2443
rect 7667 2435 7693 2443
rect 7847 2436 7873 2444
rect 8956 2444 8964 2473
rect 9047 2456 9273 2464
rect 8907 2436 8964 2444
rect 9036 2444 9044 2453
rect 9176 2446 9184 2456
rect 10147 2456 10324 2464
rect 8987 2436 9044 2444
rect 9227 2435 9293 2443
rect 9347 2435 9393 2443
rect 9667 2436 9773 2444
rect 10316 2446 10324 2456
rect 11216 2447 11224 2474
rect 9867 2436 10033 2444
rect 10447 2436 10473 2444
rect 10567 2436 10613 2444
rect 11216 2436 11233 2447
rect 11220 2433 11233 2436
rect 5107 2416 5344 2424
rect 6447 2416 6673 2424
rect 8227 2416 8273 2424
rect 8527 2416 8593 2424
rect 8727 2416 9113 2424
rect 9447 2416 9593 2424
rect 10207 2416 10273 2424
rect 10367 2416 10513 2424
rect 10967 2416 11013 2424
rect 11087 2416 11173 2424
rect 3356 2396 3473 2404
rect 3647 2396 3893 2404
rect 3987 2396 4013 2404
rect 4387 2396 5033 2404
rect 6027 2396 6153 2404
rect 7087 2396 7233 2404
rect 7627 2396 7953 2404
rect 8827 2396 8933 2404
rect 10436 2396 10753 2404
rect 807 2376 1032 2384
rect 1067 2376 1093 2384
rect 3007 2376 3233 2384
rect 3767 2376 3833 2384
rect 4527 2376 4912 2384
rect 4947 2376 4973 2384
rect 5387 2376 5433 2384
rect 5947 2376 6313 2384
rect 8267 2376 8333 2384
rect 8507 2376 9193 2384
rect 9467 2376 9513 2384
rect 9967 2376 10033 2384
rect 10436 2384 10444 2396
rect 11207 2396 11293 2404
rect 10047 2376 10444 2384
rect 10467 2376 10513 2384
rect 10947 2376 11033 2384
rect 647 2356 693 2364
rect 1367 2356 1453 2364
rect 1967 2356 2073 2364
rect 2227 2356 2764 2364
rect 787 2336 1013 2344
rect 1027 2336 1093 2344
rect 1267 2336 2373 2344
rect 2756 2344 2764 2356
rect 2787 2356 2953 2364
rect 4007 2356 4072 2364
rect 4107 2356 4273 2364
rect 4347 2356 4533 2364
rect 4687 2356 5833 2364
rect 5847 2356 6213 2364
rect 7227 2356 7433 2364
rect 8007 2356 8244 2364
rect 8236 2347 8244 2356
rect 9027 2356 9173 2364
rect 9407 2356 9433 2364
rect 10976 2356 11153 2364
rect 10976 2347 10984 2356
rect 11227 2356 11333 2364
rect 2756 2336 3553 2344
rect 3567 2336 3593 2344
rect 3787 2336 3973 2344
rect 4016 2336 4253 2344
rect 627 2316 873 2324
rect 1387 2316 1493 2324
rect 1847 2316 2193 2324
rect 2447 2316 2553 2324
rect 2627 2316 3113 2324
rect 4016 2324 4024 2336
rect 4307 2336 4733 2344
rect 4747 2336 4873 2344
rect 4927 2336 5993 2344
rect 6807 2336 6893 2344
rect 7027 2336 7533 2344
rect 8247 2336 8313 2344
rect 9087 2336 9693 2344
rect 9747 2336 10273 2344
rect 10287 2336 10593 2344
rect 10607 2336 10853 2344
rect 10867 2336 10973 2344
rect 3307 2316 4024 2324
rect 4047 2316 4213 2324
rect 4427 2316 4753 2324
rect 4967 2316 5113 2324
rect 5316 2316 5693 2324
rect 207 2296 573 2304
rect 727 2296 833 2304
rect 1047 2296 1553 2304
rect 1567 2296 1873 2304
rect 1927 2296 1993 2304
rect 2007 2296 3273 2304
rect 3336 2296 3393 2304
rect 187 2276 313 2284
rect 327 2276 533 2284
rect 887 2276 953 2284
rect 1127 2276 1633 2284
rect 1647 2276 1724 2284
rect 1716 2268 1724 2276
rect 2027 2276 2352 2284
rect 2387 2276 2413 2284
rect 2507 2276 2653 2284
rect 2667 2276 2693 2284
rect 227 2257 253 2265
rect 767 2256 1033 2264
rect 1307 2256 1513 2264
rect 1727 2257 1753 2265
rect 1807 2257 1833 2265
rect 2187 2256 2273 2264
rect 2487 2256 2644 2264
rect 147 2216 193 2224
rect 376 2224 384 2253
rect 2636 2244 2644 2256
rect 2827 2257 2893 2265
rect 2967 2256 3153 2264
rect 3167 2257 3253 2265
rect 2636 2236 2684 2244
rect 376 2216 413 2224
rect 587 2215 613 2223
rect 627 2216 753 2224
rect 967 2216 1073 2224
rect 1096 2216 1153 2224
rect 1096 2204 1104 2216
rect 1247 2215 1573 2223
rect 1587 2216 1653 2224
rect 2027 2216 2073 2224
rect 2676 2226 2684 2236
rect 2167 2215 2193 2223
rect 2387 2215 2413 2223
rect 2927 2216 3093 2224
rect 3147 2216 3293 2224
rect 3336 2226 3344 2296
rect 3707 2296 3893 2304
rect 4267 2296 4453 2304
rect 5316 2304 5324 2316
rect 6796 2324 6804 2333
rect 6647 2316 6804 2324
rect 7927 2316 7953 2324
rect 8047 2316 8093 2324
rect 8433 2324 8447 2333
rect 8433 2320 8733 2324
rect 8436 2316 8733 2320
rect 8947 2316 9053 2324
rect 10767 2316 10913 2324
rect 11107 2316 11153 2324
rect 4467 2296 5324 2304
rect 5347 2296 5513 2304
rect 5667 2296 5753 2304
rect 5807 2296 6133 2304
rect 6187 2296 6353 2304
rect 6627 2296 6953 2304
rect 7267 2296 7293 2304
rect 7307 2296 7333 2304
rect 7467 2296 7633 2304
rect 8027 2296 8173 2304
rect 9187 2296 9453 2304
rect 9507 2296 9573 2304
rect 9587 2296 9733 2304
rect 9987 2296 10253 2304
rect 11287 2296 11333 2304
rect 3427 2276 3513 2284
rect 3527 2276 3593 2284
rect 5047 2276 5173 2284
rect 5727 2276 5773 2284
rect 6667 2276 7093 2284
rect 8027 2276 8053 2284
rect 8707 2276 8793 2284
rect 8987 2276 9013 2284
rect 9767 2276 9833 2284
rect 10347 2276 10373 2284
rect 10447 2276 10493 2284
rect 11227 2276 11253 2284
rect 3367 2256 3473 2264
rect 3607 2257 3653 2265
rect 4267 2256 4433 2264
rect 3816 2244 3824 2254
rect 4456 2256 4493 2264
rect 4456 2244 4464 2256
rect 4727 2257 4792 2265
rect 4827 2256 4933 2264
rect 4987 2257 5013 2265
rect 5196 2256 5233 2264
rect 3747 2236 4464 2244
rect 3487 2216 3613 2224
rect 3707 2215 3793 2223
rect 3847 2215 4093 2223
rect 4287 2215 4353 2223
rect 4447 2215 4473 2223
rect 4527 2215 4673 2223
rect 4807 2216 5073 2224
rect 5196 2226 5204 2256
rect 5287 2256 5393 2264
rect 5447 2256 5493 2264
rect 5827 2257 5893 2265
rect 5947 2256 5993 2264
rect 6187 2257 6213 2265
rect 6507 2256 6533 2264
rect 6947 2256 7073 2264
rect 7927 2257 8133 2265
rect 8827 2256 8953 2264
rect 9207 2256 9364 2264
rect 6967 2237 6993 2245
rect 7547 2236 7753 2244
rect 7767 2236 8124 2244
rect 5456 2216 5573 2224
rect 927 2196 1104 2204
rect 1596 2196 1913 2204
rect 1596 2184 1604 2196
rect 2807 2196 4773 2204
rect 5456 2204 5464 2216
rect 5767 2216 6153 2224
rect 6227 2216 6553 2224
rect 6567 2216 6653 2224
rect 7147 2215 7193 2223
rect 7247 2216 7433 2224
rect 7787 2216 7853 2224
rect 7867 2216 8013 2224
rect 8116 2226 8124 2236
rect 8227 2236 8253 2244
rect 9356 2244 9364 2256
rect 9487 2256 9533 2264
rect 9987 2256 10173 2264
rect 10407 2256 10424 2264
rect 9936 2244 9944 2254
rect 9356 2236 9944 2244
rect 10416 2244 10424 2256
rect 10647 2256 10773 2264
rect 10987 2257 11093 2265
rect 11187 2257 11293 2265
rect 10416 2236 10533 2244
rect 8987 2215 9013 2223
rect 9496 2216 9633 2224
rect 5007 2196 5464 2204
rect 5476 2196 5713 2204
rect 1167 2176 1604 2184
rect 2147 2176 2233 2184
rect 2247 2176 2293 2184
rect 2627 2176 2693 2184
rect 2707 2176 2813 2184
rect 3287 2176 3373 2184
rect 3547 2176 3653 2184
rect 3667 2176 3953 2184
rect 3967 2176 4233 2184
rect 4247 2176 4353 2184
rect 5167 2176 5273 2184
rect 5476 2184 5484 2196
rect 5727 2196 5793 2204
rect 5867 2196 5953 2204
rect 8587 2195 8653 2203
rect 9496 2204 9504 2216
rect 9756 2226 9764 2236
rect 9767 2216 9913 2224
rect 10207 2215 10253 2223
rect 10267 2216 10353 2224
rect 10567 2215 10613 2223
rect 10707 2216 10873 2224
rect 11007 2215 11033 2223
rect 11047 2216 11233 2224
rect 9087 2196 9504 2204
rect 9527 2196 9653 2204
rect 9947 2196 10153 2204
rect 10996 2204 11004 2212
rect 10487 2196 11004 2204
rect 11107 2196 11153 2204
rect 5427 2176 5484 2184
rect 5547 2176 5673 2184
rect 6287 2176 7153 2184
rect 7227 2176 7333 2184
rect 7387 2176 7573 2184
rect 8007 2176 8413 2184
rect 8907 2176 9013 2184
rect 9907 2176 10193 2184
rect 10327 2176 10413 2184
rect 10627 2176 10752 2184
rect 10787 2176 11073 2184
rect 1347 2156 1613 2164
rect 1807 2156 1973 2164
rect 2136 2164 2144 2173
rect 1987 2156 2144 2164
rect 2156 2156 2933 2164
rect 2156 2144 2164 2156
rect 3107 2156 3693 2164
rect 4487 2156 4813 2164
rect 5187 2156 5353 2164
rect 7667 2156 8633 2164
rect 9107 2156 9953 2164
rect 9967 2156 10184 2164
rect 1887 2136 2164 2144
rect 2487 2136 2993 2144
rect 3067 2136 3733 2144
rect 4007 2136 4053 2144
rect 4067 2136 4653 2144
rect 4667 2136 5533 2144
rect 5547 2136 5813 2144
rect 6487 2136 6593 2144
rect 6787 2136 6953 2144
rect 7347 2136 8513 2144
rect 8927 2136 9064 2144
rect 707 2116 973 2124
rect 1876 2116 3213 2124
rect 287 2096 993 2104
rect 1876 2104 1884 2116
rect 3287 2116 3492 2124
rect 3527 2116 3693 2124
rect 4107 2116 4992 2124
rect 5027 2116 5493 2124
rect 8187 2116 8273 2124
rect 8567 2116 8693 2124
rect 9056 2124 9064 2136
rect 9687 2136 9933 2144
rect 10176 2144 10184 2156
rect 10547 2156 10653 2164
rect 10847 2156 10953 2164
rect 11207 2156 11293 2164
rect 10027 2136 10084 2144
rect 10176 2136 10313 2144
rect 9056 2116 9553 2124
rect 9816 2116 9853 2124
rect 1487 2096 1884 2104
rect 1907 2096 3173 2104
rect 3427 2096 3673 2104
rect 3987 2096 4413 2104
rect 5167 2096 5253 2104
rect 5887 2096 6033 2104
rect 6496 2096 7713 2104
rect 6496 2087 6504 2096
rect 8967 2096 9293 2104
rect 9816 2104 9824 2116
rect 10076 2124 10084 2136
rect 10407 2136 10493 2144
rect 10076 2116 10373 2124
rect 9667 2096 9824 2104
rect 10107 2096 10653 2104
rect 207 2076 253 2084
rect 1087 2076 1313 2084
rect 1407 2076 2573 2084
rect 2587 2076 3713 2084
rect 4047 2076 4373 2084
rect 4547 2076 5013 2084
rect 5287 2076 5333 2084
rect 5507 2076 6493 2084
rect 6627 2076 7293 2084
rect 7367 2076 7933 2084
rect 9327 2076 9833 2084
rect 9847 2076 10013 2084
rect 407 2056 1233 2064
rect 2007 2056 2053 2064
rect 2847 2056 2873 2064
rect 3047 2056 3113 2064
rect 3247 2056 3773 2064
rect 4947 2056 5193 2064
rect 5727 2056 6073 2064
rect 6167 2056 6293 2064
rect 6427 2056 6553 2064
rect 6927 2056 7373 2064
rect 7847 2056 8553 2064
rect 8667 2056 9133 2064
rect 9587 2056 9933 2064
rect 627 2036 1173 2044
rect 1327 2036 1853 2044
rect 2167 2036 2273 2044
rect 2807 2036 2953 2044
rect 3227 2036 4633 2044
rect 4787 2036 5293 2044
rect 5447 2036 5732 2044
rect 5767 2036 6033 2044
rect 6047 2036 6453 2044
rect 6467 2036 6733 2044
rect 6747 2036 6813 2044
rect 6827 2036 7393 2044
rect 7407 2036 7673 2044
rect 7716 2036 8573 2044
rect 1307 2016 1493 2024
rect 1827 2016 1853 2024
rect 2307 2016 2413 2024
rect 3907 2016 4233 2024
rect 5607 2016 5653 2024
rect 5667 2016 5953 2024
rect 5967 2016 6013 2024
rect 6907 2016 7013 2024
rect 7716 2024 7724 2036
rect 8947 2036 9113 2044
rect 9467 2036 9593 2044
rect 7427 2016 7724 2024
rect 8087 2016 8133 2024
rect 8227 2016 8493 2024
rect 8647 2016 8673 2024
rect 8827 2016 9313 2024
rect 9727 2016 10673 2024
rect 1607 1996 1893 2004
rect 2007 1996 2284 2004
rect 947 1976 1473 1984
rect 2276 1984 2284 1996
rect 2467 1996 3033 2004
rect 3087 1996 3153 2004
rect 3267 1996 3473 2004
rect 3587 1996 4433 2004
rect 4447 1996 4673 2004
rect 4727 1996 4953 2004
rect 5787 1996 5933 2004
rect 6087 1996 6113 2004
rect 6187 1996 6473 2004
rect 7187 1996 7253 2004
rect 7967 1996 8093 2004
rect 8107 1996 8233 2004
rect 8587 1996 8953 2004
rect 9127 1996 9253 2004
rect 9407 1996 9533 2004
rect 9627 1996 9833 2004
rect 10347 1996 10633 2004
rect 11087 1996 11253 2004
rect 2276 1976 2333 1984
rect 2347 1976 2373 1984
rect 6767 1976 6833 1984
rect 7007 1976 7293 1984
rect 8067 1976 8213 1984
rect 8567 1976 9193 1984
rect 9207 1976 9953 1984
rect 667 1956 713 1964
rect 727 1957 793 1965
rect 847 1957 873 1965
rect 1027 1957 1113 1965
rect 1167 1957 1293 1965
rect 1547 1957 1792 1965
rect 1827 1957 1953 1965
rect 2067 1957 2193 1965
rect 2207 1956 2253 1964
rect 2427 1956 2593 1964
rect 2647 1956 2833 1964
rect 3267 1957 3313 1965
rect 1476 1936 1873 1944
rect 187 1915 253 1923
rect 427 1915 493 1923
rect 507 1916 593 1924
rect 647 1915 693 1923
rect 767 1916 813 1924
rect 1067 1915 1153 1923
rect 1476 1926 1484 1936
rect 1207 1916 1273 1924
rect 2867 1916 2953 1924
rect 3096 1924 3104 1954
rect 3467 1956 3673 1964
rect 3827 1957 3873 1965
rect 3927 1956 3993 1964
rect 4187 1957 4273 1965
rect 4807 1957 4893 1965
rect 5007 1956 5152 1964
rect 5187 1964 5200 1967
rect 5187 1953 5204 1964
rect 3556 1936 3693 1944
rect 2967 1916 3104 1924
rect 3247 1916 3333 1924
rect 3387 1916 3433 1924
rect 3556 1926 3564 1936
rect 5196 1946 5204 1953
rect 5276 1947 5284 1973
rect 5596 1956 5633 1964
rect 5596 1944 5604 1956
rect 5807 1956 5893 1964
rect 6087 1956 6213 1964
rect 6527 1957 6573 1965
rect 6887 1957 6953 1965
rect 7087 1956 7213 1964
rect 8307 1956 8453 1964
rect 8687 1957 8753 1965
rect 8847 1957 8913 1965
rect 8967 1957 9033 1965
rect 9107 1957 9153 1965
rect 9627 1957 9673 1965
rect 9807 1956 9893 1964
rect 10056 1956 10073 1964
rect 5567 1936 5604 1944
rect 5627 1936 5733 1944
rect 7507 1936 8153 1944
rect 10056 1944 10064 1956
rect 10387 1956 10413 1964
rect 10427 1957 10473 1965
rect 10527 1957 10593 1965
rect 10787 1956 10993 1964
rect 11007 1956 11173 1964
rect 11196 1956 11213 1964
rect 9507 1936 10064 1944
rect 3847 1915 3913 1923
rect 4027 1916 4173 1924
rect 4707 1916 4793 1924
rect 4847 1916 4873 1924
rect 5907 1915 6013 1923
rect 6067 1916 6173 1924
rect 6227 1915 6253 1923
rect 6307 1915 6373 1923
rect 6387 1916 6593 1924
rect 6687 1915 6713 1923
rect 6767 1916 6873 1924
rect 7147 1916 7193 1924
rect 7407 1916 7913 1924
rect 8247 1915 8273 1923
rect 8487 1916 8653 1924
rect 8907 1916 8933 1924
rect 8947 1920 8984 1924
rect 8947 1916 8987 1920
rect 8973 1907 8987 1916
rect 9027 1916 9133 1924
rect 9387 1915 9473 1923
rect 9687 1916 9813 1924
rect 9907 1916 10113 1924
rect 10127 1916 10153 1924
rect 10407 1916 10453 1924
rect 10687 1915 10713 1923
rect 10736 1924 10744 1954
rect 11196 1944 11204 1956
rect 11156 1940 11204 1944
rect 11153 1936 11204 1940
rect 11153 1927 11167 1936
rect 10736 1916 10793 1924
rect 10967 1915 11013 1923
rect 1707 1896 1993 1904
rect 2107 1896 2133 1904
rect 2407 1896 2813 1904
rect 4487 1896 4684 1904
rect 387 1876 533 1884
rect 547 1876 733 1884
rect 1127 1876 1513 1884
rect 1947 1876 2013 1884
rect 2187 1876 2553 1884
rect 2667 1876 3073 1884
rect 3207 1876 3413 1884
rect 3567 1876 3892 1884
rect 3927 1876 3993 1884
rect 4007 1876 4213 1884
rect 4507 1876 4533 1884
rect 4676 1884 4684 1896
rect 5307 1896 5913 1904
rect 7596 1896 7653 1904
rect 4676 1876 4913 1884
rect 5147 1876 5213 1884
rect 5967 1876 6093 1884
rect 6567 1876 6913 1884
rect 7596 1884 7604 1896
rect 7947 1896 8033 1904
rect 8047 1896 8113 1904
rect 8707 1896 8733 1904
rect 9047 1896 9173 1904
rect 9187 1896 9233 1904
rect 9947 1896 10053 1904
rect 10367 1896 10533 1904
rect 10867 1896 11113 1904
rect 7147 1876 7604 1884
rect 7616 1876 8553 1884
rect 1107 1856 1133 1864
rect 2287 1856 2453 1864
rect 2476 1856 3493 1864
rect 827 1836 1813 1844
rect 2476 1844 2484 1856
rect 3507 1856 4433 1864
rect 4947 1856 5253 1864
rect 5267 1856 5713 1864
rect 5767 1856 6433 1864
rect 7616 1864 7624 1876
rect 8867 1876 9553 1884
rect 9627 1876 10093 1884
rect 10147 1876 10293 1884
rect 10507 1876 10613 1884
rect 10667 1876 10753 1884
rect 11147 1876 11193 1884
rect 7267 1856 7624 1864
rect 8127 1856 8293 1864
rect 8307 1856 8513 1864
rect 9147 1856 9293 1864
rect 9307 1856 9433 1864
rect 9887 1856 10033 1864
rect 10427 1856 10933 1864
rect 11127 1856 11233 1864
rect 2187 1836 2484 1844
rect 2507 1836 3013 1844
rect 3607 1836 4473 1844
rect 4607 1836 4913 1844
rect 5067 1836 5193 1844
rect 5387 1836 5633 1844
rect 6847 1836 6973 1844
rect 7127 1836 7993 1844
rect 8767 1836 9533 1844
rect 9547 1836 9653 1844
rect 9967 1836 10013 1844
rect 10747 1836 10813 1844
rect 1007 1816 1453 1824
rect 2027 1816 2613 1824
rect 3127 1816 3553 1824
rect 3747 1816 4173 1824
rect 4347 1816 4453 1824
rect 4527 1816 4613 1824
rect 5867 1816 6013 1824
rect 6067 1816 6213 1824
rect 6347 1816 6493 1824
rect 7507 1816 7733 1824
rect 8756 1824 8764 1833
rect 7867 1816 8764 1824
rect 9607 1816 9773 1824
rect 10427 1816 10553 1824
rect 627 1796 733 1804
rect 1147 1796 1833 1804
rect 1847 1796 1913 1804
rect 2147 1796 2212 1804
rect 2247 1796 2313 1804
rect 2467 1796 2773 1804
rect 3087 1796 3293 1804
rect 3907 1796 4993 1804
rect 5947 1796 5993 1804
rect 7813 1804 7827 1813
rect 7267 1800 7827 1804
rect 7267 1796 7824 1800
rect 7836 1796 7973 1804
rect 207 1776 293 1784
rect 307 1776 813 1784
rect 1387 1776 1413 1784
rect 1787 1776 2013 1784
rect 2027 1776 2053 1784
rect 2067 1776 2713 1784
rect 2727 1776 2893 1784
rect 2907 1776 2933 1784
rect 2947 1776 3393 1784
rect 3407 1776 3553 1784
rect 3687 1776 4473 1784
rect 5087 1776 5293 1784
rect 5607 1776 5733 1784
rect 6027 1776 6133 1784
rect 6667 1776 7193 1784
rect 7836 1784 7844 1796
rect 9267 1804 9280 1807
rect 9267 1800 9284 1804
rect 9267 1793 9287 1800
rect 9327 1796 9913 1804
rect 10107 1796 10273 1804
rect 10927 1796 11213 1804
rect 9273 1787 9287 1793
rect 7587 1776 7844 1784
rect 8587 1776 9213 1784
rect 9347 1776 9713 1784
rect 10467 1776 10613 1784
rect 10967 1776 11113 1784
rect 847 1756 973 1764
rect 1047 1756 1793 1764
rect 3787 1756 3933 1764
rect 4547 1756 4573 1764
rect 4587 1756 4933 1764
rect 5107 1756 5153 1764
rect 5247 1756 5273 1764
rect 5347 1756 5533 1764
rect 5547 1756 5573 1764
rect 5740 1764 5753 1767
rect 5736 1753 5753 1764
rect 5927 1756 5973 1764
rect 6707 1756 6813 1764
rect 7027 1756 7253 1764
rect 7727 1756 8053 1764
rect 9180 1764 9193 1767
rect 8667 1756 9193 1764
rect 9176 1753 9193 1756
rect 9956 1756 10253 1764
rect 427 1737 513 1745
rect 667 1736 773 1744
rect 1267 1736 1413 1744
rect 1467 1737 1713 1745
rect 1727 1736 1773 1744
rect 1887 1736 2053 1744
rect 2147 1737 2233 1745
rect 2327 1737 2353 1745
rect 2407 1736 2544 1744
rect 2536 1724 2544 1736
rect 2687 1737 2733 1745
rect 2596 1724 2604 1734
rect 2747 1737 2853 1745
rect 2927 1737 3033 1745
rect 3187 1737 3253 1745
rect 3267 1736 3413 1744
rect 3540 1744 3553 1747
rect 3536 1733 3553 1744
rect 3767 1737 3813 1745
rect 3907 1736 3953 1744
rect 4227 1737 4253 1745
rect 4267 1736 4393 1744
rect 4736 1740 4813 1744
rect 4733 1736 4813 1740
rect 2536 1716 2653 1724
rect 227 1696 393 1704
rect 407 1696 633 1704
rect 887 1696 1013 1704
rect 1027 1695 1133 1703
rect 1547 1695 1673 1703
rect 2387 1695 2453 1703
rect 2627 1696 2793 1704
rect 3287 1696 3373 1704
rect 3536 1706 3544 1733
rect 4733 1727 4747 1736
rect 4887 1736 4933 1744
rect 5187 1737 5513 1745
rect 5736 1744 5744 1753
rect 9176 1748 9184 1753
rect 5527 1736 5744 1744
rect 5787 1737 5873 1745
rect 4456 1720 4553 1724
rect 4453 1716 4553 1720
rect 4453 1707 4467 1716
rect 4867 1716 4904 1724
rect 3587 1695 3933 1703
rect 4896 1687 4904 1716
rect 5116 1724 5124 1734
rect 5027 1716 5124 1724
rect 5227 1716 5493 1724
rect 5876 1724 5884 1734
rect 6587 1736 7313 1744
rect 7407 1737 7473 1745
rect 7527 1737 7613 1745
rect 8227 1737 8253 1745
rect 8507 1736 8593 1744
rect 5876 1716 6024 1724
rect 5107 1696 5193 1704
rect 6016 1706 6024 1716
rect 6307 1715 6473 1723
rect 7653 1724 7667 1733
rect 7653 1720 7813 1724
rect 7656 1716 7813 1720
rect 8216 1724 8224 1734
rect 8747 1736 8793 1744
rect 8907 1737 8933 1745
rect 9227 1736 9353 1744
rect 9407 1737 9533 1745
rect 9727 1737 9893 1745
rect 9956 1744 9964 1756
rect 10347 1756 10393 1764
rect 9907 1736 9964 1744
rect 9987 1737 10113 1745
rect 10507 1736 10593 1744
rect 10607 1736 10673 1744
rect 10787 1736 10913 1744
rect 10927 1737 10993 1745
rect 11067 1737 11253 1745
rect 8216 1716 8524 1724
rect 5327 1695 5373 1703
rect 5807 1695 5853 1703
rect 6567 1696 6633 1704
rect 7007 1696 7113 1704
rect 7127 1695 7433 1703
rect 8516 1706 8524 1716
rect 7487 1696 7593 1704
rect 8867 1696 8953 1704
rect 9167 1696 9373 1704
rect 9567 1695 9593 1703
rect 9787 1696 10053 1704
rect 10307 1696 10413 1704
rect 10687 1695 10713 1703
rect 11087 1695 11133 1703
rect 11147 1695 11193 1703
rect 187 1676 253 1684
rect 267 1676 473 1684
rect 1507 1676 1753 1684
rect 1767 1676 1893 1684
rect 2887 1676 2933 1684
rect 2947 1676 3033 1684
rect 3107 1676 3153 1684
rect 3167 1676 3493 1684
rect 5407 1676 5693 1684
rect 607 1656 1093 1664
rect 1847 1656 1893 1664
rect 1907 1656 2293 1664
rect 2667 1656 3073 1664
rect 3547 1656 3653 1664
rect 4713 1664 4727 1673
rect 6107 1675 6453 1683
rect 8147 1676 8413 1684
rect 8767 1676 8813 1684
rect 9107 1676 9153 1684
rect 10887 1676 11013 1684
rect 4713 1660 4833 1664
rect 4716 1656 4833 1660
rect 5067 1656 5653 1664
rect 7567 1656 8573 1664
rect 9487 1656 9553 1664
rect 9867 1656 10213 1664
rect 10287 1656 10473 1664
rect 10767 1656 10853 1664
rect 11167 1656 11233 1664
rect 647 1636 1053 1644
rect 1247 1636 1273 1644
rect 1787 1636 2513 1644
rect 2847 1636 3873 1644
rect 3927 1636 5273 1644
rect 5987 1636 6513 1644
rect 6687 1636 6913 1644
rect 6927 1636 7333 1644
rect 7587 1636 7653 1644
rect 8596 1636 8713 1644
rect 947 1616 1273 1624
rect 1647 1616 2653 1624
rect 3067 1616 3504 1624
rect 427 1596 713 1604
rect 727 1596 813 1604
rect 1947 1596 2973 1604
rect 3496 1604 3504 1616
rect 3667 1616 3704 1624
rect 3496 1596 3673 1604
rect 3696 1604 3704 1616
rect 3947 1616 4693 1624
rect 4887 1616 5053 1624
rect 5507 1616 5993 1624
rect 6927 1616 7053 1624
rect 8167 1616 8193 1624
rect 8596 1624 8604 1636
rect 9007 1636 9173 1644
rect 10747 1636 11033 1644
rect 8207 1616 8604 1624
rect 8767 1616 8793 1624
rect 9387 1616 9813 1624
rect 9827 1616 10213 1624
rect 10527 1616 10833 1624
rect 11227 1616 11293 1624
rect 3696 1596 4193 1604
rect 5147 1596 6573 1604
rect 7167 1596 7553 1604
rect 8227 1596 8613 1604
rect 9287 1596 9373 1604
rect 9427 1596 9633 1604
rect 10727 1596 10813 1604
rect 1587 1576 3093 1584
rect 3167 1576 3653 1584
rect 3787 1576 3972 1584
rect 4007 1576 4153 1584
rect 4667 1576 4832 1584
rect 4867 1576 4933 1584
rect 5007 1576 6033 1584
rect 8807 1576 9853 1584
rect 11107 1576 11253 1584
rect 1427 1556 1553 1564
rect 1916 1556 2033 1564
rect 1916 1544 1924 1556
rect 2047 1556 2113 1564
rect 2767 1556 2833 1564
rect 3427 1556 3473 1564
rect 3587 1556 3713 1564
rect 3847 1556 4784 1564
rect 4776 1547 4784 1556
rect 4807 1556 4973 1564
rect 4996 1556 5393 1564
rect 987 1536 1924 1544
rect 2527 1536 3084 1544
rect 787 1516 1933 1524
rect 3076 1524 3084 1536
rect 3687 1536 3772 1544
rect 3807 1536 4073 1544
rect 4167 1536 4613 1544
rect 4996 1544 5004 1556
rect 6947 1556 7273 1564
rect 7387 1556 7793 1564
rect 8287 1556 8633 1564
rect 8647 1556 9133 1564
rect 9147 1556 9453 1564
rect 9647 1556 9833 1564
rect 9847 1556 10093 1564
rect 10107 1556 11073 1564
rect 4787 1536 5004 1544
rect 5687 1536 6753 1544
rect 8747 1536 8892 1544
rect 8927 1536 9093 1544
rect 9167 1536 9593 1544
rect 9987 1536 10073 1544
rect 10487 1536 10633 1544
rect 3076 1516 3553 1524
rect 3887 1516 4473 1524
rect 4707 1516 5173 1524
rect 6547 1516 7253 1524
rect 7307 1516 10373 1524
rect 207 1496 1353 1504
rect 1367 1496 1913 1504
rect 1987 1496 2313 1504
rect 2907 1496 3953 1504
rect 4607 1496 4813 1504
rect 4947 1496 5013 1504
rect 5247 1496 5293 1504
rect 5567 1496 5893 1504
rect 6007 1496 6333 1504
rect 6487 1496 6993 1504
rect 7527 1496 7873 1504
rect 9367 1496 9873 1504
rect 10167 1496 10293 1504
rect 10407 1496 10533 1504
rect 1507 1476 1593 1484
rect 1707 1476 1833 1484
rect 2547 1476 2993 1484
rect 3427 1476 4133 1484
rect 4267 1476 4873 1484
rect 4927 1476 5372 1484
rect 5407 1476 6293 1484
rect 6467 1476 7573 1484
rect 7876 1484 7884 1493
rect 7876 1476 8113 1484
rect 8247 1476 8792 1484
rect 8827 1476 8893 1484
rect 9247 1476 9324 1484
rect 747 1456 853 1464
rect 867 1456 1033 1464
rect 1516 1456 1584 1464
rect 787 1437 813 1445
rect 1087 1437 1153 1445
rect 1227 1436 1313 1444
rect 1516 1444 1524 1456
rect 1327 1436 1524 1444
rect 1576 1444 1584 1456
rect 1767 1456 2153 1464
rect 3227 1456 3253 1464
rect 3567 1456 3773 1464
rect 3827 1456 4013 1464
rect 4227 1456 4573 1464
rect 4627 1456 4733 1464
rect 4747 1456 4793 1464
rect 5247 1456 5673 1464
rect 5727 1456 5892 1464
rect 5927 1456 5953 1464
rect 6807 1456 6853 1464
rect 6907 1456 7033 1464
rect 7047 1456 7153 1464
rect 7267 1456 7493 1464
rect 8567 1456 8673 1464
rect 8847 1456 8913 1464
rect 9316 1464 9324 1476
rect 9647 1476 9733 1484
rect 9947 1476 10133 1484
rect 10347 1476 10593 1484
rect 9316 1456 9493 1464
rect 9507 1456 10153 1464
rect 10207 1456 10233 1464
rect 10587 1456 10673 1464
rect 1576 1436 1813 1444
rect 2367 1437 2413 1445
rect 2427 1437 2433 1445
rect 2567 1436 2753 1444
rect 3047 1436 3284 1444
rect 1547 1416 1973 1424
rect 107 1395 213 1403
rect 227 1396 433 1404
rect 447 1396 613 1404
rect 1067 1396 1213 1404
rect 1916 1406 1924 1416
rect 1227 1396 1253 1404
rect 1347 1395 1473 1403
rect 1567 1395 1673 1403
rect 1747 1395 1873 1403
rect 2107 1395 2213 1403
rect 2787 1396 2893 1404
rect 3027 1396 3173 1404
rect 3276 1406 3284 1436
rect 3607 1436 3733 1444
rect 3867 1436 3993 1444
rect 4107 1436 4153 1444
rect 4727 1437 4813 1445
rect 5047 1436 5073 1444
rect 5467 1436 5533 1444
rect 5787 1436 6093 1444
rect 6307 1437 7073 1445
rect 7147 1436 7233 1444
rect 7307 1436 7413 1444
rect 7427 1436 7613 1444
rect 7667 1437 7753 1445
rect 7807 1437 7833 1445
rect 8027 1436 8073 1444
rect 8127 1436 8313 1444
rect 8987 1437 9033 1445
rect 9127 1436 9253 1444
rect 9267 1437 9293 1445
rect 9427 1437 9453 1445
rect 9607 1436 9693 1444
rect 9747 1437 9793 1445
rect 10407 1436 10453 1444
rect 10467 1436 10564 1444
rect 3407 1416 3724 1424
rect 3467 1395 3593 1403
rect 3716 1404 3724 1416
rect 6756 1416 6953 1424
rect 3716 1396 3753 1404
rect 3887 1395 3933 1403
rect 3987 1396 4173 1404
rect 4447 1396 5113 1404
rect 5387 1395 5433 1403
rect 5627 1396 5653 1404
rect 5707 1395 5773 1403
rect 5927 1395 5993 1403
rect 6127 1396 6313 1404
rect 6367 1396 6433 1404
rect 6447 1396 6733 1404
rect 6756 1404 6764 1416
rect 8667 1416 8913 1424
rect 10556 1424 10564 1436
rect 10787 1437 10873 1445
rect 10636 1424 10644 1434
rect 10556 1416 10644 1424
rect 6747 1396 6764 1404
rect 7507 1396 7633 1404
rect 7907 1395 7953 1403
rect 7967 1396 8133 1404
rect 8287 1395 8613 1403
rect 8687 1396 8853 1404
rect 9067 1396 9153 1404
rect 9227 1396 9473 1404
rect 3367 1376 3593 1384
rect 4407 1376 5133 1384
rect 6827 1376 7013 1384
rect 7027 1376 7433 1384
rect 8147 1376 8333 1384
rect 9216 1384 9224 1393
rect 9587 1396 9673 1404
rect 9727 1395 9813 1403
rect 9867 1395 9913 1403
rect 9967 1396 10013 1404
rect 10267 1395 10373 1403
rect 10767 1396 10813 1404
rect 9087 1376 9224 1384
rect 10407 1376 10513 1384
rect 10887 1376 10933 1384
rect 11227 1376 11273 1384
rect 207 1356 333 1364
rect 427 1356 493 1364
rect 967 1356 1053 1364
rect 1287 1356 1393 1364
rect 1407 1356 2053 1364
rect 2727 1356 2833 1364
rect 2847 1356 3693 1364
rect 4396 1364 4404 1373
rect 4027 1356 4404 1364
rect 4416 1356 5073 1364
rect 1647 1336 1733 1344
rect 1807 1336 2533 1344
rect 2547 1336 2673 1344
rect 3187 1336 3633 1344
rect 4416 1344 4424 1356
rect 5127 1356 6773 1364
rect 6867 1356 7053 1364
rect 8027 1356 8652 1364
rect 8687 1356 8953 1364
rect 8967 1356 9013 1364
rect 9027 1356 9253 1364
rect 9427 1356 9473 1364
rect 9767 1356 10073 1364
rect 10727 1356 10813 1364
rect 3887 1336 4424 1344
rect 4607 1336 5553 1344
rect 7167 1336 7233 1344
rect 7247 1336 7313 1344
rect 8147 1336 8813 1344
rect 8827 1336 8972 1344
rect 9007 1336 9073 1344
rect 9147 1336 9653 1344
rect 9707 1336 10253 1344
rect 10587 1336 10853 1344
rect 10907 1336 10953 1344
rect 407 1316 513 1324
rect 847 1316 1572 1324
rect 1607 1316 2133 1324
rect 3027 1316 4124 1324
rect 1727 1296 1993 1304
rect 2147 1296 2833 1304
rect 3207 1296 3573 1304
rect 3687 1296 3833 1304
rect 4116 1304 4124 1316
rect 4147 1316 4233 1324
rect 4247 1316 4433 1324
rect 4827 1316 4853 1324
rect 5087 1316 6133 1324
rect 6147 1316 7133 1324
rect 7187 1316 7853 1324
rect 9427 1316 9613 1324
rect 4116 1296 4273 1304
rect 4547 1296 4993 1304
rect 5347 1296 5473 1304
rect 5907 1296 6073 1304
rect 6307 1296 6593 1304
rect 6647 1296 6773 1304
rect 9147 1296 9173 1304
rect 9647 1296 9713 1304
rect 10207 1296 10493 1304
rect 10747 1296 11073 1304
rect 11087 1296 11193 1304
rect 87 1276 833 1284
rect 1527 1276 2713 1284
rect 3007 1276 3133 1284
rect 4627 1276 4793 1284
rect 4867 1276 4893 1284
rect 5187 1276 5673 1284
rect 5687 1276 6193 1284
rect 6207 1276 6473 1284
rect 8067 1276 8093 1284
rect 8107 1276 8273 1284
rect 8407 1276 8713 1284
rect 8927 1276 9013 1284
rect 1467 1256 1633 1264
rect 1687 1256 1893 1264
rect 2447 1256 2733 1264
rect 3707 1256 3853 1264
rect 3907 1256 4253 1264
rect 4747 1256 4773 1264
rect 5027 1256 6213 1264
rect 7107 1256 7233 1264
rect 7247 1256 7253 1264
rect 7267 1256 7813 1264
rect 8767 1256 8833 1264
rect 9067 1256 9833 1264
rect 9847 1256 9913 1264
rect 9987 1256 10093 1264
rect 4527 1236 4913 1244
rect 5007 1236 5253 1244
rect 5487 1236 6093 1244
rect 6367 1236 6484 1244
rect 6476 1228 6484 1236
rect 7007 1236 7053 1244
rect 8547 1236 8613 1244
rect 8727 1236 8973 1244
rect 9387 1236 9573 1244
rect 10307 1236 10413 1244
rect 10547 1236 10633 1244
rect 567 1216 613 1224
rect 627 1217 653 1225
rect 667 1217 673 1225
rect 847 1216 1653 1224
rect 1767 1216 1793 1224
rect 1867 1217 1933 1225
rect 1987 1217 2093 1225
rect 2207 1217 2233 1225
rect 2407 1216 2544 1224
rect 2536 1204 2544 1216
rect 2567 1217 2593 1225
rect 2647 1216 2713 1224
rect 2727 1216 2973 1224
rect 2987 1217 3053 1225
rect 3107 1216 3253 1224
rect 3327 1216 3393 1224
rect 3507 1216 3553 1224
rect 3607 1217 3653 1225
rect 3767 1216 3793 1224
rect 3860 1224 3873 1227
rect 3856 1213 3873 1224
rect 4067 1216 4133 1224
rect 4407 1216 4453 1224
rect 4567 1216 4793 1224
rect 5447 1216 5493 1224
rect 5547 1217 5633 1225
rect 6487 1217 6533 1225
rect 6587 1217 6613 1225
rect 6667 1216 7193 1224
rect 7207 1217 7273 1225
rect 7667 1216 7953 1224
rect 2536 1196 3013 1204
rect 227 1176 393 1184
rect 647 1176 773 1184
rect 787 1176 813 1184
rect 1747 1175 1833 1183
rect 1907 1175 2413 1183
rect 2427 1176 2473 1184
rect 3047 1175 3073 1183
rect 3127 1175 3193 1183
rect 3267 1175 3293 1183
rect 3487 1175 3533 1183
rect 3587 1175 3613 1183
rect 3856 1186 3864 1213
rect 3927 1196 4144 1204
rect 3667 1176 3773 1184
rect 3787 1176 3824 1184
rect 1067 1156 1113 1164
rect 1607 1156 1693 1164
rect 2067 1156 2553 1164
rect 2567 1156 2913 1164
rect 3816 1164 3824 1176
rect 4087 1175 4113 1183
rect 4136 1184 4144 1196
rect 4516 1204 4524 1213
rect 4347 1196 4524 1204
rect 5087 1196 5333 1204
rect 7416 1204 7424 1214
rect 8007 1216 8033 1224
rect 8047 1217 8093 1225
rect 8507 1217 8673 1225
rect 8727 1216 8853 1224
rect 9167 1217 9213 1225
rect 9307 1217 9613 1225
rect 9667 1216 9833 1224
rect 9887 1217 9953 1225
rect 10187 1217 10273 1225
rect 10527 1216 10964 1224
rect 5527 1196 6144 1204
rect 7416 1196 7664 1204
rect 4136 1176 4693 1184
rect 4747 1175 4773 1183
rect 4887 1175 5373 1183
rect 5427 1175 5473 1183
rect 5667 1176 5753 1184
rect 5967 1175 6113 1183
rect 6136 1184 6144 1196
rect 6136 1176 6653 1184
rect 6807 1175 6833 1183
rect 7287 1176 7433 1184
rect 7507 1175 7633 1183
rect 7656 1184 7664 1196
rect 7656 1176 7673 1184
rect 7687 1175 8013 1183
rect 8247 1176 8293 1184
rect 8527 1175 8653 1183
rect 8867 1176 9193 1184
rect 9207 1176 9233 1184
rect 9347 1175 9393 1183
rect 9867 1176 10073 1184
rect 10096 1184 10104 1214
rect 10956 1204 10964 1216
rect 10987 1217 11032 1225
rect 11067 1216 11233 1224
rect 10956 1196 11184 1204
rect 10096 1176 10133 1184
rect 10227 1175 10293 1183
rect 10427 1175 10713 1183
rect 10827 1176 10933 1184
rect 11007 1175 11053 1183
rect 11176 1186 11184 1196
rect 3816 1156 3913 1164
rect 3967 1156 4553 1164
rect 4807 1156 5513 1164
rect 6267 1156 6553 1164
rect 7087 1156 7513 1164
rect 10347 1156 10893 1164
rect 10907 1156 11053 1164
rect 1207 1136 1273 1144
rect 1967 1136 2113 1144
rect 2227 1136 3873 1144
rect 4067 1136 4753 1144
rect 4767 1136 6093 1144
rect 6227 1136 6504 1144
rect 1627 1116 2173 1124
rect 2987 1116 3453 1124
rect 3827 1116 4033 1124
rect 4567 1116 4813 1124
rect 4827 1116 5073 1124
rect 5207 1116 5713 1124
rect 5856 1120 6133 1124
rect 5853 1116 6133 1120
rect 5853 1107 5867 1116
rect 6496 1124 6504 1136
rect 6767 1136 6933 1144
rect 8747 1136 8773 1144
rect 8867 1136 9293 1144
rect 9647 1136 10073 1144
rect 10367 1136 10653 1144
rect 10747 1136 10793 1144
rect 6496 1116 6973 1124
rect 6987 1116 8573 1124
rect 9407 1116 10173 1124
rect 10267 1116 10533 1124
rect 11227 1116 11273 1124
rect 3476 1096 3824 1104
rect 1827 1076 2213 1084
rect 3476 1084 3484 1096
rect 3347 1076 3484 1084
rect 3816 1084 3824 1096
rect 3947 1096 5813 1104
rect 6167 1096 6333 1104
rect 6487 1096 8133 1104
rect 9947 1096 10113 1104
rect 10127 1096 10493 1104
rect 3816 1076 4593 1084
rect 4667 1076 4713 1084
rect 5987 1076 6133 1084
rect 6627 1076 7013 1084
rect 7027 1076 7173 1084
rect 7227 1076 7553 1084
rect 9447 1076 9593 1084
rect 10307 1076 10413 1084
rect 10427 1076 10473 1084
rect 1687 1056 2993 1064
rect 3007 1056 3033 1064
rect 3247 1056 3693 1064
rect 3887 1056 4553 1064
rect 4947 1056 5933 1064
rect 6347 1056 7773 1064
rect 8527 1056 8853 1064
rect 8907 1056 9733 1064
rect 10147 1056 10613 1064
rect 1907 1036 2273 1044
rect 2287 1036 2593 1044
rect 3507 1036 3613 1044
rect 3787 1036 4353 1044
rect 4847 1036 5333 1044
rect 6067 1036 7453 1044
rect 8707 1036 8833 1044
rect 9247 1036 9473 1044
rect 9487 1036 9933 1044
rect 1467 1016 1813 1024
rect 1867 1016 3033 1024
rect 3047 1016 4573 1024
rect 4707 1016 5113 1024
rect 6867 1016 7293 1024
rect 7827 1016 8373 1024
rect 8567 1016 8993 1024
rect 9187 1016 9973 1024
rect 887 996 1233 1004
rect 1247 996 1293 1004
rect 1367 996 1893 1004
rect 2127 996 2852 1004
rect 2887 996 3813 1004
rect 4867 996 4893 1004
rect 5187 996 5572 1004
rect 5607 996 5613 1004
rect 5627 996 5973 1004
rect 7887 996 8473 1004
rect 8807 996 9113 1004
rect 9507 996 9533 1004
rect 9547 996 9653 1004
rect 9867 996 10053 1004
rect 10067 996 10133 1004
rect 10187 996 10913 1004
rect 2616 976 5513 984
rect 2616 967 2624 976
rect 6127 976 6613 984
rect 7707 976 7793 984
rect 7807 976 8713 984
rect 8727 976 9273 984
rect 9287 976 10213 984
rect 10416 976 10593 984
rect 927 956 1073 964
rect 1087 956 1193 964
rect 2247 956 2353 964
rect 2367 956 2613 964
rect 3847 956 4213 964
rect 4267 956 4893 964
rect 5376 956 5913 964
rect 5376 947 5384 956
rect 6047 956 6753 964
rect 7227 956 7293 964
rect 7907 956 8033 964
rect 8147 956 8213 964
rect 8227 956 8453 964
rect 10416 964 10424 976
rect 10867 976 11293 984
rect 9927 956 10424 964
rect 10467 956 10553 964
rect 147 936 173 944
rect 1427 936 1713 944
rect 3087 936 3233 944
rect 3547 936 3673 944
rect 4507 936 4833 944
rect 5167 936 5373 944
rect 6287 936 6373 944
rect 7007 936 7053 944
rect 7927 936 7953 944
rect 8847 936 9513 944
rect 9607 936 9853 944
rect 247 917 373 925
rect 427 917 433 925
rect 447 917 453 925
rect 607 916 793 924
rect 947 917 973 925
rect 1027 917 1153 925
rect 1167 916 1253 924
rect 1347 917 1453 925
rect 1727 917 1793 925
rect 1847 917 1893 925
rect 1947 916 2133 924
rect 187 876 233 884
rect 407 876 513 884
rect 527 876 573 884
rect 1227 876 1353 884
rect 1487 876 1573 884
rect 1587 875 1653 883
rect 1707 876 1832 884
rect 1867 876 1913 884
rect 2167 875 2253 883
rect 2396 884 2404 914
rect 2447 916 2573 924
rect 2587 916 2733 924
rect 2747 916 2813 924
rect 2827 916 3113 924
rect 3287 917 3393 925
rect 3407 916 3453 924
rect 3587 917 3733 925
rect 4007 916 4153 924
rect 4387 916 4433 924
rect 4627 924 4640 927
rect 4627 913 4644 924
rect 4827 917 4853 925
rect 4876 916 5073 924
rect 2396 876 2593 884
rect 2647 875 2713 883
rect 2727 876 2793 884
rect 2847 876 3373 884
rect 3467 875 3513 883
rect 3707 875 3753 883
rect 3807 876 3953 884
rect 4636 886 4644 913
rect 4876 904 4884 916
rect 5113 924 5127 933
rect 5113 920 5593 924
rect 5116 916 5593 920
rect 5787 916 5873 924
rect 5887 916 6013 924
rect 6267 917 6353 925
rect 6547 917 6593 925
rect 6807 916 7213 924
rect 7547 916 7873 924
rect 8607 917 8652 925
rect 8687 917 8833 925
rect 4747 896 4884 904
rect 8336 904 8344 914
rect 8967 916 9093 924
rect 9447 916 9793 924
rect 9967 916 10093 924
rect 10107 917 10133 925
rect 10347 917 10473 925
rect 6107 896 6224 904
rect 8336 896 8933 904
rect 4027 875 4053 883
rect 4407 875 4453 883
rect 4687 875 4753 883
rect 5107 876 5353 884
rect 5527 875 5993 883
rect 6047 875 6193 883
rect 6216 884 6224 896
rect 9456 896 9493 904
rect 6216 876 6273 884
rect 6447 875 6473 883
rect 6787 875 6853 883
rect 7087 876 7233 884
rect 7487 875 7533 883
rect 7687 876 7813 884
rect 7967 876 8113 884
rect 8167 876 8353 884
rect 8487 876 8573 884
rect 8587 876 8733 884
rect 9207 876 9353 884
rect 9456 884 9464 896
rect 10496 886 10504 933
rect 10527 916 10833 924
rect 10947 916 11153 924
rect 9427 876 9464 884
rect 9607 875 9633 883
rect 9747 875 9833 883
rect 9887 875 9913 883
rect 10087 876 10273 884
rect 627 856 693 864
rect 707 856 973 864
rect 2367 856 2433 864
rect 6436 864 6444 872
rect 6327 856 6444 864
rect 6567 856 6693 864
rect 7987 856 8313 864
rect 8627 856 8813 864
rect 9107 856 9213 864
rect 9227 856 9473 864
rect 11027 856 11153 864
rect 1067 836 1233 844
rect 1276 836 1473 844
rect 1276 824 1284 836
rect 1747 836 3893 844
rect 4167 836 4233 844
rect 4327 836 4813 844
rect 7307 836 8153 844
rect 8316 844 8324 853
rect 8316 836 8953 844
rect 9007 836 9713 844
rect 9727 836 9913 844
rect 10427 836 10533 844
rect 10867 836 10913 844
rect 1107 816 1284 824
rect 1807 816 1953 824
rect 1967 816 2113 824
rect 4627 816 4713 824
rect 5947 816 6213 824
rect 6787 816 7153 824
rect 7447 816 7853 824
rect 8207 816 10193 824
rect 827 796 1373 804
rect 1387 796 2333 804
rect 2347 796 2453 804
rect 5167 796 5313 804
rect 6247 796 6313 804
rect 6327 796 6553 804
rect 6627 796 7293 804
rect 7907 796 7933 804
rect 8047 796 8593 804
rect 8647 796 9173 804
rect 9287 796 9453 804
rect 9467 796 9533 804
rect 10287 796 10453 804
rect 10847 796 10953 804
rect 847 776 1333 784
rect 2547 776 2753 784
rect 3127 776 3633 784
rect 4147 776 4493 784
rect 4827 776 6113 784
rect 8007 776 8733 784
rect 10347 776 10713 784
rect 267 756 613 764
rect 2647 756 2673 764
rect 5407 756 5493 764
rect 6567 756 6593 764
rect 6707 756 6993 764
rect 7247 756 7313 764
rect 7787 756 7893 764
rect 8607 756 8993 764
rect 9047 756 9193 764
rect 9247 756 9693 764
rect 9867 756 10753 764
rect 207 736 673 744
rect 687 736 1033 744
rect 1847 736 2013 744
rect 3247 736 3873 744
rect 4127 736 4373 744
rect 5667 736 5793 744
rect 6147 736 6273 744
rect 6367 736 7013 744
rect 7027 736 8773 744
rect 10067 736 10393 744
rect 11067 736 11113 744
rect 1347 716 1473 724
rect 1887 716 2093 724
rect 2107 716 2293 724
rect 2707 716 2733 724
rect 2847 716 2973 724
rect 3107 716 3433 724
rect 4607 716 4653 724
rect 4827 716 4973 724
rect 4987 716 5053 724
rect 5287 716 5333 724
rect 5427 716 5573 724
rect 5647 716 5953 724
rect 6627 716 6813 724
rect 7527 716 8173 724
rect 8187 716 8313 724
rect 9527 716 10433 724
rect 147 697 393 705
rect 467 697 573 705
rect 1387 696 1433 704
rect 1627 696 1773 704
rect 2087 696 2213 704
rect 2407 696 2573 704
rect 2947 697 3013 705
rect 3487 696 3673 704
rect 3927 696 4153 704
rect 4227 696 4333 704
rect 4527 697 4573 705
rect 5007 696 5033 704
rect 5267 696 5473 704
rect 5527 696 5553 704
rect 5727 697 5773 705
rect 6447 697 6513 705
rect 6667 696 6733 704
rect 6987 697 7093 705
rect 7347 697 7453 705
rect 7607 696 7833 704
rect 7856 696 8113 704
rect 2536 676 3173 684
rect 147 655 213 663
rect 427 656 452 664
rect 487 655 793 663
rect 807 656 933 664
rect 987 655 1073 663
rect 1147 656 1273 664
rect 1287 656 1353 664
rect 1407 655 1452 663
rect 1487 656 1633 664
rect 1647 656 1813 664
rect 1827 655 1953 663
rect 2027 655 2053 663
rect 2107 656 2313 664
rect 2536 664 2544 676
rect 4396 676 5573 684
rect 2327 656 2544 664
rect 2567 655 2672 663
rect 2707 655 2733 663
rect 4396 666 4404 676
rect 5956 676 6033 684
rect 2827 656 2993 664
rect 3007 655 3113 663
rect 3267 656 3453 664
rect 3527 655 3653 663
rect 4607 655 4653 663
rect 4987 655 5053 663
rect 5287 656 5413 664
rect 5427 655 5453 663
rect 5956 664 5964 676
rect 7856 684 7864 696
rect 6827 676 6924 684
rect 5947 656 5964 664
rect 6916 666 6924 676
rect 7536 676 7864 684
rect 6007 656 6193 664
rect 6247 655 6273 663
rect 6387 655 6633 663
rect 6687 655 6773 663
rect 7536 666 7544 676
rect 8356 684 8364 694
rect 8427 696 8633 704
rect 8707 697 8773 705
rect 8887 696 9013 704
rect 9187 697 9253 705
rect 10207 697 10313 705
rect 10507 697 10533 705
rect 11067 697 11253 705
rect 8187 676 8364 684
rect 10447 676 10873 684
rect 10956 684 10964 694
rect 10887 676 10964 684
rect 7167 656 7533 664
rect 7927 656 7953 664
rect 8067 655 8093 663
rect 8387 655 8413 663
rect 9047 655 9073 663
rect 9127 656 9673 664
rect 9687 656 9852 664
rect 9887 655 9973 663
rect 10107 655 10153 663
rect 10227 655 10293 663
rect 10787 656 10973 664
rect 11087 655 11193 663
rect 827 636 873 644
rect 2336 636 2513 644
rect 187 616 253 624
rect 267 616 873 624
rect 1007 616 1533 624
rect 1547 616 1593 624
rect 2336 624 2344 636
rect 3907 636 4333 644
rect 4447 636 4793 644
rect 5587 636 5753 644
rect 5767 636 5804 644
rect 1787 616 2344 624
rect 2387 616 3033 624
rect 3047 616 3073 624
rect 3596 616 4093 624
rect 607 596 833 604
rect 1047 596 1153 604
rect 3596 604 3604 616
rect 4147 616 4293 624
rect 4527 616 4613 624
rect 5507 616 5773 624
rect 5796 624 5804 636
rect 5987 636 6013 644
rect 7127 636 7353 644
rect 8467 636 8793 644
rect 10347 636 10553 644
rect 5796 616 6212 624
rect 6247 616 7432 624
rect 7467 616 7793 624
rect 8047 616 8333 624
rect 8347 616 8613 624
rect 8947 616 8993 624
rect 9007 616 9313 624
rect 9727 616 10193 624
rect 10707 616 11133 624
rect 11147 616 11233 624
rect 2687 596 3604 604
rect 3627 596 3693 604
rect 4347 596 5233 604
rect 5367 596 6753 604
rect 6847 596 7953 604
rect 8107 596 8173 604
rect 1607 576 1853 584
rect 2407 576 3213 584
rect 5687 576 6624 584
rect 6616 564 6624 576
rect 7067 576 8873 584
rect 9807 576 10153 584
rect 10167 576 10633 584
rect 1447 556 1584 564
rect 6616 556 6813 564
rect 607 536 733 544
rect 1576 544 1584 556
rect 7767 556 7893 564
rect 8767 556 10333 564
rect 1576 536 2673 544
rect 2747 536 3833 544
rect 4567 536 5693 544
rect 5767 536 6593 544
rect 6607 536 8052 544
rect 8087 536 8553 544
rect 9267 536 10713 544
rect 7007 516 7353 524
rect 7587 516 7613 524
rect 7636 516 9233 524
rect 2467 496 2773 504
rect 6647 496 6793 504
rect 6807 496 7533 504
rect 7636 504 7644 516
rect 7547 496 7644 504
rect 7967 496 8173 504
rect 8307 496 8853 504
rect 8867 496 9173 504
rect 9307 496 9453 504
rect 9467 496 9553 504
rect 9567 496 9793 504
rect 9807 496 9913 504
rect 10367 496 11013 504
rect 3067 476 3093 484
rect 3107 476 3613 484
rect 3967 476 4353 484
rect 6787 476 7313 484
rect 7367 476 7933 484
rect 8587 476 9333 484
rect 10027 476 10213 484
rect 227 456 753 464
rect 1587 456 1933 464
rect 2867 456 3573 464
rect 3587 456 6733 464
rect 10287 456 10393 464
rect 10787 456 11053 464
rect 387 436 453 444
rect 2347 436 2813 444
rect 3367 436 3553 444
rect 4107 436 4193 444
rect 4247 436 4833 444
rect 5267 436 5493 444
rect 5867 436 5953 444
rect 7027 436 7133 444
rect 7827 436 7993 444
rect 8127 436 8193 444
rect 8596 436 8993 444
rect 1747 416 1833 424
rect 2807 416 3553 424
rect 3707 416 3953 424
rect 4467 416 4733 424
rect 5147 416 5553 424
rect 127 397 153 405
rect 347 397 413 405
rect 2147 396 2413 404
rect 2927 396 3193 404
rect 4167 396 4313 404
rect 1707 376 1813 384
rect 3656 384 3664 394
rect 5067 396 5193 404
rect 3656 376 3733 384
rect 4396 384 4404 394
rect 5307 396 5693 404
rect 5927 397 5993 405
rect 6427 397 6473 405
rect 6547 396 6593 404
rect 6887 397 6913 405
rect 6967 396 7093 404
rect 7207 396 7333 404
rect 7407 396 7573 404
rect 7587 396 7753 404
rect 8596 404 8604 436
rect 9587 436 10013 444
rect 10087 436 10493 444
rect 10507 436 10593 444
rect 8627 416 9293 424
rect 9347 416 9653 424
rect 9667 416 9753 424
rect 10347 416 10813 424
rect 11107 416 11133 424
rect 8407 396 8604 404
rect 4396 376 4493 384
rect 7996 384 8004 394
rect 8396 384 8404 394
rect 8667 396 8793 404
rect 8807 396 8873 404
rect 8967 397 9033 405
rect 9047 396 9153 404
rect 9467 396 9813 404
rect 9887 396 10093 404
rect 10407 397 10473 405
rect 10767 397 10853 405
rect 10987 397 11053 405
rect 4636 376 5504 384
rect 7996 376 8404 384
rect 8996 376 9393 384
rect 107 356 173 364
rect 407 356 533 364
rect 887 355 1013 363
rect 2167 355 2213 363
rect 2347 355 2393 363
rect 2487 355 2653 363
rect 2847 355 2873 363
rect 3127 356 3233 364
rect 4636 366 4644 376
rect 3587 355 3613 363
rect 3947 356 4133 364
rect 4387 355 4453 363
rect 4527 355 4593 363
rect 4827 355 4893 363
rect 4947 355 5073 363
rect 5207 355 5273 363
rect 5496 364 5504 376
rect 5496 356 5533 364
rect 5667 355 5713 363
rect 6007 356 6373 364
rect 6387 355 6433 363
rect 6487 356 6553 364
rect 6567 356 6613 364
rect 6807 355 6833 363
rect 6927 356 7113 364
rect 7127 355 7393 363
rect 7567 356 7613 364
rect 7687 355 7733 363
rect 7787 355 7813 363
rect 7927 356 7973 364
rect 8127 355 8173 363
rect 8647 356 8753 364
rect 8996 364 9004 376
rect 9256 366 9264 376
rect 10396 376 10693 384
rect 8827 356 9004 364
rect 9027 356 9213 364
rect 9827 355 9853 363
rect 9947 356 10073 364
rect 10087 355 10113 363
rect 10396 364 10404 376
rect 10387 356 10404 364
rect 10427 355 10453 363
rect 10627 356 10752 364
rect 10787 356 10833 364
rect 10887 355 10973 363
rect 1147 336 1233 344
rect 2447 336 2853 344
rect 3267 336 3604 344
rect 767 316 1053 324
rect 1067 316 1333 324
rect 1967 316 3293 324
rect 3596 324 3604 336
rect 5107 336 5393 344
rect 5407 336 5473 344
rect 8747 336 8813 344
rect 8867 336 9433 344
rect 9447 336 9673 344
rect 9687 336 9733 344
rect 9907 336 10053 344
rect 3596 316 3673 324
rect 3747 316 4633 324
rect 4827 316 5033 324
rect 5547 316 5933 324
rect 6287 316 6773 324
rect 7087 316 7193 324
rect 7367 316 7673 324
rect 7867 316 8673 324
rect 9867 316 10293 324
rect 11087 316 11153 324
rect 607 296 1313 304
rect 1327 296 2193 304
rect 2667 296 2793 304
rect 2867 296 3253 304
rect 3767 296 4313 304
rect 5967 296 6793 304
rect 7927 296 8133 304
rect 8147 296 8373 304
rect 8387 296 8513 304
rect 8627 296 8953 304
rect 9187 296 9393 304
rect 9587 296 10333 304
rect 427 276 833 284
rect 847 276 913 284
rect 927 276 1253 284
rect 2627 276 3253 284
rect 3267 276 3373 284
rect 3567 276 4813 284
rect 4867 276 5233 284
rect 6367 276 6953 284
rect 9147 276 9653 284
rect 767 256 793 264
rect 1227 256 4413 264
rect 4907 256 5173 264
rect 5527 256 5893 264
rect 5907 256 6313 264
rect 7107 256 7433 264
rect 7447 256 8113 264
rect 8127 256 8433 264
rect 8607 256 8853 264
rect 9407 256 9453 264
rect 9747 256 10473 264
rect 3307 236 3753 244
rect 3967 236 4173 244
rect 5487 236 6353 244
rect 6867 236 7933 244
rect 7947 236 8093 244
rect 8227 236 8493 244
rect 8507 236 9333 244
rect 9607 236 11053 244
rect 127 216 173 224
rect 187 216 413 224
rect 827 216 973 224
rect 1707 216 2093 224
rect 2107 216 2293 224
rect 2407 216 2813 224
rect 2887 216 3273 224
rect 7327 216 7913 224
rect 4667 196 4953 204
rect 5907 196 6133 204
rect 8727 196 8913 204
rect 9447 196 9553 204
rect 227 176 333 184
rect 347 176 593 184
rect 947 176 1404 184
rect 1396 168 1404 176
rect 2567 177 2613 185
rect 2847 177 2913 185
rect 3327 177 3473 185
rect 1127 155 1213 163
rect 1267 157 1333 165
rect 1407 156 2133 164
rect 2147 157 2733 165
rect 3516 164 3524 174
rect 3567 176 3693 184
rect 3747 177 3793 185
rect 4107 177 4133 185
rect 4187 176 4253 184
rect 4096 164 4104 174
rect 4307 176 4373 184
rect 4427 177 4473 185
rect 4627 176 4893 184
rect 4967 177 5093 185
rect 5167 177 5213 185
rect 5707 177 5753 185
rect 5867 177 5893 185
rect 6167 176 6313 184
rect 3516 156 4104 164
rect 407 136 453 144
rect 627 136 753 144
rect 767 136 793 144
rect 2427 136 2553 144
rect 2647 135 2713 143
rect 2927 136 3033 144
rect 3207 135 3233 143
rect 3507 136 3713 144
rect 3767 136 3933 144
rect 4207 135 4233 143
rect 4327 135 4393 143
rect 4447 136 4493 144
rect 4507 136 4853 144
rect 4927 135 5133 143
rect 5327 136 5493 144
rect 5727 136 5853 144
rect 5927 136 6013 144
rect 6127 136 6273 144
rect 6336 146 6344 193
rect 6427 176 6573 184
rect 6807 176 6953 184
rect 7067 176 7233 184
rect 7247 176 7313 184
rect 7487 177 7513 185
rect 7667 176 7853 184
rect 7907 177 8153 185
rect 8527 176 8744 184
rect 8736 164 8744 176
rect 8767 176 8893 184
rect 8987 176 9133 184
rect 9207 176 9393 184
rect 9407 176 9573 184
rect 8736 156 9593 164
rect 6387 135 6413 143
rect 6647 136 6773 144
rect 6787 135 6853 143
rect 6967 135 6993 143
rect 7187 135 7253 143
rect 7267 136 7633 144
rect 7647 136 7833 144
rect 7887 136 7933 144
rect 9456 146 9464 156
rect 10147 157 10173 165
rect 10227 155 10373 163
rect 8587 135 8733 143
rect 8787 135 8873 143
rect 8927 135 8953 143
rect 9327 135 9413 143
rect 9647 136 9713 144
rect 9807 135 9873 143
rect 10027 135 10053 143
rect 10747 135 10873 143
rect 11147 135 11333 143
rect 207 116 473 124
rect 1807 116 2093 124
rect 2607 116 2753 124
rect 4167 116 4293 124
rect 5247 116 5653 124
rect 8087 116 8153 124
rect 8167 116 8413 124
rect 8427 116 9173 124
rect 9187 116 9213 124
rect 10107 116 10233 124
rect 10547 115 10673 123
rect 847 96 913 104
rect 3807 96 4633 104
rect 6567 96 6933 104
rect 6947 96 8033 104
rect 8447 96 8993 104
rect 9347 96 9933 104
rect 10767 96 11313 104
rect 1287 76 1733 84
rect 1747 76 1853 84
rect 1967 76 4253 84
rect 6447 76 8633 84
rect 8887 76 8973 84
rect 9147 76 9313 84
rect 9567 76 9673 84
rect 1587 56 3553 64
rect 4487 56 5173 64
rect 6827 56 7093 64
rect 7467 56 8533 64
rect 8547 56 8613 64
rect 8747 56 9533 64
rect 9547 56 9693 64
rect 7847 36 8113 44
rect 8127 36 8573 44
rect 8907 36 9733 44
rect 9787 36 11093 44
rect 7047 16 7513 24
rect 7527 16 7673 24
rect 7687 16 8593 24
rect 8987 16 9633 24
use INVX1  _1668_ ~/ETRI050_DesignKit/devel/Ref_Design/CPU_6502/layout/digital_ETRI
timestamp 1701862152
transform 1 0 6830 0 -1 3390
box -12 -8 52 272
use NAND2X1  _1669_ ~/ETRI050_DesignKit/devel/Ref_Design/CPU_6502/layout/digital_ETRI
timestamp 1702508443
transform -1 0 6930 0 -1 790
box -12 -8 72 272
use OAI21X1  _1670_ ~/ETRI050_DesignKit/devel/Ref_Design/CPU_6502/layout/digital_ETRI
timestamp 1702508443
transform 1 0 6670 0 -1 2870
box -12 -8 92 272
use INVX1  _1671_
timestamp 1701862152
transform -1 0 6490 0 -1 8590
box -12 -8 52 272
use NAND2X1  _1672_
timestamp 1702508443
transform 1 0 6030 0 -1 10670
box -12 -8 72 272
use OAI21X1  _1673_
timestamp 1702508443
transform 1 0 6430 0 1 8590
box -12 -8 92 272
use INVX8  _1674_ ~/ETRI050_DesignKit/devel/Ref_Design/CPU_6502/layout/digital_ETRI
timestamp 1701862152
transform -1 0 6590 0 -1 9110
box -12 -8 114 272
use OR2X2  _1675_ ~/ETRI050_DesignKit/devel/Ref_Design/CPU_6502/layout/digital_ETRI
timestamp 1702508443
transform 1 0 150 0 -1 5470
box -12 -8 92 272
use OAI21X1  _1676_
timestamp 1702508443
transform -1 0 470 0 -1 5470
box -12 -8 92 272
use INVX1  _1677_
timestamp 1701862152
transform -1 0 670 0 1 5470
box -12 -8 52 272
use INVX1  _1678_
timestamp 1701862152
transform 1 0 170 0 -1 10670
box -12 -8 52 272
use NAND2X1  _1679_
timestamp 1702508443
transform -1 0 430 0 -1 11190
box -12 -8 72 272
use OAI21X1  _1680_
timestamp 1702508443
transform 1 0 370 0 -1 10670
box -12 -8 92 272
use INVX1  _1681_
timestamp 1701862152
transform -1 0 210 0 -1 7030
box -12 -8 52 272
use NAND2X1  _1682_
timestamp 1702508443
transform -1 0 210 0 1 7030
box -12 -8 72 272
use OAI21X1  _1683_
timestamp 1702508443
transform 1 0 170 0 1 6510
box -12 -8 92 272
use OR2X2  _1684_
timestamp 1702508443
transform 1 0 1050 0 -1 11190
box -12 -8 92 272
use OAI21X1  _1685_
timestamp 1702508443
transform -1 0 1370 0 -1 11190
box -12 -8 92 272
use INVX1  _1686_
timestamp 1701862152
transform -1 0 1130 0 1 10670
box -12 -8 52 272
use OR2X2  _1687_
timestamp 1702508443
transform 1 0 1530 0 -1 11190
box -12 -8 92 272
use OAI21X1  _1688_
timestamp 1702508443
transform -1 0 1850 0 -1 11190
box -12 -8 92 272
use INVX1  _1689_
timestamp 1701862152
transform -1 0 2070 0 1 10150
box -12 -8 52 272
use MUX2X1  _1690_ ~/ETRI050_DesignKit/devel/Ref_Design/CPU_6502/layout/digital_ETRI
timestamp 1701862152
transform 1 0 2190 0 1 9110
box -12 -8 114 272
use INVX1  _1691_
timestamp 1701862152
transform -1 0 2250 0 -1 9110
box -12 -8 52 272
use INVX1  _1692_
timestamp 1701862152
transform 1 0 170 0 1 790
box -12 -8 52 272
use NAND2X1  _1693_
timestamp 1702508443
transform 1 0 170 0 -1 1310
box -12 -8 72 272
use INVX1  _1694_
timestamp 1701862152
transform 1 0 590 0 -1 270
box -12 -8 52 272
use NAND2X1  _1695_
timestamp 1702508443
transform -1 0 850 0 -1 270
box -12 -8 72 272
use NOR2X1  _1696_ ~/ETRI050_DesignKit/devel/Ref_Design/CPU_6502/layout/digital_ETRI
timestamp 1701862152
transform 1 0 1230 0 1 2870
box -12 -8 74 272
use INVX2  _1697_ ~/ETRI050_DesignKit/devel/Ref_Design/CPU_6502/layout/digital_ETRI
timestamp 1701862152
transform -1 0 2890 0 -1 2870
box -12 -8 52 272
use NOR2X1  _1698_
timestamp 1701862152
transform -1 0 2030 0 1 3390
box -12 -8 74 272
use NAND2X1  _1699_
timestamp 1702508443
transform 1 0 3910 0 1 3390
box -12 -8 72 272
use NOR2X1  _1700_
timestamp 1701862152
transform -1 0 2750 0 -1 3910
box -12 -8 74 272
use AND2X2  _1701_ ~/ETRI050_DesignKit/devel/Ref_Design/CPU_6502/layout/digital_ETRI
timestamp 1701862152
transform -1 0 1310 0 1 270
box -12 -8 94 272
use NOR2X1  _1702_
timestamp 1701862152
transform 1 0 1010 0 1 270
box -12 -8 74 272
use NAND3X1  _1703_ ~/ETRI050_DesignKit/devel/Ref_Design/CPU_6502/layout/digital_ETRI
timestamp 1702508443
transform -1 0 1550 0 1 1830
box -12 -8 92 272
use NOR2X1  _1704_
timestamp 1701862152
transform -1 0 9270 0 1 2870
box -12 -8 74 272
use INVX4  _1705_ ~/ETRI050_DesignKit/devel/Ref_Design/CPU_6502/layout/digital_ETRI
timestamp 1701862152
transform 1 0 9870 0 -1 790
box -12 -8 72 272
use NOR2X1  _1706_
timestamp 1701862152
transform -1 0 8130 0 -1 4950
box -12 -8 74 272
use INVX1  _1707_
timestamp 1701862152
transform 1 0 8530 0 -1 4950
box -12 -8 52 272
use INVX1  _1708_
timestamp 1701862152
transform 1 0 5150 0 -1 5990
box -12 -8 52 272
use INVX1  _1709_
timestamp 1701862152
transform -1 0 11270 0 1 5990
box -12 -8 52 272
use INVX1  _1710_
timestamp 1701862152
transform 1 0 5530 0 -1 5470
box -12 -8 52 272
use NAND2X1  _1711_
timestamp 1702508443
transform -1 0 5390 0 -1 5990
box -12 -8 72 272
use OAI21X1  _1712_
timestamp 1702508443
transform -1 0 5250 0 1 5470
box -12 -8 92 272
use OAI21X1  _1713_
timestamp 1702508443
transform 1 0 8050 0 1 4430
box -12 -8 92 272
use NAND2X1  _1714_
timestamp 1702508443
transform 1 0 7850 0 1 4950
box -12 -8 72 272
use OAI21X1  _1715_
timestamp 1702508443
transform -1 0 8150 0 1 4950
box -12 -8 92 272
use NAND2X1  _1716_
timestamp 1702508443
transform -1 0 8350 0 1 4430
box -12 -8 72 272
use OAI21X1  _1717_
timestamp 1702508443
transform -1 0 8150 0 1 1310
box -12 -8 92 272
use OAI21X1  _1718_
timestamp 1702508443
transform -1 0 6090 0 1 5990
box -12 -8 92 272
use INVX1  _1719_
timestamp 1701862152
transform -1 0 6890 0 -1 5990
box -12 -8 52 272
use AOI21X1  _1720_ ~/ETRI050_DesignKit/devel/Ref_Design/CPU_6502/layout/digital_ETRI
timestamp 1702508443
transform -1 0 6930 0 1 5470
box -12 -8 92 272
use OAI21X1  _1721_
timestamp 1702508443
transform -1 0 7170 0 1 5470
box -12 -8 92 272
use MUX2X1  _1722_
timestamp 1701862152
transform -1 0 7890 0 1 4430
box -12 -8 114 272
use OAI21X1  _1723_
timestamp 1702508443
transform 1 0 8030 0 1 1830
box -12 -8 92 272
use NOR2X1  _1724_
timestamp 1701862152
transform -1 0 8110 0 -1 1310
box -12 -8 74 272
use INVX1  _1725_
timestamp 1701862152
transform 1 0 6670 0 1 5990
box -12 -8 52 272
use AOI21X1  _1726_
timestamp 1702508443
transform 1 0 6850 0 1 5990
box -12 -8 92 272
use OAI21X1  _1727_
timestamp 1702508443
transform -1 0 7170 0 1 5990
box -12 -8 92 272
use NAND2X1  _1728_
timestamp 1702508443
transform 1 0 7810 0 1 5990
box -12 -8 72 272
use OAI21X1  _1729_
timestamp 1702508443
transform -1 0 7810 0 -1 5990
box -12 -8 92 272
use NAND2X1  _1730_
timestamp 1702508443
transform -1 0 8270 0 1 3390
box -12 -8 72 272
use NAND2X1  _1731_
timestamp 1702508443
transform -1 0 8130 0 -1 270
box -12 -8 72 272
use NAND2X1  _1732_
timestamp 1702508443
transform -1 0 8090 0 1 5470
box -12 -8 72 272
use OAI21X1  _1733_
timestamp 1702508443
transform -1 0 8310 0 1 5470
box -12 -8 92 272
use NAND2X1  _1734_
timestamp 1702508443
transform 1 0 8230 0 -1 5470
box -12 -8 72 272
use NAND2X1  _1735_
timestamp 1702508443
transform 1 0 8690 0 -1 5470
box -12 -8 72 272
use OAI21X1  _1736_
timestamp 1702508443
transform 1 0 8530 0 1 4950
box -12 -8 92 272
use AND2X2  _1737_
timestamp 1701862152
transform -1 0 8670 0 -1 3910
box -12 -8 94 272
use NAND2X1  _1738_
timestamp 1702508443
transform 1 0 9010 0 1 790
box -12 -8 72 272
use NOR2X1  _1739_
timestamp 1701862152
transform -1 0 9270 0 -1 790
box -12 -8 74 272
use NAND2X1  _1740_
timestamp 1702508443
transform 1 0 6590 0 1 270
box -12 -8 72 272
use OAI22X1  _1741_ ~/ETRI050_DesignKit/devel/Ref_Design/CPU_6502/layout/digital_ETRI
timestamp 1701862152
transform 1 0 6470 0 1 790
box -12 -8 112 272
use INVX1  _1742_
timestamp 1701862152
transform -1 0 6450 0 -1 790
box -12 -8 52 272
use NAND2X1  _1743_
timestamp 1702508443
transform -1 0 2470 0 -1 3390
box -12 -8 72 272
use INVX4  _1744_
timestamp 1701862152
transform 1 0 410 0 -1 4950
box -12 -8 72 272
use NAND2X1  _1745_
timestamp 1702508443
transform 1 0 2230 0 -1 3910
box -12 -8 72 272
use NOR2X1  _1746_
timestamp 1701862152
transform -1 0 5290 0 -1 3390
box -12 -8 74 272
use INVX1  _1747_
timestamp 1701862152
transform -1 0 430 0 -1 270
box -12 -8 52 272
use NOR2X1  _1748_
timestamp 1701862152
transform -1 0 630 0 1 270
box -12 -8 74 272
use NAND2X1  _1749_
timestamp 1702508443
transform -1 0 1090 0 1 1310
box -12 -8 72 272
use NOR2X1  _1750_
timestamp 1701862152
transform -1 0 1310 0 1 1310
box -12 -8 74 272
use NAND2X1  _1751_
timestamp 1702508443
transform -1 0 4670 0 -1 2870
box -12 -8 72 272
use OAI22X1  _1752_
timestamp 1701862152
transform 1 0 4830 0 -1 2870
box -12 -8 112 272
use INVX1  _1753_
timestamp 1701862152
transform -1 0 4470 0 1 790
box -12 -8 52 272
use INVX1  _1754_
timestamp 1701862152
transform 1 0 390 0 -1 790
box -12 -8 52 272
use NOR2X1  _1755_
timestamp 1701862152
transform -1 0 630 0 -1 790
box -12 -8 74 272
use NOR2X1  _1756_
timestamp 1701862152
transform -1 0 230 0 -1 270
box -12 -8 74 272
use NAND2X1  _1757_
timestamp 1702508443
transform 1 0 790 0 -1 790
box -12 -8 72 272
use INVX2  _1758_
timestamp 1701862152
transform 1 0 170 0 1 2350
box -12 -8 52 272
use NOR2X1  _1759_
timestamp 1701862152
transform -1 0 2710 0 -1 2870
box -12 -8 74 272
use INVX1  _1760_
timestamp 1701862152
transform 1 0 3050 0 -1 2870
box -12 -8 52 272
use INVX8  _1761_
timestamp 1701862152
transform -1 0 3450 0 -1 3390
box -12 -8 114 272
use NAND2X1  _1762_
timestamp 1702508443
transform -1 0 210 0 1 270
box -12 -8 72 272
use NAND2X1  _1763_
timestamp 1702508443
transform 1 0 170 0 -1 790
box -12 -8 72 272
use NOR2X1  _1764_
timestamp 1701862152
transform 1 0 610 0 1 1310
box -12 -8 74 272
use INVX1  _1765_
timestamp 1701862152
transform 1 0 1470 0 1 1310
box -12 -8 52 272
use NOR2X1  _1766_
timestamp 1701862152
transform -1 0 3310 0 -1 1830
box -12 -8 74 272
use INVX8  _1767_
timestamp 1701862152
transform 1 0 1570 0 -1 4430
box -12 -8 114 272
use NAND2X1  _1768_
timestamp 1702508443
transform 1 0 390 0 -1 1310
box -12 -8 72 272
use NOR2X1  _1769_
timestamp 1701862152
transform -1 0 650 0 1 1830
box -12 -8 74 272
use NAND2X1  _1770_
timestamp 1702508443
transform 1 0 2190 0 -1 3390
box -12 -8 72 272
use OAI21X1  _1771_
timestamp 1702508443
transform -1 0 2530 0 -1 3910
box -12 -8 92 272
use NOR2X1  _1772_
timestamp 1701862152
transform -1 0 3170 0 -1 3910
box -12 -8 74 272
use OAI21X1  _1773_
timestamp 1702508443
transform 1 0 4030 0 1 2870
box -12 -8 92 272
use AOI21X1  _1774_
timestamp 1702508443
transform -1 0 5470 0 -1 2350
box -12 -8 92 272
use NAND2X1  _1775_
timestamp 1702508443
transform 1 0 370 0 1 790
box -12 -8 72 272
use NOR2X1  _1776_
timestamp 1701862152
transform -1 0 450 0 1 1310
box -12 -8 74 272
use INVX2  _1777_
timestamp 1701862152
transform 1 0 810 0 -1 1830
box -12 -8 52 272
use NOR2X1  _1778_
timestamp 1701862152
transform -1 0 4590 0 1 5470
box -12 -8 74 272
use INVX2  _1779_
timestamp 1701862152
transform -1 0 6210 0 -1 5470
box -12 -8 52 272
use OAI21X1  _1780_
timestamp 1702508443
transform 1 0 4910 0 1 2870
box -12 -8 92 272
use INVX1  _1781_
timestamp 1701862152
transform 1 0 4490 0 1 2870
box -12 -8 52 272
use NOR2X1  _1782_
timestamp 1701862152
transform -1 0 230 0 1 1310
box -12 -8 74 272
use OAI21X1  _1783_
timestamp 1702508443
transform -1 0 1530 0 1 2870
box -12 -8 92 272
use OAI21X1  _1784_
timestamp 1702508443
transform -1 0 5210 0 1 2870
box -12 -8 92 272
use OR2X2  _1785_
timestamp 1702508443
transform 1 0 5090 0 -1 2870
box -12 -8 92 272
use OAI21X1  _1786_
timestamp 1702508443
transform -1 0 5230 0 -1 2350
box -12 -8 92 272
use INVX1  _1787_
timestamp 1701862152
transform 1 0 5150 0 1 2350
box -12 -8 52 272
use NOR2X1  _1788_
timestamp 1701862152
transform -1 0 4990 0 -1 2350
box -12 -8 74 272
use INVX1  _1789_
timestamp 1701862152
transform 1 0 170 0 1 1830
box -12 -8 52 272
use NOR2X1  _1790_
timestamp 1701862152
transform -1 0 450 0 -1 2350
box -12 -8 74 272
use NAND2X1  _1791_
timestamp 1702508443
transform -1 0 2250 0 -1 2350
box -12 -8 72 272
use NOR2X1  _1792_
timestamp 1701862152
transform -1 0 3610 0 -1 2350
box -12 -8 74 272
use NAND2X1  _1793_
timestamp 1702508443
transform -1 0 4730 0 1 1830
box -12 -8 72 272
use AND2X2  _1794_
timestamp 1701862152
transform 1 0 1010 0 1 1830
box -12 -8 94 272
use NAND2X1  _1795_
timestamp 1702508443
transform -1 0 2310 0 1 2350
box -12 -8 72 272
use AOI21X1  _1796_
timestamp 1702508443
transform -1 0 1950 0 -1 1830
box -12 -8 92 272
use AOI21X1  _1797_
timestamp 1702508443
transform 1 0 2110 0 -1 1830
box -12 -8 92 272
use NAND2X1  _1798_
timestamp 1702508443
transform 1 0 1030 0 -1 1310
box -12 -8 72 272
use NOR2X1  _1799_
timestamp 1701862152
transform 1 0 3830 0 1 3910
box -12 -8 74 272
use AOI21X1  _1800_
timestamp 1702508443
transform 1 0 3530 0 1 1830
box -12 -8 92 272
use NAND2X1  _1801_
timestamp 1702508443
transform -1 0 1310 0 1 1830
box -12 -8 72 272
use NOR2X1  _1802_
timestamp 1701862152
transform -1 0 3850 0 1 2350
box -12 -8 74 272
use OAI21X1  _1803_
timestamp 1702508443
transform -1 0 4090 0 1 2350
box -12 -8 92 272
use OAI21X1  _1804_
timestamp 1702508443
transform -1 0 4330 0 1 2350
box -12 -8 92 272
use INVX1  _1805_
timestamp 1701862152
transform 1 0 5570 0 1 2350
box -12 -8 52 272
use NOR2X1  _1806_
timestamp 1701862152
transform -1 0 4990 0 1 2350
box -12 -8 74 272
use NOR2X1  _1807_
timestamp 1701862152
transform -1 0 5410 0 1 2350
box -12 -8 74 272
use NAND3X1  _1808_
timestamp 1702508443
transform 1 0 4890 0 1 1830
box -12 -8 92 272
use INVX2  _1809_
timestamp 1701862152
transform -1 0 7270 0 -1 270
box -12 -8 52 272
use NOR2X1  _1810_
timestamp 1701862152
transform -1 0 7270 0 1 1310
box -12 -8 74 272
use NOR2X1  _1811_
timestamp 1701862152
transform 1 0 7570 0 -1 1830
box -12 -8 74 272
use NAND2X1  _1812_
timestamp 1702508443
transform -1 0 7690 0 -1 1310
box -12 -8 72 272
use INVX1  _1813_
timestamp 1701862152
transform 1 0 9210 0 1 790
box -12 -8 52 272
use NOR2X1  _1814_
timestamp 1701862152
transform -1 0 8310 0 -1 1830
box -12 -8 74 272
use NAND2X1  _1815_
timestamp 1702508443
transform 1 0 8470 0 1 2350
box -12 -8 72 272
use INVX2  _1816_
timestamp 1701862152
transform -1 0 9770 0 -1 2350
box -12 -8 52 272
use NAND2X1  _1817_
timestamp 1702508443
transform -1 0 9510 0 1 1310
box -12 -8 72 272
use INVX1  _1818_
timestamp 1701862152
transform -1 0 9690 0 1 270
box -12 -8 52 272
use OAI21X1  _1819_
timestamp 1702508443
transform -1 0 8550 0 -1 1830
box -12 -8 92 272
use OAI21X1  _1820_
timestamp 1702508443
transform -1 0 8630 0 1 1310
box -12 -8 92 272
use AOI21X1  _1821_
timestamp 1702508443
transform -1 0 5050 0 1 1310
box -12 -8 92 272
use AND2X2  _1822_
timestamp 1701862152
transform -1 0 4870 0 -1 790
box -12 -8 94 272
use NAND3X1  _1823_
timestamp 1702508443
transform -1 0 4410 0 -1 790
box -12 -8 92 272
use NOR2X1  _1824_
timestamp 1701862152
transform 1 0 4730 0 1 2350
box -12 -8 74 272
use NAND2X1  _1825_
timestamp 1702508443
transform 1 0 5790 0 1 1830
box -12 -8 72 272
use INVX1  _1826_
timestamp 1701862152
transform 1 0 8290 0 -1 270
box -12 -8 52 272
use NOR2X1  _1827_
timestamp 1701862152
transform 1 0 9430 0 -1 790
box -12 -8 74 272
use NAND3X1  _1828_
timestamp 1702508443
transform 1 0 8570 0 1 270
box -12 -8 92 272
use OAI21X1  _1829_
timestamp 1702508443
transform 1 0 5890 0 1 270
box -12 -8 92 272
use NAND2X1  _1830_
timestamp 1702508443
transform 1 0 3330 0 1 4430
box -12 -8 72 272
use NAND2X1  _1831_
timestamp 1702508443
transform -1 0 8150 0 -1 790
box -12 -8 72 272
use OAI22X1  _1832_
timestamp 1701862152
transform 1 0 6610 0 -1 790
box -12 -8 112 272
use NOR2X1  _1833_
timestamp 1701862152
transform -1 0 850 0 1 270
box -12 -8 74 272
use NAND2X1  _1834_
timestamp 1702508443
transform 1 0 1250 0 -1 1310
box -12 -8 72 272
use NOR2X1  _1835_
timestamp 1701862152
transform -1 0 2650 0 -1 1310
box -12 -8 74 272
use NAND2X1  _1836_
timestamp 1702508443
transform 1 0 1190 0 1 790
box -12 -8 72 272
use OAI21X1  _1837_
timestamp 1702508443
transform -1 0 2650 0 1 790
box -12 -8 92 272
use OAI21X1  _1838_
timestamp 1702508443
transform 1 0 2330 0 1 790
box -12 -8 92 272
use NAND2X1  _1839_
timestamp 1702508443
transform -1 0 430 0 1 270
box -12 -8 72 272
use NOR2X1  _1840_
timestamp 1701862152
transform -1 0 1070 0 1 2870
box -12 -8 74 272
use NAND2X1  _1841_
timestamp 1702508443
transform 1 0 3810 0 1 2870
box -12 -8 72 272
use NOR2X1  _1842_
timestamp 1701862152
transform -1 0 3090 0 -1 1830
box -12 -8 74 272
use NAND2X1  _1843_
timestamp 1702508443
transform -1 0 4070 0 -1 2350
box -12 -8 72 272
use OAI21X1  _1844_
timestamp 1702508443
transform 1 0 3930 0 -1 2870
box -12 -8 92 272
use NOR2X1  _1845_
timestamp 1701862152
transform -1 0 1910 0 -1 4950
box -12 -8 74 272
use NAND2X1  _1846_
timestamp 1702508443
transform 1 0 4230 0 1 4430
box -12 -8 72 272
use NAND2X1  _1847_
timestamp 1702508443
transform 1 0 3550 0 1 4430
box -12 -8 72 272
use OAI21X1  _1848_
timestamp 1702508443
transform 1 0 3990 0 1 4430
box -12 -8 92 272
use NOR2X1  _1849_
timestamp 1701862152
transform -1 0 4230 0 -1 2870
box -12 -8 74 272
use NAND2X1  _1850_
timestamp 1702508443
transform -1 0 1030 0 1 790
box -12 -8 72 272
use INVX2  _1851_
timestamp 1701862152
transform 1 0 1670 0 -1 1830
box -12 -8 52 272
use NAND2X1  _1852_
timestamp 1702508443
transform -1 0 2530 0 1 2350
box -12 -8 72 272
use NOR2X1  _1853_
timestamp 1701862152
transform 1 0 170 0 -1 2350
box -12 -8 74 272
use AOI21X1  _1854_
timestamp 1702508443
transform 1 0 2410 0 -1 2350
box -12 -8 92 272
use AOI21X1  _1855_
timestamp 1702508443
transform -1 0 2730 0 -1 2350
box -12 -8 92 272
use OAI21X1  _1856_
timestamp 1702508443
transform 1 0 1570 0 -1 790
box -12 -8 92 272
use OAI21X1  _1857_
timestamp 1702508443
transform -1 0 2810 0 -1 790
box -12 -8 92 272
use AOI21X1  _1858_
timestamp 1702508443
transform 1 0 2510 0 -1 790
box -12 -8 92 272
use NOR2X1  _1859_
timestamp 1701862152
transform 1 0 2290 0 -1 790
box -12 -8 74 272
use OAI21X1  _1860_
timestamp 1702508443
transform -1 0 1890 0 -1 790
box -12 -8 92 272
use OAI21X1  _1861_
timestamp 1702508443
transform -1 0 2130 0 -1 790
box -12 -8 92 272
use AND2X2  _1862_
timestamp 1701862152
transform -1 0 2210 0 1 270
box -12 -8 94 272
use NAND3X1  _1863_
timestamp 1702508443
transform 1 0 2370 0 1 270
box -12 -8 92 272
use NOR3X1  _1864_ ~/ETRI050_DesignKit/devel/Ref_Design/CPU_6502/layout/digital_ETRI
timestamp 1701862152
transform 1 0 3590 0 1 270
box -12 -8 172 272
use NOR2X1  _1865_
timestamp 1701862152
transform 1 0 7410 0 -1 1310
box -12 -8 74 272
use AOI22X1  _1866_ ~/ETRI050_DesignKit/devel/Ref_Design/CPU_6502/layout/digital_ETRI
timestamp 1701862152
transform 1 0 3770 0 -1 1310
box -14 -8 114 272
use NAND2X1  _1867_
timestamp 1702508443
transform 1 0 1230 0 -1 1830
box -12 -8 72 272
use INVX1  _1868_
timestamp 1701862152
transform 1 0 1670 0 1 1310
box -12 -8 52 272
use OAI21X1  _1869_
timestamp 1702508443
transform 1 0 2090 0 1 1310
box -12 -8 92 272
use OAI21X1  _1870_
timestamp 1702508443
transform -1 0 1770 0 -1 1310
box -12 -8 92 272
use AND2X2  _1871_
timestamp 1701862152
transform -1 0 2890 0 -1 1310
box -12 -8 94 272
use NOR2X1  _1872_
timestamp 1701862152
transform -1 0 630 0 1 790
box -12 -8 74 272
use INVX2  _1873_
timestamp 1701862152
transform 1 0 790 0 1 790
box -12 -8 52 272
use OAI21X1  _1874_
timestamp 1702508443
transform -1 0 1490 0 1 790
box -12 -8 92 272
use NOR3X1  _1875_
timestamp 1701862152
transform 1 0 1010 0 -1 790
box -12 -8 172 272
use OAI21X1  _1876_
timestamp 1702508443
transform 1 0 1330 0 -1 790
box -12 -8 92 272
use NOR2X1  _1877_
timestamp 1701862152
transform 1 0 2270 0 1 4950
box -12 -8 74 272
use INVX1  _1878_
timestamp 1701862152
transform 1 0 610 0 -1 1310
box -12 -8 52 272
use NAND2X1  _1879_
timestamp 1702508443
transform 1 0 810 0 1 1310
box -12 -8 72 272
use OAI21X1  _1880_
timestamp 1702508443
transform -1 0 2150 0 -1 4950
box -12 -8 92 272
use OAI21X1  _1881_
timestamp 1702508443
transform -1 0 2390 0 -1 4950
box -12 -8 92 272
use NOR3X1  _1882_
timestamp 1701862152
transform 1 0 1650 0 -1 3390
box -12 -8 172 272
use NOR3X1  _1883_
timestamp 1701862152
transform 1 0 1130 0 -1 3390
box -12 -8 172 272
use XOR2X1  _1884_ ~/ETRI050_DesignKit/devel/Ref_Design/CPU_6502/layout/digital_ETRI
timestamp 1702508443
transform -1 0 4250 0 1 3390
box -12 -8 132 272
use AND2X2  _1885_
timestamp 1701862152
transform -1 0 3930 0 -1 3390
box -12 -8 94 272
use AOI22X1  _1886_
timestamp 1701862152
transform 1 0 3590 0 -1 3390
box -14 -8 114 272
use AND2X2  _1887_
timestamp 1701862152
transform -1 0 3650 0 1 2870
box -12 -8 94 272
use NAND3X1  _1888_
timestamp 1702508443
transform -1 0 2690 0 1 270
box -12 -8 92 272
use NAND2X1  _1889_
timestamp 1702508443
transform 1 0 1770 0 -1 2870
box -12 -8 72 272
use INVX1  _1890_
timestamp 1701862152
transform -1 0 430 0 -1 1830
box -12 -8 52 272
use NAND2X1  _1891_
timestamp 1702508443
transform 1 0 170 0 -1 1830
box -12 -8 72 272
use NOR2X1  _1892_
timestamp 1701862152
transform 1 0 5010 0 -1 3390
box -12 -8 74 272
use NAND2X1  _1893_
timestamp 1702508443
transform 1 0 3990 0 1 1830
box -12 -8 72 272
use OAI21X1  _1894_
timestamp 1702508443
transform 1 0 4210 0 1 1830
box -12 -8 92 272
use INVX2  _1895_
timestamp 1701862152
transform -1 0 1970 0 1 1830
box -12 -8 52 272
use NAND2X1  _1896_
timestamp 1702508443
transform 1 0 1970 0 -1 2350
box -12 -8 72 272
use INVX1  _1897_
timestamp 1701862152
transform 1 0 3590 0 1 2350
box -12 -8 52 272
use NAND2X1  _1898_
timestamp 1702508443
transform 1 0 3370 0 1 2350
box -12 -8 72 272
use OAI21X1  _1899_
timestamp 1702508443
transform -1 0 3410 0 -1 2350
box -12 -8 92 272
use NOR2X1  _1900_
timestamp 1701862152
transform -1 0 4230 0 -1 1830
box -12 -8 74 272
use NAND2X1  _1901_
timestamp 1702508443
transform -1 0 850 0 1 1830
box -12 -8 72 272
use INVX1  _1902_
timestamp 1701862152
transform 1 0 5130 0 1 1830
box -12 -8 52 272
use OAI21X1  _1903_
timestamp 1702508443
transform 1 0 3450 0 1 1310
box -12 -8 92 272
use OAI21X1  _1904_
timestamp 1702508443
transform -1 0 3610 0 -1 1310
box -12 -8 92 272
use NAND2X1  _1905_
timestamp 1702508443
transform 1 0 3090 0 1 270
box -12 -8 72 272
use INVX1  _1906_
timestamp 1701862152
transform 1 0 370 0 1 2350
box -12 -8 52 272
use NOR2X1  _1907_
timestamp 1701862152
transform -1 0 3170 0 -1 2350
box -12 -8 74 272
use INVX1  _1908_
timestamp 1701862152
transform 1 0 6530 0 -1 2350
box -12 -8 52 272
use NOR2X1  _1909_
timestamp 1701862152
transform -1 0 6190 0 -1 2350
box -12 -8 74 272
use AOI22X1  _1910_
timestamp 1701862152
transform -1 0 5730 0 -1 2350
box -14 -8 114 272
use NOR2X1  _1911_
timestamp 1701862152
transform -1 0 850 0 1 2870
box -12 -8 74 272
use NAND2X1  _1912_
timestamp 1702508443
transform -1 0 3450 0 1 3910
box -12 -8 72 272
use NOR2X1  _1913_
timestamp 1701862152
transform -1 0 1170 0 -1 2870
box -12 -8 74 272
use NAND2X1  _1914_
timestamp 1702508443
transform -1 0 1610 0 1 3390
box -12 -8 72 272
use INVX1  _1915_
timestamp 1701862152
transform 1 0 2630 0 1 3390
box -12 -8 52 272
use NAND2X1  _1916_
timestamp 1702508443
transform -1 0 3550 0 1 3390
box -12 -8 72 272
use OAI21X1  _1917_
timestamp 1702508443
transform -1 0 4850 0 -1 3390
box -12 -8 92 272
use NAND2X1  _1918_
timestamp 1702508443
transform 1 0 1830 0 1 4950
box -12 -8 72 272
use NAND2X1  _1919_
timestamp 1702508443
transform -1 0 1390 0 -1 2870
box -12 -8 72 272
use INVX1  _1920_
timestamp 1701862152
transform -1 0 5150 0 1 4430
box -12 -8 52 272
use NAND2X1  _1921_
timestamp 1702508443
transform 1 0 4890 0 1 4430
box -12 -8 72 272
use OAI21X1  _1922_
timestamp 1702508443
transform -1 0 4730 0 1 4430
box -12 -8 92 272
use NOR2X1  _1923_
timestamp 1701862152
transform 1 0 4550 0 -1 3390
box -12 -8 74 272
use NAND2X1  _1924_
timestamp 1702508443
transform 1 0 2050 0 1 4950
box -12 -8 72 272
use INVX1  _1925_
timestamp 1701862152
transform 1 0 6190 0 -1 4430
box -12 -8 52 272
use NAND2X1  _1926_
timestamp 1702508443
transform 1 0 810 0 -1 1310
box -12 -8 72 272
use OAI21X1  _1927_
timestamp 1702508443
transform 1 0 3050 0 -1 1310
box -12 -8 92 272
use OAI21X1  _1928_
timestamp 1702508443
transform -1 0 3370 0 -1 1310
box -12 -8 92 272
use NAND3X1  _1929_
timestamp 1702508443
transform 1 0 3490 0 1 790
box -12 -8 92 272
use NOR3X1  _1930_
timestamp 1701862152
transform 1 0 3290 0 1 270
box -12 -8 172 272
use NAND2X1  _1931_
timestamp 1702508443
transform 1 0 3910 0 1 270
box -12 -8 72 272
use NOR2X1  _1932_
timestamp 1701862152
transform -1 0 4190 0 1 270
box -12 -8 74 272
use INVX1  _1933_
timestamp 1701862152
transform -1 0 1970 0 1 270
box -12 -8 52 272
use NAND2X1  _1934_
timestamp 1702508443
transform -1 0 5610 0 1 790
box -12 -8 72 272
use INVX1  _1935_
timestamp 1701862152
transform 1 0 5690 0 -1 270
box -12 -8 52 272
use NAND2X1  _1936_
timestamp 1702508443
transform -1 0 8490 0 1 3390
box -12 -8 72 272
use NAND2X1  _1937_
timestamp 1702508443
transform -1 0 7690 0 -1 270
box -12 -8 72 272
use NOR2X1  _1938_
timestamp 1701862152
transform -1 0 7910 0 -1 270
box -12 -8 74 272
use NAND2X1  _1939_
timestamp 1702508443
transform -1 0 6830 0 -1 270
box -12 -8 72 272
use NOR2X1  _1940_
timestamp 1701862152
transform -1 0 5950 0 -1 270
box -12 -8 74 272
use NAND2X1  _1941_
timestamp 1702508443
transform 1 0 5930 0 -1 790
box -12 -8 72 272
use INVX1  _1942_
timestamp 1701862152
transform 1 0 4910 0 -1 1310
box -12 -8 52 272
use NOR2X1  _1943_
timestamp 1701862152
transform 1 0 8170 0 1 270
box -12 -8 74 272
use NOR2X1  _1944_
timestamp 1701862152
transform -1 0 8430 0 1 270
box -12 -8 74 272
use NAND2X1  _1945_
timestamp 1702508443
transform 1 0 7950 0 1 270
box -12 -8 72 272
use NOR2X1  _1946_
timestamp 1701862152
transform -1 0 6190 0 1 270
box -12 -8 74 272
use AOI22X1  _1947_
timestamp 1701862152
transform -1 0 6250 0 -1 790
box -14 -8 114 272
use NAND3X1  _1948_
timestamp 1702508443
transform 1 0 5450 0 -1 790
box -12 -8 92 272
use NAND2X1  _1949_
timestamp 1702508443
transform 1 0 4690 0 -1 1310
box -12 -8 72 272
use NAND3X1  _1950_
timestamp 1702508443
transform -1 0 8390 0 -1 790
box -12 -8 92 272
use NAND2X1  _1951_
timestamp 1702508443
transform 1 0 610 0 -1 2350
box -12 -8 72 272
use NAND2X1  _1952_
timestamp 1702508443
transform -1 0 5810 0 1 2350
box -12 -8 72 272
use OAI21X1  _1953_
timestamp 1702508443
transform 1 0 5890 0 -1 2350
box -12 -8 92 272
use INVX1  _1954_
timestamp 1701862152
transform 1 0 8270 0 -1 1310
box -12 -8 52 272
use NAND2X1  _1955_
timestamp 1702508443
transform -1 0 8850 0 1 1310
box -12 -8 72 272
use INVX1  _1956_
timestamp 1701862152
transform -1 0 6370 0 -1 1310
box -12 -8 52 272
use AOI21X1  _1957_
timestamp 1702508443
transform -1 0 6170 0 -1 1310
box -12 -8 92 272
use NAND3X1  _1958_
timestamp 1702508443
transform 1 0 5370 0 -1 1310
box -12 -8 92 272
use INVX1  _1959_
timestamp 1701862152
transform 1 0 5790 0 -1 2870
box -12 -8 52 272
use NOR2X1  _1960_
timestamp 1701862152
transform -1 0 6290 0 -1 2870
box -12 -8 74 272
use OAI21X1  _1961_
timestamp 1702508443
transform -1 0 4570 0 1 2350
box -12 -8 92 272
use NAND3X1  _1962_
timestamp 1702508443
transform 1 0 5970 0 1 2350
box -12 -8 92 272
use NOR2X1  _1963_
timestamp 1701862152
transform 1 0 5430 0 1 1310
box -12 -8 74 272
use INVX2  _1964_
timestamp 1701862152
transform 1 0 9250 0 1 1310
box -12 -8 52 272
use NAND2X1  _1965_
timestamp 1702508443
transform 1 0 7650 0 1 790
box -12 -8 72 272
use NOR2X1  _1966_
timestamp 1701862152
transform -1 0 7790 0 1 270
box -12 -8 74 272
use AND2X2  _1967_
timestamp 1701862152
transform -1 0 6890 0 1 270
box -12 -8 94 272
use AOI22X1  _1968_
timestamp 1701862152
transform 1 0 5610 0 -1 1310
box -14 -8 114 272
use OAI21X1  _1969_
timestamp 1702508443
transform 1 0 5810 0 1 2870
box -12 -8 92 272
use OAI21X1  _1970_
timestamp 1702508443
transform 1 0 5450 0 -1 3390
box -12 -8 92 272
use AND2X2  _1971_
timestamp 1701862152
transform 1 0 5890 0 1 3910
box -12 -8 94 272
use INVX1  _1972_
timestamp 1701862152
transform 1 0 5830 0 1 4950
box -12 -8 52 272
use NOR2X1  _1973_
timestamp 1701862152
transform -1 0 6190 0 -1 3910
box -12 -8 74 272
use OAI21X1  _1974_
timestamp 1702508443
transform 1 0 6350 0 -1 3910
box -12 -8 92 272
use MUX2X1  _1975_
timestamp 1701862152
transform -1 0 6230 0 1 3910
box -12 -8 114 272
use OAI21X1  _1976_
timestamp 1702508443
transform -1 0 6670 0 -1 3910
box -12 -8 92 272
use XOR2X1  _1977_
timestamp 1702508443
transform 1 0 6930 0 1 2870
box -12 -8 132 272
use NOR2X1  _1978_
timestamp 1701862152
transform -1 0 6510 0 -1 2870
box -12 -8 74 272
use INVX1  _1979_
timestamp 1701862152
transform 1 0 6510 0 1 2870
box -12 -8 52 272
use NOR2X1  _1980_
timestamp 1701862152
transform 1 0 6710 0 1 2870
box -12 -8 74 272
use AOI21X1  _1981_
timestamp 1702508443
transform 1 0 6270 0 1 2870
box -12 -8 92 272
use NAND3X1  _1982_
timestamp 1702508443
transform -1 0 5810 0 -1 1830
box -12 -8 92 272
use NOR3X1  _1983_
timestamp 1701862152
transform -1 0 4990 0 -1 270
box -12 -8 172 272
use NOR2X1  _1984_
timestamp 1701862152
transform -1 0 6590 0 -1 1310
box -12 -8 74 272
use AOI22X1  _1985_
timestamp 1701862152
transform 1 0 5110 0 -1 1310
box -14 -8 114 272
use OAI21X1  _1986_
timestamp 1702508443
transform 1 0 8310 0 1 790
box -12 -8 92 272
use NAND2X1  _1987_
timestamp 1702508443
transform 1 0 6990 0 1 1310
box -12 -8 72 272
use INVX1  _1988_
timestamp 1701862152
transform -1 0 7450 0 1 1310
box -12 -8 52 272
use INVX1  _1989_
timestamp 1701862152
transform 1 0 2810 0 -1 5470
box -12 -8 52 272
use OAI21X1  _1990_
timestamp 1702508443
transform 1 0 2130 0 1 1830
box -12 -8 92 272
use OAI21X1  _1991_
timestamp 1702508443
transform -1 0 2910 0 1 1830
box -12 -8 92 272
use OAI21X1  _1992_
timestamp 1702508443
transform -1 0 4310 0 -1 2350
box -12 -8 92 272
use OAI21X1  _1993_
timestamp 1702508443
transform -1 0 4550 0 -1 2350
box -12 -8 92 272
use NAND3X1  _1994_
timestamp 1702508443
transform 1 0 2590 0 1 1830
box -12 -8 92 272
use NAND3X1  _1995_
timestamp 1702508443
transform 1 0 3050 0 1 1830
box -12 -8 92 272
use AOI21X1  _1996_
timestamp 1702508443
transform -1 0 6810 0 1 790
box -12 -8 92 272
use AND2X2  _1997_
timestamp 1701862152
transform -1 0 5150 0 1 790
box -12 -8 94 272
use NAND3X1  _1998_
timestamp 1702508443
transform 1 0 4350 0 1 270
box -12 -8 92 272
use INVX1  _1999_
timestamp 1701862152
transform -1 0 3970 0 -1 270
box -12 -8 52 272
use NOR2X1  _2000_
timestamp 1701862152
transform -1 0 4670 0 -1 270
box -12 -8 74 272
use AND2X2  _2001_
timestamp 1701862152
transform -1 0 6070 0 -1 2870
box -12 -8 94 272
use OAI21X1  _2002_
timestamp 1702508443
transform -1 0 2010 0 1 2870
box -12 -8 92 272
use NOR2X1  _2003_
timestamp 1701862152
transform 1 0 1430 0 -1 3390
box -12 -8 74 272
use AOI21X1  _2004_
timestamp 1702508443
transform 1 0 2870 0 -1 3390
box -12 -8 92 272
use OAI21X1  _2005_
timestamp 1702508443
transform -1 0 3210 0 1 2870
box -12 -8 92 272
use NAND3X1  _2006_
timestamp 1702508443
transform 1 0 2890 0 1 2870
box -12 -8 92 272
use NAND2X1  _2007_
timestamp 1702508443
transform 1 0 6910 0 -1 2870
box -12 -8 72 272
use NAND3X1  _2008_
timestamp 1702508443
transform 1 0 590 0 -1 1830
box -12 -8 92 272
use NOR2X1  _2009_
timestamp 1701862152
transform -1 0 4150 0 -1 3390
box -12 -8 74 272
use OAI21X1  _2010_
timestamp 1702508443
transform -1 0 4450 0 -1 2870
box -12 -8 92 272
use INVX1  _2011_
timestamp 1701862152
transform -1 0 2170 0 1 790
box -12 -8 52 272
use OAI21X1  _2012_
timestamp 1702508443
transform 1 0 1650 0 1 790
box -12 -8 92 272
use OAI21X1  _2013_
timestamp 1702508443
transform -1 0 1970 0 1 790
box -12 -8 92 272
use INVX1  _2014_
timestamp 1701862152
transform 1 0 4570 0 1 1310
box -12 -8 52 272
use OAI21X1  _2015_
timestamp 1702508443
transform 1 0 3290 0 1 1830
box -12 -8 92 272
use OAI21X1  _2016_
timestamp 1702508443
transform -1 0 3850 0 1 1830
box -12 -8 92 272
use OAI21X1  _2017_
timestamp 1702508443
transform -1 0 5350 0 -1 1830
box -12 -8 92 272
use NOR2X1  _2018_
timestamp 1701862152
transform 1 0 5070 0 -1 1830
box -12 -8 74 272
use NAND3X1  _2019_
timestamp 1702508443
transform -1 0 5650 0 -1 2870
box -12 -8 92 272
use AOI21X1  _2020_
timestamp 1702508443
transform -1 0 5410 0 -1 2870
box -12 -8 92 272
use NAND2X1  _2021_
timestamp 1702508443
transform -1 0 7030 0 -1 1310
box -12 -8 72 272
use NAND2X1  _2022_
timestamp 1702508443
transform -1 0 7270 0 1 790
box -12 -8 72 272
use INVX1  _2023_
timestamp 1701862152
transform 1 0 8270 0 1 1830
box -12 -8 52 272
use OAI21X1  _2024_
timestamp 1702508443
transform -1 0 8530 0 1 1830
box -12 -8 92 272
use NOR2X1  _2025_
timestamp 1701862152
transform 1 0 9650 0 -1 790
box -12 -8 74 272
use AOI21X1  _2026_
timestamp 1702508443
transform -1 0 8850 0 1 790
box -12 -8 92 272
use NAND3X1  _2027_
timestamp 1702508443
transform -1 0 7050 0 1 790
box -12 -8 92 272
use INVX1  _2028_
timestamp 1701862152
transform 1 0 7090 0 -1 790
box -12 -8 52 272
use NAND2X1  _2029_
timestamp 1702508443
transform 1 0 7530 0 1 270
box -12 -8 72 272
use NOR2X1  _2030_
timestamp 1701862152
transform -1 0 7250 0 -1 1310
box -12 -8 74 272
use NAND3X1  _2031_
timestamp 1702508443
transform 1 0 7530 0 -1 790
box -12 -8 92 272
use INVX1  _2032_
timestamp 1701862152
transform -1 0 8830 0 1 270
box -12 -8 52 272
use OR2X2  _2033_
timestamp 1702508443
transform 1 0 8310 0 1 1310
box -12 -8 92 272
use NOR2X1  _2034_
timestamp 1701862152
transform -1 0 9030 0 -1 1310
box -12 -8 74 272
use NAND2X1  _2035_
timestamp 1702508443
transform -1 0 8610 0 1 790
box -12 -8 72 272
use NAND2X1  _2036_
timestamp 1702508443
transform -1 0 8770 0 -1 1830
box -12 -8 72 272
use NOR2X1  _2037_
timestamp 1701862152
transform -1 0 8830 0 -1 790
box -12 -8 74 272
use NAND2X1  _2038_
timestamp 1702508443
transform 1 0 8090 0 1 790
box -12 -8 72 272
use OAI21X1  _2039_
timestamp 1702508443
transform 1 0 7850 0 1 790
box -12 -8 92 272
use NOR3X1  _2040_
timestamp 1701862152
transform -1 0 7930 0 -1 790
box -12 -8 172 272
use OAI21X1  _2041_
timestamp 1702508443
transform -1 0 7070 0 -1 270
box -12 -8 92 272
use NAND2X1  _2042_
timestamp 1702508443
transform 1 0 8990 0 -1 790
box -12 -8 72 272
use NOR2X1  _2043_
timestamp 1701862152
transform 1 0 7310 0 1 270
box -12 -8 74 272
use AOI22X1  _2044_
timestamp 1701862152
transform 1 0 7050 0 1 270
box -14 -8 114 272
use AND2X2  _2045_
timestamp 1701862152
transform -1 0 6430 0 1 270
box -12 -8 94 272
use OAI21X1  _2046_
timestamp 1702508443
transform 1 0 6530 0 -1 270
box -12 -8 92 272
use NAND3X1  _2047_
timestamp 1702508443
transform -1 0 6390 0 -1 270
box -12 -8 92 272
use INVX1  _2048_
timestamp 1701862152
transform -1 0 6150 0 -1 270
box -12 -8 52 272
use NAND3X1  _2049_
timestamp 1702508443
transform -1 0 7370 0 -1 790
box -12 -8 92 272
use NOR2X1  _2050_
timestamp 1701862152
transform 1 0 1550 0 -1 2870
box -12 -8 74 272
use INVX1  _2051_
timestamp 1701862152
transform 1 0 6350 0 -1 2350
box -12 -8 52 272
use OAI22X1  _2052_
timestamp 1701862152
transform -1 0 6330 0 1 790
box -12 -8 112 272
use OAI21X1  _2053_
timestamp 1702508443
transform -1 0 4510 0 1 1830
box -12 -8 92 272
use OAI21X1  _2054_
timestamp 1702508443
transform 1 0 2970 0 1 1310
box -12 -8 92 272
use OAI21X1  _2055_
timestamp 1702508443
transform -1 0 3290 0 1 1310
box -12 -8 92 272
use NOR2X1  _2056_
timestamp 1701862152
transform -1 0 1990 0 -1 1310
box -12 -8 74 272
use NAND2X1  _2057_
timestamp 1702508443
transform 1 0 2810 0 1 790
box -12 -8 72 272
use NAND3X1  _2058_
timestamp 1702508443
transform 1 0 3730 0 1 790
box -12 -8 92 272
use NOR2X1  _2059_
timestamp 1701862152
transform 1 0 3970 0 1 790
box -12 -8 74 272
use NAND3X1  _2060_
timestamp 1702508443
transform -1 0 4270 0 1 790
box -12 -8 92 272
use INVX1  _2061_
timestamp 1701862152
transform -1 0 3070 0 -1 270
box -12 -8 52 272
use OR2X2  _2062_
timestamp 1702508443
transform 1 0 2850 0 1 270
box -12 -8 92 272
use OR2X2  _2063_
timestamp 1702508443
transform 1 0 3230 0 -1 270
box -12 -8 92 272
use NOR2X1  _2064_
timestamp 1701862152
transform 1 0 3470 0 -1 270
box -12 -8 74 272
use NAND3X1  _2065_
timestamp 1702508443
transform -1 0 3770 0 -1 270
box -12 -8 92 272
use NOR2X1  _2066_
timestamp 1701862152
transform -1 0 5530 0 -1 270
box -12 -8 74 272
use NOR2X1  _2067_
timestamp 1701862152
transform 1 0 7430 0 1 790
box -12 -8 74 272
use AOI22X1  _2068_
timestamp 1701862152
transform 1 0 5970 0 1 790
box -14 -8 114 272
use OAI21X1  _2069_
timestamp 1702508443
transform 1 0 3470 0 -1 1830
box -12 -8 92 272
use OAI21X1  _2070_
timestamp 1702508443
transform -1 0 4010 0 -1 1830
box -12 -8 92 272
use NAND2X1  _2071_
timestamp 1702508443
transform -1 0 5830 0 1 790
box -12 -8 72 272
use OAI21X1  _2072_
timestamp 1702508443
transform -1 0 7910 0 1 1310
box -12 -8 92 272
use OAI22X1  _2073_
timestamp 1701862152
transform 1 0 6730 0 1 1310
box -12 -8 112 272
use NOR2X1  _2074_
timestamp 1701862152
transform 1 0 1870 0 1 1310
box -12 -8 74 272
use NAND2X1  _2075_
timestamp 1702508443
transform -1 0 2370 0 1 1310
box -12 -8 72 272
use OAI21X1  _2076_
timestamp 1702508443
transform -1 0 2450 0 -1 1310
box -12 -8 92 272
use OR2X2  _2077_
timestamp 1702508443
transform 1 0 4250 0 -1 1310
box -12 -8 92 272
use NAND2X1  _2078_
timestamp 1702508443
transform -1 0 2430 0 1 1830
box -12 -8 72 272
use NAND2X1  _2079_
timestamp 1702508443
transform -1 0 1070 0 -1 1830
box -12 -8 72 272
use OAI21X1  _2080_
timestamp 1702508443
transform 1 0 2350 0 -1 1830
box -12 -8 92 272
use INVX1  _2081_
timestamp 1701862152
transform 1 0 2590 0 -1 1830
box -12 -8 52 272
use AOI22X1  _2082_
timestamp 1701862152
transform -1 0 2890 0 -1 1830
box -14 -8 114 272
use NOR2X1  _2083_
timestamp 1701862152
transform 1 0 4470 0 -1 1310
box -12 -8 74 272
use NAND3X1  _2084_
timestamp 1702508443
transform -1 0 5390 0 1 790
box -12 -8 92 272
use NOR3X1  _2085_
timestamp 1701862152
transform -1 0 5310 0 -1 270
box -12 -8 172 272
use NAND3X1  _2086_
timestamp 1702508443
transform -1 0 4450 0 -1 270
box -12 -8 92 272
use NAND2X1  _2087_
timestamp 1702508443
transform -1 0 4910 0 1 790
box -12 -8 72 272
use INVX1  _2088_
timestamp 1701862152
transform -1 0 5730 0 1 270
box -12 -8 52 272
use NOR2X1  _2089_
timestamp 1701862152
transform 1 0 5470 0 1 270
box -12 -8 74 272
use NAND2X1  _2090_
timestamp 1702508443
transform -1 0 5070 0 -1 790
box -12 -8 72 272
use NAND2X1  _2091_
timestamp 1702508443
transform 1 0 3270 0 1 790
box -12 -8 72 272
use NOR2X1  _2092_
timestamp 1701862152
transform 1 0 2830 0 -1 270
box -12 -8 74 272
use NAND3X1  _2093_
timestamp 1702508443
transform -1 0 3050 0 -1 790
box -12 -8 92 272
use INVX1  _2094_
timestamp 1701862152
transform 1 0 2390 0 -1 270
box -12 -8 52 272
use NAND3X1  _2095_
timestamp 1702508443
transform 1 0 2590 0 -1 270
box -12 -8 92 272
use NOR2X1  _2096_
timestamp 1701862152
transform -1 0 5090 0 1 270
box -12 -8 74 272
use NAND3X1  _2097_
timestamp 1702508443
transform -1 0 5310 0 1 270
box -12 -8 92 272
use NOR2X1  _2098_
timestamp 1701862152
transform 1 0 4810 0 1 270
box -12 -8 74 272
use OAI21X1  _2099_
timestamp 1702508443
transform 1 0 4130 0 -1 270
box -12 -8 92 272
use NAND2X1  _2100_
timestamp 1702508443
transform -1 0 6030 0 -1 1830
box -12 -8 72 272
use INVX1  _2101_
timestamp 1701862152
transform -1 0 5930 0 1 1310
box -12 -8 52 272
use OAI21X1  _2102_
timestamp 1702508443
transform -1 0 6370 0 1 1310
box -12 -8 92 272
use NAND2X1  _2103_
timestamp 1702508443
transform 1 0 5870 0 -1 1310
box -12 -8 72 272
use NOR2X1  _2104_
timestamp 1701862152
transform -1 0 6130 0 1 1310
box -12 -8 74 272
use NOR2X1  _2105_
timestamp 1701862152
transform -1 0 4450 0 -1 1830
box -12 -8 74 272
use NAND3X1  _2106_
timestamp 1702508443
transform 1 0 4090 0 -1 790
box -12 -8 92 272
use NAND2X1  _2107_
timestamp 1702508443
transform -1 0 3710 0 -1 790
box -12 -8 72 272
use NAND3X1  _2108_
timestamp 1702508443
transform 1 0 3030 0 1 790
box -12 -8 92 272
use NOR2X1  _2109_
timestamp 1701862152
transform -1 0 3490 0 -1 790
box -12 -8 74 272
use NAND2X1  _2110_
timestamp 1702508443
transform 1 0 3210 0 -1 790
box -12 -8 72 272
use NOR2X1  _2111_
timestamp 1701862152
transform -1 0 3930 0 -1 790
box -12 -8 74 272
use NAND3X1  _2112_
timestamp 1702508443
transform -1 0 5290 0 -1 790
box -12 -8 92 272
use NOR2X1  _2113_
timestamp 1701862152
transform -1 0 5270 0 1 1310
box -12 -8 74 272
use NAND3X1  _2114_
timestamp 1702508443
transform -1 0 5730 0 1 1310
box -12 -8 92 272
use AND2X2  _2115_
timestamp 1701862152
transform -1 0 5770 0 -1 790
box -12 -8 94 272
use INVX1  _2116_
timestamp 1701862152
transform 1 0 2530 0 1 1310
box -12 -8 52 272
use OAI21X1  _2117_
timestamp 1702508443
transform 1 0 2730 0 1 1310
box -12 -8 92 272
use NAND3X1  _2118_
timestamp 1702508443
transform 1 0 3910 0 1 1310
box -12 -8 92 272
use NOR2X1  _2119_
timestamp 1701862152
transform -1 0 4190 0 1 1310
box -12 -8 74 272
use NAND2X1  _2120_
timestamp 1702508443
transform 1 0 4030 0 -1 1310
box -12 -8 72 272
use NOR2X1  _2121_
timestamp 1701862152
transform -1 0 4650 0 1 270
box -12 -8 74 272
use INVX1  _2122_
timestamp 1701862152
transform -1 0 2970 0 1 2350
box -12 -8 52 272
use NOR2X1  _2123_
timestamp 1701862152
transform 1 0 2890 0 -1 2350
box -12 -8 74 272
use NAND3X1  _2124_
timestamp 1702508443
transform -1 0 3850 0 -1 2350
box -12 -8 92 272
use OAI21X1  _2125_
timestamp 1702508443
transform 1 0 5910 0 -1 3390
box -12 -8 92 272
use OAI21X1  _2126_
timestamp 1702508443
transform 1 0 5570 0 1 2870
box -12 -8 92 272
use AOI21X1  _2127_
timestamp 1702508443
transform -1 0 6130 0 1 2870
box -12 -8 92 272
use NOR2X1  _2128_
timestamp 1701862152
transform 1 0 4690 0 1 2870
box -12 -8 74 272
use NAND2X1  _2129_
timestamp 1702508443
transform 1 0 5370 0 1 2870
box -12 -8 72 272
use NOR2X1  _2130_
timestamp 1701862152
transform -1 0 4770 0 -1 2350
box -12 -8 74 272
use NAND2X1  _2131_
timestamp 1702508443
transform 1 0 4770 0 1 1310
box -12 -8 72 272
use NOR2X1  _2132_
timestamp 1701862152
transform -1 0 4690 0 1 790
box -12 -8 74 272
use NAND3X1  _2133_
timestamp 1702508443
transform 1 0 4550 0 -1 790
box -12 -8 92 272
use OAI21X1  _2134_
timestamp 1702508443
transform 1 0 3690 0 -1 2870
box -12 -8 92 272
use OAI21X1  _2135_
timestamp 1702508443
transform 1 0 4310 0 -1 3390
box -12 -8 92 272
use INVX1  _2136_
timestamp 1701862152
transform -1 0 2870 0 1 3390
box -12 -8 52 272
use NAND3X1  _2137_
timestamp 1702508443
transform 1 0 2410 0 1 3390
box -12 -8 92 272
use OAI21X1  _2138_
timestamp 1702508443
transform 1 0 3210 0 -1 4430
box -12 -8 92 272
use OAI21X1  _2139_
timestamp 1702508443
transform -1 0 3050 0 -1 4430
box -12 -8 92 272
use NOR2X1  _2140_
timestamp 1701862152
transform 1 0 2910 0 1 4430
box -12 -8 74 272
use NAND2X1  _2141_
timestamp 1702508443
transform -1 0 3170 0 1 4430
box -12 -8 72 272
use NOR2X1  _2142_
timestamp 1701862152
transform 1 0 3030 0 1 3390
box -12 -8 74 272
use INVX1  _2143_
timestamp 1701862152
transform -1 0 7550 0 -1 3390
box -12 -8 52 272
use OAI21X1  _2144_
timestamp 1702508443
transform 1 0 2170 0 1 2870
box -12 -8 92 272
use INVX1  _2145_
timestamp 1701862152
transform -1 0 10170 0 -1 2870
box -12 -8 52 272
use AOI21X1  _2146_
timestamp 1702508443
transform -1 0 7790 0 -1 3390
box -12 -8 92 272
use INVX1  _2147_
timestamp 1701862152
transform 1 0 7690 0 -1 3910
box -12 -8 52 272
use NAND2X1  _2148_
timestamp 1702508443
transform 1 0 7510 0 1 3390
box -12 -8 72 272
use OAI21X1  _2149_
timestamp 1702508443
transform 1 0 7730 0 1 3390
box -12 -8 92 272
use OAI21X1  _2150_
timestamp 1702508443
transform -1 0 8050 0 1 3390
box -12 -8 92 272
use OAI21X1  _2151_
timestamp 1702508443
transform 1 0 7270 0 -1 3390
box -12 -8 92 272
use OAI21X1  _2152_
timestamp 1702508443
transform 1 0 7030 0 -1 3390
box -12 -8 92 272
use NAND3X1  _2153_
timestamp 1702508443
transform -1 0 6230 0 -1 3390
box -12 -8 92 272
use INVX2  _2154_
timestamp 1701862152
transform 1 0 2930 0 -1 7030
box -12 -8 52 272
use INVX2  _2155_
timestamp 1701862152
transform 1 0 6470 0 1 5990
box -12 -8 52 272
use OAI21X1  _2156_
timestamp 1702508443
transform -1 0 4770 0 1 3910
box -12 -8 92 272
use NOR2X1  _2157_
timestamp 1701862152
transform -1 0 4890 0 -1 4430
box -12 -8 74 272
use OAI21X1  _2158_
timestamp 1702508443
transform -1 0 2770 0 1 2350
box -12 -8 92 272
use OAI21X1  _2159_
timestamp 1702508443
transform 1 0 3610 0 1 3910
box -12 -8 92 272
use NOR2X1  _2160_
timestamp 1701862152
transform -1 0 3970 0 -1 4430
box -12 -8 74 272
use INVX1  _2161_
timestamp 1701862152
transform -1 0 4090 0 1 3910
box -12 -8 52 272
use INVX1  _2162_
timestamp 1701862152
transform -1 0 4530 0 1 3910
box -12 -8 52 272
use OAI21X1  _2163_
timestamp 1702508443
transform 1 0 3810 0 -1 3910
box -12 -8 92 272
use INVX2  _2164_
timestamp 1701862152
transform -1 0 670 0 -1 4950
box -12 -8 52 272
use OAI22X1  _2165_
timestamp 1701862152
transform -1 0 3430 0 -1 3910
box -12 -8 112 272
use NOR2X1  _2166_
timestamp 1701862152
transform 1 0 4050 0 -1 3910
box -12 -8 74 272
use NAND3X1  _2167_
timestamp 1702508443
transform 1 0 4250 0 1 3910
box -12 -8 92 272
use NAND2X1  _2168_
timestamp 1702508443
transform 1 0 3170 0 1 3910
box -12 -8 72 272
use OAI21X1  _2169_
timestamp 1702508443
transform 1 0 2530 0 -1 4430
box -12 -8 92 272
use NOR2X1  _2170_
timestamp 1701862152
transform -1 0 2810 0 -1 4430
box -12 -8 74 272
use NAND3X1  _2171_
timestamp 1702508443
transform 1 0 4130 0 -1 4430
box -12 -8 92 272
use NOR2X1  _2172_
timestamp 1701862152
transform 1 0 4370 0 -1 4430
box -12 -8 74 272
use NAND3X1  _2173_
timestamp 1702508443
transform -1 0 4670 0 -1 4430
box -12 -8 92 272
use OAI22X1  _2174_
timestamp 1701862152
transform 1 0 6110 0 1 7030
box -12 -8 112 272
use INVX2  _2175_
timestamp 1701862152
transform -1 0 2630 0 1 8070
box -12 -8 52 272
use INVX2  _2176_
timestamp 1701862152
transform -1 0 6550 0 -1 8070
box -12 -8 52 272
use OAI22X1  _2177_
timestamp 1701862152
transform 1 0 5030 0 1 8070
box -12 -8 112 272
use INVX1  _2178_
timestamp 1701862152
transform -1 0 4250 0 -1 8590
box -12 -8 52 272
use OAI22X1  _2179_
timestamp 1701862152
transform -1 0 6130 0 -1 8070
box -12 -8 112 272
use INVX2  _2180_
timestamp 1701862152
transform -1 0 3090 0 -1 9630
box -12 -8 52 272
use INVX2  _2181_
timestamp 1701862152
transform 1 0 5130 0 1 7550
box -12 -8 52 272
use OAI22X1  _2182_
timestamp 1701862152
transform 1 0 5650 0 -1 10150
box -12 -8 112 272
use INVX1  _2183_
timestamp 1701862152
transform -1 0 3650 0 1 10150
box -12 -8 52 272
use INVX1  _2184_
timestamp 1701862152
transform 1 0 4430 0 1 8070
box -12 -8 52 272
use OAI22X1  _2185_
timestamp 1701862152
transform 1 0 6050 0 1 10150
box -12 -8 112 272
use INVX2  _2186_
timestamp 1701862152
transform 1 0 3610 0 1 10670
box -12 -8 52 272
use OAI22X1  _2187_
timestamp 1701862152
transform -1 0 5610 0 -1 10670
box -12 -8 112 272
use INVX2  _2188_
timestamp 1701862152
transform 1 0 2210 0 -1 10670
box -12 -8 52 272
use OAI22X1  _2189_
timestamp 1701862152
transform 1 0 5770 0 -1 10670
box -12 -8 112 272
use INVX1  _2190_
timestamp 1701862152
transform -1 0 2950 0 1 10150
box -12 -8 52 272
use OAI22X1  _2191_
timestamp 1701862152
transform -1 0 5490 0 -1 10150
box -12 -8 112 272
use INVX1  _2192_
timestamp 1701862152
transform -1 0 11210 0 1 3910
box -12 -8 52 272
use OAI21X1  _2193_
timestamp 1702508443
transform 1 0 1330 0 -1 3910
box -12 -8 92 272
use INVX1  _2194_
timestamp 1701862152
transform 1 0 1130 0 -1 3910
box -12 -8 52 272
use NAND3X1  _2195_
timestamp 1702508443
transform 1 0 2710 0 1 3910
box -12 -8 92 272
use NOR2X1  _2196_
timestamp 1701862152
transform 1 0 2950 0 1 3910
box -12 -8 74 272
use OAI21X1  _2197_
timestamp 1702508443
transform 1 0 5430 0 1 3910
box -12 -8 92 272
use NOR2X1  _2198_
timestamp 1701862152
transform 1 0 370 0 1 1830
box -12 -8 74 272
use NAND2X1  _2199_
timestamp 1702508443
transform -1 0 2950 0 -1 3910
box -12 -8 72 272
use NAND3X1  _2200_
timestamp 1702508443
transform 1 0 5450 0 -1 3910
box -12 -8 92 272
use NOR2X1  _2201_
timestamp 1701862152
transform -1 0 5730 0 1 3910
box -12 -8 74 272
use INVX4  _2202_
timestamp 1701862152
transform -1 0 8310 0 -1 4430
box -12 -8 72 272
use OAI21X1  _2203_
timestamp 1702508443
transform -1 0 5050 0 -1 3910
box -12 -8 92 272
use OAI21X1  _2204_
timestamp 1702508443
transform 1 0 5210 0 -1 3910
box -12 -8 92 272
use NOR3X1  _2205_
timestamp 1701862152
transform -1 0 9210 0 -1 3910
box -12 -8 172 272
use NAND3X1  _2206_
timestamp 1702508443
transform 1 0 9130 0 1 3910
box -12 -8 92 272
use OR2X2  _2207_
timestamp 1702508443
transform 1 0 9610 0 -1 3910
box -12 -8 92 272
use AOI21X1  _2208_
timestamp 1702508443
transform -1 0 9930 0 -1 3910
box -12 -8 92 272
use OAI21X1  _2209_
timestamp 1702508443
transform -1 0 9730 0 1 4430
box -12 -8 92 272
use INVX2  _2210_
timestamp 1701862152
transform -1 0 10690 0 -1 4950
box -12 -8 52 272
use OAI21X1  _2211_
timestamp 1702508443
transform 1 0 9370 0 -1 3910
box -12 -8 92 272
use NAND2X1  _2212_
timestamp 1702508443
transform -1 0 8990 0 1 3910
box -12 -8 72 272
use AOI21X1  _2213_
timestamp 1702508443
transform -1 0 9450 0 1 3910
box -12 -8 92 272
use NAND3X1  _2214_
timestamp 1702508443
transform -1 0 9630 0 -1 4430
box -12 -8 92 272
use OAI21X1  _2215_
timestamp 1702508443
transform 1 0 9790 0 -1 4430
box -12 -8 92 272
use NAND3X1  _2216_
timestamp 1702508443
transform -1 0 9610 0 -1 7030
box -12 -8 92 272
use AND2X2  _2217_
timestamp 1701862152
transform 1 0 9330 0 -1 4430
box -12 -8 94 272
use INVX1  _2218_
timestamp 1701862152
transform -1 0 9870 0 1 3910
box -12 -8 52 272
use OR2X2  _2219_
timestamp 1702508443
transform 1 0 10030 0 1 3910
box -12 -8 92 272
use AOI21X1  _2220_
timestamp 1702508443
transform 1 0 10410 0 -1 4950
box -12 -8 92 272
use NAND2X1  _2221_
timestamp 1702508443
transform -1 0 9810 0 -1 7030
box -12 -8 72 272
use OR2X2  _2222_
timestamp 1702508443
transform 1 0 10150 0 1 4430
box -12 -8 92 272
use OR2X2  _2223_
timestamp 1702508443
transform -1 0 10110 0 -1 4430
box -12 -8 92 272
use AOI22X1  _2224_
timestamp 1701862152
transform -1 0 9990 0 1 4430
box -14 -8 114 272
use AOI22X1  _2225_
timestamp 1701862152
transform 1 0 10150 0 -1 4950
box -14 -8 114 272
use AOI22X1  _2226_
timestamp 1701862152
transform 1 0 9030 0 -1 7030
box -14 -8 114 272
use NAND3X1  _2227_
timestamp 1702508443
transform -1 0 9370 0 -1 7030
box -12 -8 92 272
use INVX1  _2228_
timestamp 1701862152
transform -1 0 5850 0 -1 7030
box -12 -8 52 272
use OAI21X1  _2229_
timestamp 1702508443
transform 1 0 4410 0 1 3390
box -12 -8 92 272
use OR2X2  _2230_
timestamp 1702508443
transform -1 0 4570 0 -1 3910
box -12 -8 92 272
use NOR2X1  _2231_
timestamp 1701862152
transform -1 0 4330 0 -1 3910
box -12 -8 74 272
use OAI21X1  _2232_
timestamp 1702508443
transform 1 0 1690 0 1 2870
box -12 -8 92 272
use AOI21X1  _2233_
timestamp 1702508443
transform 1 0 2410 0 1 2870
box -12 -8 92 272
use AND2X2  _2234_
timestamp 1701862152
transform -1 0 2730 0 1 2870
box -12 -8 94 272
use INVX1  _2235_
timestamp 1701862152
transform 1 0 6410 0 1 3390
box -12 -8 52 272
use AOI21X1  _2236_
timestamp 1702508443
transform -1 0 5770 0 -1 3910
box -12 -8 92 272
use NAND3X1  _2237_
timestamp 1702508443
transform -1 0 4810 0 -1 3910
box -12 -8 92 272
use INVX2  _2238_
timestamp 1701862152
transform 1 0 4810 0 -1 4950
box -12 -8 52 272
use NOR2X1  _2239_
timestamp 1701862152
transform 1 0 2930 0 1 4950
box -12 -8 74 272
use NAND2X1  _2240_
timestamp 1702508443
transform 1 0 2490 0 1 3910
box -12 -8 72 272
use OAI21X1  _2241_
timestamp 1702508443
transform -1 0 2570 0 1 4950
box -12 -8 92 272
use OAI21X1  _2242_
timestamp 1702508443
transform 1 0 2550 0 -1 4950
box -12 -8 92 272
use NOR2X1  _2243_
timestamp 1701862152
transform 1 0 2710 0 1 4950
box -12 -8 74 272
use NAND3X1  _2244_
timestamp 1702508443
transform 1 0 3150 0 1 4950
box -12 -8 92 272
use INVX1  _2245_
timestamp 1701862152
transform 1 0 2990 0 1 5990
box -12 -8 52 272
use AOI21X1  _2246_
timestamp 1702508443
transform 1 0 3010 0 -1 4950
box -12 -8 92 272
use OAI22X1  _2247_
timestamp 1701862152
transform -1 0 3210 0 -1 6510
box -12 -8 112 272
use AOI21X1  _2248_
timestamp 1702508443
transform 1 0 3590 0 -1 7030
box -12 -8 92 272
use OAI21X1  _2249_
timestamp 1702508443
transform 1 0 6370 0 1 7030
box -12 -8 92 272
use NAND2X1  _2250_
timestamp 1702508443
transform -1 0 10690 0 -1 7550
box -12 -8 72 272
use AOI22X1  _2251_
timestamp 1701862152
transform -1 0 10810 0 1 8070
box -14 -8 114 272
use NAND3X1  _2252_
timestamp 1702508443
transform -1 0 11090 0 -1 8070
box -12 -8 92 272
use NAND3X1  _2253_
timestamp 1702508443
transform -1 0 10850 0 -1 8070
box -12 -8 92 272
use INVX1  _2254_
timestamp 1701862152
transform 1 0 5490 0 1 8070
box -12 -8 52 272
use NAND2X1  _2255_
timestamp 1702508443
transform 1 0 3110 0 1 7030
box -12 -8 72 272
use OAI21X1  _2256_
timestamp 1702508443
transform -1 0 5290 0 1 7030
box -12 -8 92 272
use AOI21X1  _2257_
timestamp 1702508443
transform 1 0 5150 0 -1 7550
box -12 -8 92 272
use OAI21X1  _2258_
timestamp 1702508443
transform 1 0 5810 0 -1 8590
box -12 -8 92 272
use NAND2X1  _2259_
timestamp 1702508443
transform 1 0 10430 0 -1 7550
box -12 -8 72 272
use AOI22X1  _2260_
timestamp 1701862152
transform 1 0 10010 0 1 8070
box -14 -8 114 272
use NAND3X1  _2261_
timestamp 1702508443
transform -1 0 10370 0 1 7550
box -12 -8 92 272
use NAND3X1  _2262_
timestamp 1702508443
transform -1 0 10130 0 1 7550
box -12 -8 92 272
use INVX1  _2263_
timestamp 1701862152
transform 1 0 5570 0 1 7550
box -12 -8 52 272
use INVX1  _2264_
timestamp 1701862152
transform 1 0 1710 0 -1 6510
box -12 -8 52 272
use NOR2X1  _2265_
timestamp 1701862152
transform 1 0 1910 0 -1 6510
box -12 -8 74 272
use INVX1  _2266_
timestamp 1701862152
transform 1 0 4010 0 1 6510
box -12 -8 52 272
use OAI21X1  _2267_
timestamp 1702508443
transform -1 0 3830 0 -1 7550
box -12 -8 92 272
use AOI21X1  _2268_
timestamp 1702508443
transform 1 0 4450 0 -1 7550
box -12 -8 92 272
use OAI21X1  _2269_
timestamp 1702508443
transform 1 0 5770 0 1 7550
box -12 -8 92 272
use NAND2X1  _2270_
timestamp 1702508443
transform 1 0 8690 0 1 7550
box -12 -8 72 272
use AOI22X1  _2271_
timestamp 1701862152
transform -1 0 9050 0 -1 8070
box -14 -8 114 272
use NAND3X1  _2272_
timestamp 1702508443
transform -1 0 9270 0 -1 8070
box -12 -8 92 272
use NAND3X1  _2273_
timestamp 1702508443
transform -1 0 8790 0 -1 8070
box -12 -8 92 272
use INVX1  _2274_
timestamp 1701862152
transform -1 0 6110 0 -1 9630
box -12 -8 52 272
use NAND2X1  _2275_
timestamp 1702508443
transform -1 0 2430 0 1 8070
box -12 -8 72 272
use OAI21X1  _2276_
timestamp 1702508443
transform -1 0 3330 0 1 8070
box -12 -8 92 272
use AOI21X1  _2277_
timestamp 1702508443
transform -1 0 3810 0 -1 8590
box -12 -8 92 272
use OAI21X1  _2278_
timestamp 1702508443
transform 1 0 6650 0 1 9110
box -12 -8 92 272
use NAND2X1  _2279_
timestamp 1702508443
transform -1 0 10370 0 1 5990
box -12 -8 72 272
use AOI22X1  _2280_
timestamp 1701862152
transform 1 0 10530 0 1 5990
box -14 -8 114 272
use NAND3X1  _2281_
timestamp 1702508443
transform -1 0 10870 0 -1 5990
box -12 -8 92 272
use NAND3X1  _2282_
timestamp 1702508443
transform -1 0 10650 0 -1 6510
box -12 -8 92 272
use INVX1  _2283_
timestamp 1701862152
transform 1 0 6050 0 -1 8590
box -12 -8 52 272
use NAND2X1  _2284_
timestamp 1702508443
transform -1 0 2210 0 1 8070
box -12 -8 72 272
use OAI21X1  _2285_
timestamp 1702508443
transform -1 0 4290 0 1 8070
box -12 -8 92 272
use AOI21X1  _2286_
timestamp 1702508443
transform 1 0 5110 0 -1 8590
box -12 -8 92 272
use OAI21X1  _2287_
timestamp 1702508443
transform -1 0 6270 0 1 8590
box -12 -8 92 272
use NAND2X1  _2288_
timestamp 1702508443
transform -1 0 8970 0 1 7550
box -12 -8 72 272
use AOI22X1  _2289_
timestamp 1701862152
transform 1 0 8590 0 1 8070
box -14 -8 114 272
use NAND3X1  _2290_
timestamp 1702508443
transform -1 0 10150 0 -1 8070
box -12 -8 92 272
use NAND3X1  _2291_
timestamp 1702508443
transform -1 0 8930 0 1 8070
box -12 -8 92 272
use INVX1  _2292_
timestamp 1701862152
transform -1 0 6330 0 -1 9110
box -12 -8 52 272
use NAND2X1  _2293_
timestamp 1702508443
transform -1 0 2670 0 -1 8590
box -12 -8 72 272
use OAI21X1  _2294_
timestamp 1702508443
transform -1 0 4150 0 1 8590
box -12 -8 92 272
use AOI21X1  _2295_
timestamp 1702508443
transform 1 0 5030 0 1 8590
box -12 -8 92 272
use OAI21X1  _2296_
timestamp 1702508443
transform 1 0 6750 0 -1 9110
box -12 -8 92 272
use NAND2X1  _2297_
timestamp 1702508443
transform -1 0 9690 0 -1 5990
box -12 -8 72 272
use AOI22X1  _2298_
timestamp 1701862152
transform -1 0 10170 0 -1 5470
box -14 -8 114 272
use NAND3X1  _2299_
timestamp 1702508443
transform -1 0 9490 0 -1 6510
box -12 -8 92 272
use NAND3X1  _2300_
timestamp 1702508443
transform 1 0 9630 0 1 5990
box -12 -8 92 272
use INVX1  _2301_
timestamp 1701862152
transform 1 0 5650 0 1 9630
box -12 -8 52 272
use INVX1  _2302_
timestamp 1701862152
transform -1 0 3590 0 -1 9110
box -12 -8 52 272
use NOR2X1  _2303_
timestamp 1701862152
transform 1 0 2690 0 1 9110
box -12 -8 74 272
use INVX1  _2304_
timestamp 1701862152
transform 1 0 2890 0 -1 9110
box -12 -8 52 272
use OAI21X1  _2305_
timestamp 1702508443
transform -1 0 3930 0 1 8590
box -12 -8 92 272
use AOI21X1  _2306_
timestamp 1702508443
transform 1 0 4550 0 1 8590
box -12 -8 92 272
use OAI21X1  _2307_
timestamp 1702508443
transform 1 0 6410 0 1 9110
box -12 -8 92 272
use NAND2X1  _2308_
timestamp 1702508443
transform -1 0 9010 0 -1 6510
box -12 -8 72 272
use AOI22X1  _2309_
timestamp 1701862152
transform -1 0 8770 0 1 5990
box -14 -8 114 272
use NAND3X1  _2310_
timestamp 1702508443
transform -1 0 9250 0 -1 6510
box -12 -8 92 272
use NAND3X1  _2311_
timestamp 1702508443
transform -1 0 8810 0 -1 6510
box -12 -8 92 272
use INVX1  _2312_
timestamp 1701862152
transform -1 0 5670 0 -1 9630
box -12 -8 52 272
use INVX1  _2313_
timestamp 1701862152
transform -1 0 1950 0 1 8590
box -12 -8 52 272
use NOR2X1  _2314_
timestamp 1701862152
transform 1 0 1530 0 -1 8590
box -12 -8 74 272
use INVX1  _2315_
timestamp 1701862152
transform 1 0 1950 0 -1 8590
box -12 -8 52 272
use OAI21X1  _2316_
timestamp 1702508443
transform -1 0 4390 0 1 8590
box -12 -8 92 272
use AOI21X1  _2317_
timestamp 1702508443
transform 1 0 4790 0 1 8590
box -12 -8 92 272
use OAI21X1  _2318_
timestamp 1702508443
transform 1 0 6890 0 1 9110
box -12 -8 92 272
use INVX1  _2319_
timestamp 1701862152
transform -1 0 11230 0 1 4430
box -12 -8 52 272
use OAI21X1  _2320_
timestamp 1702508443
transform 1 0 5190 0 1 3910
box -12 -8 92 272
use INVX2  _2321_
timestamp 1701862152
transform 1 0 6610 0 1 3910
box -12 -8 52 272
use NAND3X1  _2322_
timestamp 1702508443
transform -1 0 8050 0 1 3910
box -12 -8 92 272
use OAI21X1  _2323_
timestamp 1702508443
transform 1 0 8010 0 -1 4430
box -12 -8 92 272
use INVX1  _2324_
timestamp 1701862152
transform -1 0 11270 0 -1 2870
box -12 -8 52 272
use OAI21X1  _2325_
timestamp 1702508443
transform -1 0 8290 0 1 3910
box -12 -8 92 272
use INVX1  _2326_
timestamp 1701862152
transform -1 0 3290 0 -1 4950
box -12 -8 52 272
use OAI21X1  _2327_
timestamp 1702508443
transform -1 0 3530 0 -1 4950
box -12 -8 92 272
use INVX2  _2328_
timestamp 1701862152
transform 1 0 3950 0 -1 5470
box -12 -8 52 272
use OAI21X1  _2329_
timestamp 1702508443
transform 1 0 3710 0 -1 5470
box -12 -8 92 272
use NOR2X1  _2330_
timestamp 1701862152
transform 1 0 3830 0 1 4950
box -12 -8 74 272
use AOI22X1  _2331_
timestamp 1701862152
transform 1 0 4930 0 1 3910
box -14 -8 114 272
use NAND2X1  _2332_
timestamp 1702508443
transform -1 0 4310 0 1 4950
box -12 -8 72 272
use INVX1  _2333_
timestamp 1701862152
transform -1 0 11250 0 -1 4430
box -12 -8 52 272
use NOR2X1  _2334_
timestamp 1701862152
transform 1 0 9110 0 -1 4430
box -12 -8 74 272
use OAI21X1  _2335_
timestamp 1702508443
transform 1 0 5290 0 -1 5470
box -12 -8 92 272
use INVX1  _2336_
timestamp 1701862152
transform -1 0 5170 0 1 5990
box -12 -8 52 272
use INVX1  _2337_
timestamp 1701862152
transform 1 0 4630 0 1 3390
box -12 -8 52 272
use OAI21X1  _2338_
timestamp 1702508443
transform 1 0 3250 0 1 3390
box -12 -8 92 272
use OAI21X1  _2339_
timestamp 1702508443
transform 1 0 4830 0 1 3390
box -12 -8 92 272
use NAND2X1  _2340_
timestamp 1702508443
transform 1 0 5070 0 1 3390
box -12 -8 72 272
use INVX1  _2341_
timestamp 1701862152
transform -1 0 670 0 1 5990
box -12 -8 52 272
use OAI21X1  _2342_
timestamp 1702508443
transform 1 0 2750 0 1 5470
box -12 -8 92 272
use INVX2  _2343_
timestamp 1701862152
transform -1 0 4710 0 1 6510
box -12 -8 52 272
use OAI21X1  _2344_
timestamp 1702508443
transform -1 0 5010 0 1 5470
box -12 -8 92 272
use INVX1  _2345_
timestamp 1701862152
transform -1 0 4790 0 1 5470
box -12 -8 52 272
use OAI21X1  _2346_
timestamp 1702508443
transform -1 0 4990 0 -1 5990
box -12 -8 92 272
use NAND2X1  _2347_
timestamp 1702508443
transform -1 0 5830 0 -1 5990
box -12 -8 72 272
use OAI21X1  _2348_
timestamp 1702508443
transform 1 0 5350 0 -1 6510
box -12 -8 92 272
use AOI21X1  _2349_
timestamp 1702508443
transform -1 0 5190 0 -1 6510
box -12 -8 92 272
use OAI21X1  _2350_
timestamp 1702508443
transform -1 0 4610 0 -1 6510
box -12 -8 92 272
use INVX1  _2351_
timestamp 1701862152
transform 1 0 5690 0 1 7030
box -12 -8 52 272
use OAI21X1  _2352_
timestamp 1702508443
transform -1 0 5950 0 1 7030
box -12 -8 92 272
use INVX1  _2353_
timestamp 1701862152
transform -1 0 870 0 1 7030
box -12 -8 52 272
use NAND2X1  _2354_
timestamp 1702508443
transform 1 0 5550 0 -1 5990
box -12 -8 72 272
use OAI21X1  _2355_
timestamp 1702508443
transform 1 0 5450 0 1 7030
box -12 -8 92 272
use AOI21X1  _2356_
timestamp 1702508443
transform -1 0 5010 0 -1 7550
box -12 -8 92 272
use OAI21X1  _2357_
timestamp 1702508443
transform 1 0 4810 0 1 8070
box -12 -8 92 272
use INVX1  _2358_
timestamp 1701862152
transform 1 0 5290 0 1 8070
box -12 -8 52 272
use OAI21X1  _2359_
timestamp 1702508443
transform -1 0 5650 0 -1 8590
box -12 -8 92 272
use INVX1  _2360_
timestamp 1701862152
transform -1 0 870 0 -1 6510
box -12 -8 52 272
use NAND2X1  _2361_
timestamp 1702508443
transform -1 0 5390 0 1 5990
box -12 -8 72 272
use OAI21X1  _2362_
timestamp 1702508443
transform 1 0 5350 0 1 6510
box -12 -8 92 272
use AOI21X1  _2363_
timestamp 1702508443
transform 1 0 5370 0 -1 7030
box -12 -8 92 272
use OAI21X1  _2364_
timestamp 1702508443
transform 1 0 5370 0 -1 8070
box -12 -8 92 272
use INVX1  _2365_
timestamp 1701862152
transform 1 0 5610 0 -1 8070
box -12 -8 52 272
use OAI21X1  _2366_
timestamp 1702508443
transform -1 0 5870 0 -1 8070
box -12 -8 92 272
use INVX1  _2367_
timestamp 1701862152
transform 1 0 2790 0 -1 7550
box -12 -8 52 272
use NAND2X1  _2368_
timestamp 1702508443
transform -1 0 5670 0 -1 7030
box -12 -8 72 272
use OAI21X1  _2369_
timestamp 1702508443
transform 1 0 5330 0 1 7550
box -12 -8 92 272
use AOI21X1  _2370_
timestamp 1702508443
transform -1 0 5430 0 -1 8590
box -12 -8 92 272
use OAI21X1  _2371_
timestamp 1702508443
transform 1 0 6050 0 -1 9110
box -12 -8 92 272
use INVX1  _2372_
timestamp 1701862152
transform 1 0 6210 0 1 9110
box -12 -8 52 272
use OAI21X1  _2373_
timestamp 1702508443
transform -1 0 6350 0 -1 9630
box -12 -8 92 272
use INVX1  _2374_
timestamp 1701862152
transform 1 0 150 0 -1 9110
box -12 -8 52 272
use OAI21X1  _2375_
timestamp 1702508443
transform -1 0 4370 0 1 5470
box -12 -8 92 272
use OAI22X1  _2376_
timestamp 1701862152
transform 1 0 4650 0 -1 5990
box -12 -8 112 272
use AOI21X1  _2377_
timestamp 1702508443
transform -1 0 4130 0 -1 6510
box -12 -8 92 272
use OAI21X1  _2378_
timestamp 1702508443
transform 1 0 3810 0 -1 6510
box -12 -8 92 272
use AOI21X1  _2379_
timestamp 1702508443
transform -1 0 5190 0 1 6510
box -12 -8 92 272
use OAI21X1  _2380_
timestamp 1702508443
transform -1 0 4970 0 -1 8590
box -12 -8 92 272
use AOI22X1  _2381_
timestamp 1701862152
transform 1 0 3950 0 -1 8590
box -14 -8 114 272
use OAI21X1  _2382_
timestamp 1702508443
transform -1 0 4730 0 -1 8590
box -12 -8 92 272
use NOR2X1  _2383_
timestamp 1701862152
transform -1 0 5790 0 1 8590
box -12 -8 74 272
use OAI21X1  _2384_
timestamp 1702508443
transform -1 0 6030 0 1 8590
box -12 -8 92 272
use INVX1  _2385_
timestamp 1701862152
transform 1 0 1350 0 -1 10150
box -12 -8 52 272
use NAND2X1  _2386_
timestamp 1702508443
transform 1 0 5610 0 -1 7550
box -12 -8 72 272
use OAI21X1  _2387_
timestamp 1702508443
transform 1 0 5590 0 -1 9110
box -12 -8 92 272
use AOI21X1  _2388_
timestamp 1702508443
transform -1 0 5430 0 -1 9110
box -12 -8 92 272
use OAI21X1  _2389_
timestamp 1702508443
transform -1 0 5230 0 -1 9630
box -12 -8 92 272
use INVX1  _2390_
timestamp 1701862152
transform 1 0 5230 0 1 9630
box -12 -8 52 272
use OAI21X1  _2391_
timestamp 1702508443
transform -1 0 5510 0 1 9630
box -12 -8 92 272
use INVX1  _2392_
timestamp 1701862152
transform 1 0 1550 0 -1 10150
box -12 -8 52 272
use NAND2X1  _2393_
timestamp 1702508443
transform -1 0 5450 0 -1 7550
box -12 -8 72 272
use OAI21X1  _2394_
timestamp 1702508443
transform 1 0 5490 0 1 8590
box -12 -8 92 272
use AOI21X1  _2395_
timestamp 1702508443
transform -1 0 5890 0 -1 9110
box -12 -8 92 272
use OAI21X1  _2396_
timestamp 1702508443
transform 1 0 5770 0 1 9110
box -12 -8 92 272
use INVX1  _2397_
timestamp 1701862152
transform 1 0 6010 0 1 9110
box -12 -8 52 272
use OAI21X1  _2398_
timestamp 1702508443
transform 1 0 5830 0 -1 9630
box -12 -8 92 272
use OAI21X1  _2399_
timestamp 1702508443
transform -1 0 3330 0 -1 5470
box -12 -8 92 272
use NOR2X1  _2400_
timestamp 1701862152
transform -1 0 3490 0 1 5990
box -12 -8 74 272
use INVX2  _2401_
timestamp 1701862152
transform 1 0 3370 0 -1 6510
box -12 -8 52 272
use OAI21X1  _2402_
timestamp 1702508443
transform -1 0 2370 0 -1 4430
box -12 -8 92 272
use AND2X2  _2403_
timestamp 1701862152
transform -1 0 2750 0 1 4430
box -12 -8 94 272
use NAND3X1  _2404_
timestamp 1702508443
transform -1 0 3090 0 -1 5470
box -12 -8 92 272
use AOI21X1  _2405_
timestamp 1702508443
transform 1 0 2410 0 -1 2870
box -12 -8 92 272
use NAND3X1  _2406_
timestamp 1702508443
transform 1 0 3110 0 -1 3390
box -12 -8 92 272
use NOR2X1  _2407_
timestamp 1701862152
transform -1 0 3290 0 1 5470
box -12 -8 74 272
use AOI21X1  _2408_
timestamp 1702508443
transform 1 0 870 0 -1 2870
box -12 -8 92 272
use OAI21X1  _2409_
timestamp 1702508443
transform 1 0 890 0 -1 3910
box -12 -8 92 272
use OAI21X1  _2410_
timestamp 1702508443
transform 1 0 1270 0 1 4430
box -12 -8 92 272
use OAI21X1  _2411_
timestamp 1702508443
transform -1 0 910 0 -1 4950
box -12 -8 92 272
use NOR2X1  _2412_
timestamp 1701862152
transform 1 0 2530 0 -1 5990
box -12 -8 74 272
use OAI21X1  _2413_
timestamp 1702508443
transform 1 0 2990 0 1 5470
box -12 -8 92 272
use OAI21X1  _2414_
timestamp 1702508443
transform 1 0 4150 0 -1 5470
box -12 -8 92 272
use INVX2  _2415_
timestamp 1701862152
transform -1 0 4110 0 1 7030
box -12 -8 52 272
use INVX1  _2416_
timestamp 1701862152
transform 1 0 4050 0 1 4950
box -12 -8 52 272
use OAI21X1  _2417_
timestamp 1702508443
transform 1 0 4370 0 -1 5470
box -12 -8 92 272
use NAND2X1  _2418_
timestamp 1702508443
transform -1 0 1690 0 -1 4950
box -12 -8 72 272
use NAND3X1  _2419_
timestamp 1702508443
transform 1 0 2230 0 1 4430
box -12 -8 92 272
use NOR2X1  _2420_
timestamp 1701862152
transform 1 0 3890 0 1 5990
box -12 -8 74 272
use NAND3X1  _2421_
timestamp 1702508443
transform -1 0 3730 0 1 5990
box -12 -8 92 272
use NOR2X1  _2422_
timestamp 1701862152
transform -1 0 3590 0 -1 5990
box -12 -8 74 272
use NAND2X1  _2423_
timestamp 1702508443
transform -1 0 3810 0 -1 5990
box -12 -8 72 272
use NAND2X1  _2424_
timestamp 1702508443
transform 1 0 3310 0 -1 5990
box -12 -8 72 272
use INVX1  _2425_
timestamp 1701862152
transform 1 0 4430 0 1 5990
box -12 -8 52 272
use NOR2X1  _2426_
timestamp 1701862152
transform 1 0 4050 0 -1 7030
box -12 -8 74 272
use AOI22X1  _2427_
timestamp 1701862152
transform 1 0 4870 0 1 5990
box -14 -8 114 272
use OAI21X1  _2428_
timestamp 1702508443
transform 1 0 4630 0 1 5990
box -12 -8 92 272
use AOI21X1  _2429_
timestamp 1702508443
transform -1 0 4370 0 -1 6510
box -12 -8 92 272
use OAI21X1  _2430_
timestamp 1702508443
transform 1 0 4870 0 1 6510
box -12 -8 92 272
use AOI21X1  _2431_
timestamp 1702508443
transform -1 0 5030 0 -1 7030
box -12 -8 92 272
use INVX1  _2432_
timestamp 1701862152
transform 1 0 5170 0 -1 7030
box -12 -8 52 272
use OR2X2  _2433_
timestamp 1702508443
transform -1 0 4510 0 -1 8070
box -12 -8 92 272
use INVX2  _2434_
timestamp 1701862152
transform 1 0 4930 0 1 7550
box -12 -8 52 272
use OAI21X1  _2435_
timestamp 1702508443
transform 1 0 4270 0 1 7030
box -12 -8 92 272
use OAI21X1  _2436_
timestamp 1702508443
transform -1 0 4770 0 -1 7550
box -12 -8 92 272
use AOI21X1  _2437_
timestamp 1702508443
transform -1 0 4750 0 -1 8070
box -12 -8 92 272
use OAI21X1  _2438_
timestamp 1702508443
transform -1 0 4990 0 -1 8070
box -12 -8 92 272
use AOI21X1  _2439_
timestamp 1702508443
transform -1 0 5210 0 -1 8070
box -12 -8 92 272
use INVX1  _2440_
timestamp 1701862152
transform 1 0 4710 0 1 10150
box -12 -8 52 272
use OAI21X1  _2441_
timestamp 1702508443
transform 1 0 3990 0 -1 7550
box -12 -8 92 272
use OAI21X1  _2442_
timestamp 1702508443
transform -1 0 4270 0 -1 8070
box -12 -8 92 272
use AOI21X1  _2443_
timestamp 1702508443
transform -1 0 4050 0 1 8070
box -12 -8 92 272
use OAI21X1  _2444_
timestamp 1702508443
transform 1 0 3730 0 1 8070
box -12 -8 92 272
use AOI21X1  _2445_
timestamp 1702508443
transform -1 0 4770 0 1 7550
box -12 -8 92 272
use INVX1  _2446_
timestamp 1701862152
transform 1 0 4610 0 1 8070
box -12 -8 52 272
use INVX1  _2447_
timestamp 1701862152
transform 1 0 4370 0 1 9110
box -12 -8 52 272
use OAI22X1  _2448_
timestamp 1701862152
transform 1 0 5030 0 1 9110
box -12 -8 112 272
use AOI21X1  _2449_
timestamp 1702508443
transform 1 0 5290 0 1 9110
box -12 -8 92 272
use OAI21X1  _2450_
timestamp 1702508443
transform 1 0 5530 0 1 9110
box -12 -8 92 272
use AOI21X1  _2451_
timestamp 1702508443
transform -1 0 5470 0 -1 9630
box -12 -8 92 272
use INVX1  _2452_
timestamp 1701862152
transform -1 0 5350 0 -1 10670
box -12 -8 52 272
use INVX1  _2453_
timestamp 1701862152
transform 1 0 3870 0 -1 10150
box -12 -8 52 272
use AOI22X1  _2454_
timestamp 1701862152
transform 1 0 3970 0 1 7550
box -14 -8 114 272
use OAI21X1  _2455_
timestamp 1702508443
transform 1 0 3950 0 -1 8070
box -12 -8 92 272
use AOI21X1  _2456_
timestamp 1702508443
transform -1 0 3790 0 -1 8070
box -12 -8 92 272
use OAI21X1  _2457_
timestamp 1702508443
transform 1 0 3490 0 1 8070
box -12 -8 92 272
use AOI21X1  _2458_
timestamp 1702508443
transform -1 0 4490 0 -1 8590
box -12 -8 92 272
use INVX1  _2459_
timestamp 1701862152
transform -1 0 4610 0 -1 11190
box -12 -8 52 272
use INVX1  _2460_
timestamp 1701862152
transform 1 0 4230 0 -1 10670
box -12 -8 52 272
use OAI22X1  _2461_
timestamp 1701862152
transform 1 0 4390 0 -1 9110
box -12 -8 112 272
use AOI21X1  _2462_
timestamp 1702508443
transform -1 0 4730 0 -1 9110
box -12 -8 92 272
use OAI21X1  _2463_
timestamp 1702508443
transform -1 0 4970 0 -1 9110
box -12 -8 92 272
use AOI21X1  _2464_
timestamp 1702508443
transform -1 0 5210 0 -1 9110
box -12 -8 92 272
use INVX1  _2465_
timestamp 1701862152
transform -1 0 5030 0 -1 11190
box -12 -8 52 272
use INVX1  _2466_
timestamp 1701862152
transform -1 0 4110 0 -1 10150
box -12 -8 52 272
use OAI22X1  _2467_
timestamp 1701862152
transform -1 0 4270 0 -1 9630
box -12 -8 112 272
use AOI21X1  _2468_
timestamp 1702508443
transform -1 0 4490 0 -1 9630
box -12 -8 92 272
use OAI21X1  _2469_
timestamp 1702508443
transform -1 0 4370 0 1 9630
box -12 -8 92 272
use AOI21X1  _2470_
timestamp 1702508443
transform -1 0 4610 0 1 9630
box -12 -8 92 272
use INVX1  _2471_
timestamp 1701862152
transform -1 0 5150 0 -1 10670
box -12 -8 52 272
use INVX1  _2472_
timestamp 1701862152
transform 1 0 4090 0 1 9630
box -12 -8 52 272
use OAI22X1  _2473_
timestamp 1701862152
transform 1 0 4650 0 -1 9630
box -12 -8 112 272
use AOI21X1  _2474_
timestamp 1702508443
transform -1 0 4990 0 -1 9630
box -12 -8 92 272
use OAI21X1  _2475_
timestamp 1702508443
transform 1 0 4750 0 1 9630
box -12 -8 92 272
use AOI21X1  _2476_
timestamp 1702508443
transform -1 0 5070 0 1 9630
box -12 -8 92 272
use INVX1  _2477_
timestamp 1701862152
transform 1 0 4950 0 1 10670
box -12 -8 52 272
use OAI21X1  _2478_
timestamp 1702508443
transform 1 0 3190 0 1 5990
box -12 -8 92 272
use AOI22X1  _2479_
timestamp 1701862152
transform -1 0 2830 0 1 5990
box -14 -8 114 272
use OAI21X1  _2480_
timestamp 1702508443
transform -1 0 2830 0 -1 5990
box -12 -8 92 272
use NOR3X1  _2481_
timestamp 1701862152
transform -1 0 3150 0 -1 5990
box -12 -8 172 272
use OAI21X1  _2482_
timestamp 1702508443
transform 1 0 1590 0 -1 5990
box -12 -8 92 272
use OAI21X1  _2483_
timestamp 1702508443
transform 1 0 2390 0 1 6510
box -12 -8 92 272
use INVX1  _2484_
timestamp 1701862152
transform -1 0 2050 0 1 6510
box -12 -8 52 272
use INVX1  _2485_
timestamp 1701862152
transform -1 0 2250 0 1 6510
box -12 -8 52 272
use AOI22X1  _2486_
timestamp 1701862152
transform 1 0 2430 0 -1 7030
box -14 -8 114 272
use OAI21X1  _2487_
timestamp 1702508443
transform 1 0 2190 0 -1 7030
box -12 -8 92 272
use NOR2X1  _2488_
timestamp 1701862152
transform -1 0 2030 0 -1 7030
box -12 -8 74 272
use OAI21X1  _2489_
timestamp 1702508443
transform 1 0 1490 0 -1 7030
box -12 -8 92 272
use OAI21X1  _2490_
timestamp 1702508443
transform -1 0 1130 0 1 5470
box -12 -8 92 272
use INVX1  _2491_
timestamp 1701862152
transform 1 0 1290 0 1 5470
box -12 -8 52 272
use AOI21X1  _2492_
timestamp 1702508443
transform -1 0 2210 0 -1 6510
box -12 -8 92 272
use OAI21X1  _2493_
timestamp 1702508443
transform 1 0 2030 0 1 5990
box -12 -8 92 272
use NOR2X1  _2494_
timestamp 1701862152
transform -1 0 1630 0 1 5990
box -12 -8 74 272
use OAI21X1  _2495_
timestamp 1702508443
transform 1 0 1330 0 1 5990
box -12 -8 92 272
use OAI21X1  _2496_
timestamp 1702508443
transform 1 0 1730 0 -1 7030
box -12 -8 92 272
use INVX1  _2497_
timestamp 1701862152
transform -1 0 1930 0 -1 7550
box -12 -8 52 272
use INVX1  _2498_
timestamp 1701862152
transform 1 0 870 0 1 8070
box -12 -8 52 272
use AOI22X1  _2499_
timestamp 1701862152
transform 1 0 2550 0 1 7550
box -14 -8 114 272
use OAI21X1  _2500_
timestamp 1702508443
transform 1 0 1970 0 1 7550
box -12 -8 92 272
use NOR2X1  _2501_
timestamp 1701862152
transform 1 0 1750 0 1 7550
box -12 -8 74 272
use OAI21X1  _2502_
timestamp 1702508443
transform -1 0 1350 0 1 7550
box -12 -8 92 272
use INVX1  _2503_
timestamp 1701862152
transform -1 0 1550 0 1 8070
box -12 -8 52 272
use NAND2X1  _2504_
timestamp 1702508443
transform -1 0 1990 0 1 8070
box -12 -8 72 272
use OAI21X1  _2505_
timestamp 1702508443
transform 1 0 1270 0 1 8070
box -12 -8 92 272
use OAI21X1  _2506_
timestamp 1702508443
transform -1 0 1870 0 -1 8070
box -12 -8 92 272
use OAI21X1  _2507_
timestamp 1702508443
transform 1 0 1550 0 -1 8070
box -12 -8 92 272
use NOR2X1  _2508_
timestamp 1701862152
transform 1 0 1070 0 1 8070
box -12 -8 74 272
use OAI21X1  _2509_
timestamp 1702508443
transform 1 0 630 0 -1 8590
box -12 -8 92 272
use INVX1  _2510_
timestamp 1701862152
transform -1 0 1590 0 1 9110
box -12 -8 52 272
use OAI21X1  _2511_
timestamp 1702508443
transform -1 0 1570 0 -1 9630
box -12 -8 92 272
use INVX1  _2512_
timestamp 1701862152
transform 1 0 1050 0 -1 9630
box -12 -8 52 272
use INVX1  _2513_
timestamp 1701862152
transform -1 0 1090 0 1 8590
box -12 -8 52 272
use AOI22X1  _2514_
timestamp 1701862152
transform 1 0 2150 0 -1 8590
box -14 -8 114 272
use OAI21X1  _2515_
timestamp 1702508443
transform 1 0 1270 0 -1 9110
box -12 -8 92 272
use NOR2X1  _2516_
timestamp 1701862152
transform -1 0 1150 0 1 9110
box -12 -8 74 272
use OAI21X1  _2517_
timestamp 1702508443
transform -1 0 930 0 1 9110
box -12 -8 92 272
use OAI21X1  _2518_
timestamp 1702508443
transform 1 0 1730 0 -1 9630
box -12 -8 92 272
use INVX1  _2519_
timestamp 1701862152
transform 1 0 1810 0 1 9630
box -12 -8 52 272
use AOI21X1  _2520_
timestamp 1702508443
transform -1 0 2730 0 -1 9110
box -12 -8 92 272
use OAI21X1  _2521_
timestamp 1702508443
transform 1 0 2410 0 -1 9110
box -12 -8 92 272
use NOR2X1  _2522_
timestamp 1701862152
transform -1 0 2070 0 1 9630
box -12 -8 74 272
use OAI21X1  _2523_
timestamp 1702508443
transform -1 0 2310 0 1 9630
box -12 -8 92 272
use OAI21X1  _2524_
timestamp 1702508443
transform -1 0 2050 0 -1 9110
box -12 -8 92 272
use INVX1  _2525_
timestamp 1701862152
transform 1 0 870 0 -1 8590
box -12 -8 52 272
use AOI21X1  _2526_
timestamp 1702508443
transform -1 0 1810 0 -1 8590
box -12 -8 92 272
use OAI21X1  _2527_
timestamp 1702508443
transform -1 0 1370 0 -1 8590
box -12 -8 92 272
use NOR2X1  _2528_
timestamp 1701862152
transform -1 0 1130 0 -1 8590
box -12 -8 74 272
use OAI21X1  _2529_
timestamp 1702508443
transform -1 0 1390 0 1 9110
box -12 -8 92 272
use AND2X2  _2530_
timestamp 1701862152
transform -1 0 7650 0 -1 6510
box -12 -8 94 272
use AND2X2  _2531_
timestamp 1701862152
transform 1 0 8010 0 1 7550
box -12 -8 94 272
use INVX1  _2532_
timestamp 1701862152
transform -1 0 9930 0 1 2870
box -12 -8 52 272
use NOR2X1  _2533_
timestamp 1701862152
transform -1 0 9030 0 1 4430
box -12 -8 74 272
use INVX8  _2534_
timestamp 1701862152
transform -1 0 9450 0 -1 5470
box -12 -8 114 272
use OAI21X1  _2535_
timestamp 1702508443
transform 1 0 170 0 -1 4950
box -12 -8 92 272
use NOR2X1  _2536_
timestamp 1701862152
transform 1 0 730 0 1 4950
box -12 -8 74 272
use NAND2X1  _2537_
timestamp 1702508443
transform 1 0 870 0 1 3390
box -12 -8 72 272
use OAI21X1  _2538_
timestamp 1702508443
transform -1 0 490 0 -1 3910
box -12 -8 92 272
use NOR3X1  _2539_
timestamp 1701862152
transform -1 0 330 0 1 4950
box -12 -8 172 272
use NAND3X1  _2540_
timestamp 1702508443
transform 1 0 3130 0 1 2350
box -12 -8 92 272
use NOR2X1  _2541_
timestamp 1701862152
transform -1 0 3410 0 1 2870
box -12 -8 74 272
use NAND2X1  _2542_
timestamp 1702508443
transform -1 0 2430 0 -1 6510
box -12 -8 72 272
use NAND2X1  _2543_
timestamp 1702508443
transform 1 0 950 0 1 4950
box -12 -8 72 272
use OAI22X1  _2544_
timestamp 1701862152
transform 1 0 1510 0 1 4430
box -12 -8 112 272
use NAND3X1  _2545_
timestamp 1702508443
transform 1 0 1370 0 -1 5470
box -12 -8 92 272
use NAND3X1  _2546_
timestamp 1702508443
transform -1 0 2170 0 -1 5470
box -12 -8 92 272
use NAND3X1  _2547_
timestamp 1702508443
transform 1 0 2050 0 -1 4430
box -12 -8 92 272
use OAI21X1  _2548_
timestamp 1702508443
transform 1 0 1150 0 1 4950
box -12 -8 92 272
use INVX1  _2549_
timestamp 1701862152
transform 1 0 1390 0 1 4950
box -12 -8 52 272
use OAI21X1  _2550_
timestamp 1702508443
transform -1 0 1930 0 -1 5470
box -12 -8 92 272
use INVX2  _2551_
timestamp 1701862152
transform 1 0 2650 0 -1 9630
box -12 -8 52 272
use NOR2X1  _2552_
timestamp 1701862152
transform 1 0 3490 0 -1 5470
box -12 -8 74 272
use AOI22X1  _2553_
timestamp 1701862152
transform -1 0 2950 0 -1 6510
box -14 -8 114 272
use OAI21X1  _2554_
timestamp 1702508443
transform -1 0 3390 0 1 6510
box -12 -8 92 272
use NOR2X1  _2555_
timestamp 1701862152
transform -1 0 3590 0 1 6510
box -12 -8 74 272
use NAND2X1  _2556_
timestamp 1702508443
transform -1 0 2930 0 1 6510
box -12 -8 72 272
use AOI22X1  _2557_
timestamp 1701862152
transform 1 0 2590 0 -1 6510
box -14 -8 114 272
use INVX1  _2558_
timestamp 1701862152
transform 1 0 3330 0 -1 7550
box -12 -8 52 272
use NAND2X1  _2559_
timestamp 1702508443
transform 1 0 3530 0 -1 7550
box -12 -8 72 272
use OAI22X1  _2560_
timestamp 1701862152
transform -1 0 3670 0 1 7030
box -12 -8 112 272
use OAI21X1  _2561_
timestamp 1702508443
transform -1 0 1670 0 1 4950
box -12 -8 92 272
use OAI21X1  _2562_
timestamp 1702508443
transform 1 0 3330 0 1 7030
box -12 -8 92 272
use INVX1  _2563_
timestamp 1701862152
transform 1 0 3870 0 1 5470
box -12 -8 52 272
use AOI22X1  _2564_
timestamp 1701862152
transform -1 0 3850 0 1 6510
box -14 -8 114 272
use AND2X2  _2565_
timestamp 1701862152
transform 1 0 3830 0 1 7030
box -12 -8 94 272
use OAI21X1  _2566_
timestamp 1702508443
transform 1 0 3290 0 1 7550
box -12 -8 92 272
use NOR2X1  _2567_
timestamp 1701862152
transform 1 0 3250 0 -1 8070
box -12 -8 74 272
use NAND2X1  _2568_
timestamp 1702508443
transform -1 0 3110 0 -1 8590
box -12 -8 72 272
use NAND2X1  _2569_
timestamp 1702508443
transform 1 0 2830 0 -1 8590
box -12 -8 72 272
use OAI22X1  _2570_
timestamp 1701862152
transform 1 0 2990 0 -1 8070
box -12 -8 112 272
use NAND2X1  _2571_
timestamp 1702508443
transform -1 0 4010 0 -1 9630
box -12 -8 72 272
use NOR2X1  _2572_
timestamp 1701862152
transform -1 0 4030 0 -1 5990
box -12 -8 74 272
use NAND2X1  _2573_
timestamp 1702508443
transform -1 0 3890 0 -1 7030
box -12 -8 72 272
use OAI21X1  _2574_
timestamp 1702508443
transform 1 0 3570 0 -1 6510
box -12 -8 92 272
use AOI21X1  _2575_
timestamp 1702508443
transform 1 0 3470 0 -1 8070
box -12 -8 92 272
use OAI21X1  _2576_
timestamp 1702508443
transform -1 0 3570 0 -1 8590
box -12 -8 92 272
use XOR2X1  _2577_
timestamp 1702508443
transform 1 0 3370 0 1 9110
box -12 -8 132 272
use OAI21X1  _2578_
timestamp 1702508443
transform 1 0 3890 0 1 9110
box -12 -8 92 272
use INVX1  _2579_
timestamp 1701862152
transform -1 0 2890 0 -1 9630
box -12 -8 52 272
use INVX2  _2580_
timestamp 1701862152
transform -1 0 4250 0 -1 9110
box -12 -8 52 272
use OAI21X1  _2581_
timestamp 1702508443
transform -1 0 4210 0 1 9110
box -12 -8 92 272
use AOI21X1  _2582_
timestamp 1702508443
transform 1 0 3650 0 1 9110
box -12 -8 92 272
use OAI21X1  _2583_
timestamp 1702508443
transform 1 0 3150 0 1 9110
box -12 -8 92 272
use AOI21X1  _2584_
timestamp 1702508443
transform 1 0 2910 0 1 9110
box -12 -8 92 272
use NAND2X1  _2585_
timestamp 1702508443
transform 1 0 3990 0 -1 9110
box -12 -8 72 272
use NAND2X1  _2586_
timestamp 1702508443
transform 1 0 3170 0 1 9630
box -12 -8 72 272
use AOI22X1  _2587_
timestamp 1701862152
transform 1 0 3750 0 -1 9110
box -14 -8 114 272
use NAND3X1  _2588_
timestamp 1702508443
transform 1 0 3350 0 1 8590
box -12 -8 92 272
use NAND2X1  _2589_
timestamp 1702508443
transform 1 0 3190 0 -1 10150
box -12 -8 72 272
use OAI22X1  _2590_
timestamp 1701862152
transform 1 0 2930 0 -1 10150
box -12 -8 112 272
use NAND2X1  _2591_
timestamp 1702508443
transform -1 0 3730 0 -1 11190
box -12 -8 72 272
use OAI21X1  _2592_
timestamp 1702508443
transform -1 0 3790 0 -1 9630
box -12 -8 92 272
use AOI21X1  _2593_
timestamp 1702508443
transform -1 0 3330 0 -1 9630
box -12 -8 92 272
use OAI21X1  _2594_
timestamp 1702508443
transform -1 0 3490 0 -1 10150
box -12 -8 92 272
use XOR2X1  _2595_
timestamp 1702508443
transform 1 0 3150 0 -1 11190
box -12 -8 132 272
use OAI21X1  _2596_
timestamp 1702508443
transform 1 0 3430 0 -1 11190
box -12 -8 92 272
use INVX1  _2597_
timestamp 1701862152
transform 1 0 2890 0 -1 10670
box -12 -8 52 272
use OAI21X1  _2598_
timestamp 1702508443
transform -1 0 3690 0 1 9630
box -12 -8 92 272
use AOI21X1  _2599_
timestamp 1702508443
transform -1 0 3450 0 1 9630
box -12 -8 92 272
use OAI21X1  _2600_
timestamp 1702508443
transform -1 0 3190 0 1 10150
box -12 -8 92 272
use AOI21X1  _2601_
timestamp 1702508443
transform 1 0 3090 0 -1 10670
box -12 -8 92 272
use NAND2X1  _2602_
timestamp 1702508443
transform -1 0 3390 0 -1 10670
box -12 -8 72 272
use NAND2X1  _2603_
timestamp 1702508443
transform 1 0 3550 0 -1 10670
box -12 -8 72 272
use AOI22X1  _2604_
timestamp 1701862152
transform 1 0 3350 0 1 10150
box -14 -8 114 272
use INVX1  _2605_
timestamp 1701862152
transform 1 0 2470 0 1 10670
box -12 -8 52 272
use OAI21X1  _2606_
timestamp 1702508443
transform 1 0 2650 0 1 10670
box -12 -8 92 272
use OAI22X1  _2607_
timestamp 1701862152
transform -1 0 2990 0 1 10670
box -12 -8 112 272
use OAI21X1  _2608_
timestamp 1702508443
transform -1 0 3930 0 1 9630
box -12 -8 92 272
use AOI21X1  _2609_
timestamp 1702508443
transform -1 0 2550 0 1 9630
box -12 -8 92 272
use OAI21X1  _2610_
timestamp 1702508443
transform -1 0 2770 0 -1 10150
box -12 -8 92 272
use AOI21X1  _2611_
timestamp 1702508443
transform -1 0 2490 0 -1 10670
box -12 -8 92 272
use NAND3X1  _2612_
timestamp 1702508443
transform 1 0 2650 0 -1 10670
box -12 -8 92 272
use NAND2X1  _2613_
timestamp 1702508443
transform 1 0 1970 0 1 10670
box -12 -8 72 272
use OAI22X1  _2614_
timestamp 1701862152
transform 1 0 1950 0 -1 10670
box -12 -8 112 272
use NAND2X1  _2615_
timestamp 1702508443
transform -1 0 2530 0 -1 11190
box -12 -8 72 272
use OAI21X1  _2616_
timestamp 1702508443
transform -1 0 3570 0 -1 9630
box -12 -8 92 272
use AOI21X1  _2617_
timestamp 1702508443
transform 1 0 2410 0 -1 9630
box -12 -8 92 272
use OAI21X1  _2618_
timestamp 1702508443
transform -1 0 2750 0 1 10150
box -12 -8 92 272
use XOR2X1  _2619_
timestamp 1702508443
transform 1 0 2190 0 1 10670
box -12 -8 132 272
use OAI21X1  _2620_
timestamp 1702508443
transform 1 0 2230 0 -1 11190
box -12 -8 92 272
use AOI21X1  _2621_
timestamp 1702508443
transform -1 0 1550 0 1 5470
box -12 -8 92 272
use OAI22X1  _2622_
timestamp 1701862152
transform -1 0 1430 0 -1 5990
box -12 -8 112 272
use NAND3X1  _2623_
timestamp 1702508443
transform 1 0 2570 0 -1 5470
box -12 -8 92 272
use NAND3X1  _2624_
timestamp 1702508443
transform -1 0 2590 0 1 5470
box -12 -8 92 272
use NAND3X1  _2625_
timestamp 1702508443
transform 1 0 2330 0 -1 5470
box -12 -8 92 272
use NOR3X1  _2626_
timestamp 1701862152
transform -1 0 1210 0 -1 5470
box -12 -8 172 272
use AOI22X1  _2627_
timestamp 1701862152
transform -1 0 1670 0 1 3910
box -14 -8 114 272
use NOR3X1  _2628_
timestamp 1701862152
transform 1 0 1250 0 1 3910
box -12 -8 172 272
use INVX1  _2629_
timestamp 1701862152
transform -1 0 890 0 -1 5470
box -12 -8 52 272
use NAND3X1  _2630_
timestamp 1702508443
transform 1 0 850 0 -1 5990
box -12 -8 92 272
use AND2X2  _2631_
timestamp 1701862152
transform -1 0 910 0 1 5990
box -12 -8 94 272
use NAND2X1  _2632_
timestamp 1702508443
transform 1 0 2230 0 1 10150
box -12 -8 72 272
use NAND2X1  _2633_
timestamp 1702508443
transform -1 0 2510 0 1 10150
box -12 -8 72 272
use AOI22X1  _2634_
timestamp 1701862152
transform 1 0 2430 0 -1 10150
box -14 -8 114 272
use NAND2X1  _2635_
timestamp 1702508443
transform 1 0 2210 0 -1 10150
box -12 -8 72 272
use NOR2X1  _2636_
timestamp 1701862152
transform -1 0 870 0 -1 10150
box -12 -8 74 272
use AND2X2  _2637_
timestamp 1701862152
transform -1 0 710 0 1 6510
box -12 -8 94 272
use NOR2X1  _2638_
timestamp 1701862152
transform -1 0 470 0 1 6510
box -12 -8 74 272
use OAI21X1  _2639_
timestamp 1702508443
transform -1 0 470 0 -1 6510
box -12 -8 92 272
use OAI21X1  _2640_
timestamp 1702508443
transform -1 0 470 0 1 5990
box -12 -8 92 272
use INVX1  _2641_
timestamp 1701862152
transform 1 0 170 0 -1 7550
box -12 -8 52 272
use AOI21X1  _2642_
timestamp 1702508443
transform -1 0 570 0 1 4950
box -12 -8 92 272
use AOI22X1  _2643_
timestamp 1701862152
transform -1 0 2710 0 1 6510
box -14 -8 114 272
use NAND3X1  _2644_
timestamp 1702508443
transform 1 0 2690 0 -1 7030
box -12 -8 92 272
use AOI21X1  _2645_
timestamp 1702508443
transform 1 0 2870 0 1 7030
box -12 -8 92 272
use OAI21X1  _2646_
timestamp 1702508443
transform 1 0 2170 0 1 7030
box -12 -8 92 272
use INVX1  _2647_
timestamp 1701862152
transform 1 0 850 0 1 7550
box -12 -8 52 272
use AOI21X1  _2648_
timestamp 1702508443
transform 1 0 390 0 1 7550
box -12 -8 92 272
use NAND2X1  _2649_
timestamp 1702508443
transform 1 0 370 0 -1 7550
box -12 -8 72 272
use NOR2X1  _2650_
timestamp 1701862152
transform -1 0 870 0 -1 7550
box -12 -8 74 272
use OAI21X1  _2651_
timestamp 1702508443
transform 1 0 590 0 -1 7550
box -12 -8 92 272
use OAI21X1  _2652_
timestamp 1702508443
transform 1 0 590 0 1 7030
box -12 -8 92 272
use NOR2X1  _2653_
timestamp 1701862152
transform 1 0 170 0 1 7550
box -12 -8 74 272
use NAND2X1  _2654_
timestamp 1702508443
transform -1 0 690 0 1 7550
box -12 -8 72 272
use INVX1  _2655_
timestamp 1701862152
transform 1 0 1970 0 1 7030
box -12 -8 52 272
use AOI21X1  _2656_
timestamp 1702508443
transform 1 0 1610 0 -1 5470
box -12 -8 92 272
use OAI22X1  _2657_
timestamp 1701862152
transform -1 0 1870 0 1 5990
box -12 -8 112 272
use NAND3X1  _2658_
timestamp 1702508443
transform -1 0 2350 0 1 5470
box -12 -8 92 272
use NAND3X1  _2659_
timestamp 1702508443
transform 1 0 2050 0 -1 5990
box -12 -8 92 272
use NAND3X1  _2660_
timestamp 1702508443
transform -1 0 2110 0 1 5470
box -12 -8 92 272
use NOR3X1  _2661_
timestamp 1701862152
transform -1 0 1870 0 1 5470
box -12 -8 172 272
use NAND3X1  _2662_
timestamp 1702508443
transform 1 0 830 0 1 5470
box -12 -8 92 272
use AND2X2  _2663_
timestamp 1701862152
transform -1 0 1170 0 -1 5990
box -12 -8 94 272
use INVX1  _2664_
timestamp 1701862152
transform 1 0 830 0 -1 7030
box -12 -8 52 272
use NOR2X1  _2665_
timestamp 1701862152
transform 1 0 1270 0 -1 7030
box -12 -8 74 272
use OAI21X1  _2666_
timestamp 1702508443
transform 1 0 1490 0 1 7030
box -12 -8 92 272
use OAI22X1  _2667_
timestamp 1701862152
transform 1 0 1030 0 -1 7030
box -12 -8 112 272
use AOI22X1  _2668_
timestamp 1701862152
transform -1 0 2910 0 1 7550
box -14 -8 114 272
use NAND3X1  _2669_
timestamp 1702508443
transform 1 0 2770 0 -1 8070
box -12 -8 92 272
use AOI21X1  _2670_
timestamp 1702508443
transform 1 0 2030 0 -1 8070
box -12 -8 92 272
use OAI21X1  _2671_
timestamp 1702508443
transform -1 0 1590 0 1 7550
box -12 -8 92 272
use INVX1  _2672_
timestamp 1701862152
transform 1 0 1230 0 -1 7550
box -12 -8 52 272
use OAI21X1  _2673_
timestamp 1702508443
transform -1 0 1510 0 -1 7550
box -12 -8 92 272
use NAND3X1  _2674_
timestamp 1702508443
transform 1 0 1730 0 1 7030
box -12 -8 92 272
use NAND3X1  _2675_
timestamp 1702508443
transform 1 0 1670 0 -1 7550
box -12 -8 92 272
use OAI21X1  _2676_
timestamp 1702508443
transform -1 0 2170 0 -1 7550
box -12 -8 92 272
use AOI22X1  _2677_
timestamp 1701862152
transform 1 0 2510 0 -1 8070
box -14 -8 114 272
use NAND3X1  _2678_
timestamp 1702508443
transform -1 0 2350 0 -1 8070
box -12 -8 92 272
use AOI21X1  _2679_
timestamp 1702508443
transform -1 0 1770 0 1 8070
box -12 -8 92 272
use OAI21X1  _2680_
timestamp 1702508443
transform -1 0 470 0 -1 8590
box -12 -8 92 272
use NOR2X1  _2681_
timestamp 1701862152
transform 1 0 1030 0 -1 7550
box -12 -8 74 272
use NAND3X1  _2682_
timestamp 1702508443
transform -1 0 470 0 -1 8070
box -12 -8 92 272
use NOR2X1  _2683_
timestamp 1701862152
transform -1 0 230 0 -1 9630
box -12 -8 74 272
use INVX1  _2684_
timestamp 1701862152
transform -1 0 210 0 1 10150
box -12 -8 52 272
use AOI22X1  _2685_
timestamp 1701862152
transform 1 0 1070 0 1 5990
box -14 -8 114 272
use NAND3X1  _2686_
timestamp 1702508443
transform 1 0 1030 0 1 7550
box -12 -8 92 272
use NOR3X1  _2687_
timestamp 1701862152
transform -1 0 1190 0 -1 10150
box -12 -8 172 272
use NOR2X1  _2688_
timestamp 1701862152
transform 1 0 170 0 -1 10150
box -12 -8 74 272
use OAI21X1  _2689_
timestamp 1702508443
transform 1 0 390 0 -1 9630
box -12 -8 92 272
use OAI21X1  _2690_
timestamp 1702508443
transform 1 0 390 0 1 9110
box -12 -8 92 272
use AOI22X1  _2691_
timestamp 1701862152
transform 1 0 2850 0 1 8590
box -14 -8 114 272
use NAND3X1  _2692_
timestamp 1702508443
transform 1 0 2610 0 1 8590
box -12 -8 92 272
use AOI21X1  _2693_
timestamp 1702508443
transform -1 0 1330 0 -1 9630
box -12 -8 92 272
use OAI21X1  _2694_
timestamp 1702508443
transform 1 0 830 0 -1 9630
box -12 -8 92 272
use OAI21X1  _2695_
timestamp 1702508443
transform 1 0 170 0 1 9630
box -12 -8 92 272
use INVX1  _2696_
timestamp 1701862152
transform -1 0 670 0 -1 10150
box -12 -8 52 272
use NAND3X1  _2697_
timestamp 1702508443
transform 1 0 390 0 -1 10150
box -12 -8 92 272
use NAND3X1  _2698_
timestamp 1702508443
transform 1 0 410 0 1 9630
box -12 -8 92 272
use NAND2X1  _2699_
timestamp 1702508443
transform 1 0 630 0 -1 9630
box -12 -8 72 272
use AND2X2  _2700_
timestamp 1701862152
transform 1 0 650 0 1 9630
box -12 -8 94 272
use NAND2X1  _2701_
timestamp 1702508443
transform -1 0 890 0 -1 10670
box -12 -8 72 272
use AOI22X1  _2702_
timestamp 1701862152
transform 1 0 3590 0 1 8590
box -14 -8 114 272
use NAND3X1  _2703_
timestamp 1702508443
transform -1 0 3190 0 1 8590
box -12 -8 92 272
use AOI21X1  _2704_
timestamp 1702508443
transform -1 0 1670 0 1 9630
box -12 -8 92 272
use OAI21X1  _2705_
timestamp 1702508443
transform 1 0 1350 0 1 9630
box -12 -8 92 272
use NOR2X1  _2706_
timestamp 1701862152
transform 1 0 370 0 1 10150
box -12 -8 74 272
use NAND2X1  _2707_
timestamp 1702508443
transform -1 0 650 0 1 10150
box -12 -8 72 272
use XOR2X1  _2708_
timestamp 1702508443
transform 1 0 790 0 1 10150
box -12 -8 132 272
use OAI21X1  _2709_
timestamp 1702508443
transform -1 0 690 0 -1 10670
box -12 -8 92 272
use NAND2X1  _2710_
timestamp 1702508443
transform 1 0 1810 0 1 10150
box -12 -8 72 272
use AOI22X1  _2711_
timestamp 1701862152
transform 1 0 2350 0 1 8590
box -14 -8 114 272
use NAND3X1  _2712_
timestamp 1702508443
transform -1 0 2190 0 1 8590
box -12 -8 92 272
use AOI21X1  _2713_
timestamp 1702508443
transform -1 0 2050 0 -1 9630
box -12 -8 92 272
use OAI21X1  _2714_
timestamp 1702508443
transform 1 0 1750 0 -1 10150
box -12 -8 92 272
use NAND3X1  _2715_
timestamp 1702508443
transform 1 0 1070 0 1 10150
box -12 -8 92 272
use XOR2X1  _2716_
timestamp 1702508443
transform 1 0 1290 0 1 10150
box -12 -8 132 272
use OAI21X1  _2717_
timestamp 1702508443
transform 1 0 1570 0 1 10150
box -12 -8 92 272
use INVX1  _2718_
timestamp 1701862152
transform -1 0 10170 0 1 4950
box -12 -8 52 272
use NAND3X1  _2719_
timestamp 1702508443
transform -1 0 9970 0 1 4950
box -12 -8 92 272
use OAI21X1  _2720_
timestamp 1702508443
transform -1 0 4750 0 1 4950
box -12 -8 92 272
use INVX1  _2721_
timestamp 1701862152
transform -1 0 7470 0 -1 2350
box -12 -8 52 272
use INVX2  _2722_
timestamp 1701862152
transform 1 0 10090 0 -1 790
box -12 -8 52 272
use NAND2X1  _2723_
timestamp 1702508443
transform -1 0 7230 0 1 1830
box -12 -8 72 272
use OAI21X1  _2724_
timestamp 1702508443
transform -1 0 7270 0 -1 2350
box -12 -8 92 272
use NAND2X1  _2725_
timestamp 1702508443
transform 1 0 7070 0 1 3390
box -12 -8 72 272
use OAI21X1  _2726_
timestamp 1702508443
transform -1 0 7370 0 1 3390
box -12 -8 92 272
use NAND2X1  _2727_
timestamp 1702508443
transform -1 0 5570 0 1 3390
box -12 -8 72 272
use OAI21X1  _2728_
timestamp 1702508443
transform -1 0 5810 0 1 3390
box -12 -8 92 272
use INVX2  _2729_
timestamp 1701862152
transform -1 0 6870 0 -1 3910
box -12 -8 52 272
use OAI22X1  _2730_
timestamp 1701862152
transform 1 0 8330 0 -1 3910
box -12 -8 112 272
use INVX1  _2731_
timestamp 1701862152
transform 1 0 9370 0 1 1830
box -12 -8 52 272
use NOR2X1  _2732_
timestamp 1701862152
transform 1 0 7810 0 1 1830
box -12 -8 74 272
use NAND2X1  _2733_
timestamp 1702508443
transform 1 0 8690 0 1 2350
box -12 -8 72 272
use OAI21X1  _2734_
timestamp 1702508443
transform 1 0 7270 0 -1 5470
box -12 -8 92 272
use OAI21X1  _2735_
timestamp 1702508443
transform 1 0 7350 0 -1 2870
box -12 -8 92 272
use NAND2X1  _2736_
timestamp 1702508443
transform -1 0 7670 0 1 1310
box -12 -8 72 272
use OR2X2  _2737_
timestamp 1702508443
transform 1 0 8670 0 1 1830
box -12 -8 92 272
use OAI21X1  _2738_
timestamp 1702508443
transform -1 0 8130 0 -1 2870
box -12 -8 92 272
use INVX1  _2739_
timestamp 1701862152
transform -1 0 7910 0 1 2870
box -12 -8 52 272
use NOR2X1  _2740_
timestamp 1701862152
transform -1 0 6710 0 -1 1830
box -12 -8 74 272
use NAND2X1  _2741_
timestamp 1702508443
transform 1 0 6870 0 -1 1830
box -12 -8 72 272
use OAI22X1  _2742_
timestamp 1701862152
transform -1 0 8390 0 -1 2870
box -12 -8 112 272
use OAI21X1  _2743_
timestamp 1702508443
transform -1 0 8390 0 1 2870
box -12 -8 92 272
use NOR2X1  _2744_
timestamp 1701862152
transform -1 0 7490 0 -1 270
box -12 -8 74 272
use NAND2X1  _2745_
timestamp 1702508443
transform -1 0 7430 0 1 1830
box -12 -8 72 272
use OAI21X1  _2746_
timestamp 1702508443
transform 1 0 8070 0 1 2870
box -12 -8 92 272
use INVX1  _2747_
timestamp 1701862152
transform -1 0 7890 0 -1 2350
box -12 -8 52 272
use OAI22X1  _2748_
timestamp 1701862152
transform 1 0 8050 0 -1 2350
box -12 -8 112 272
use OAI21X1  _2749_
timestamp 1702508443
transform 1 0 6010 0 1 1830
box -12 -8 92 272
use NAND2X1  _2750_
timestamp 1702508443
transform -1 0 6810 0 -1 1310
box -12 -8 72 272
use OAI21X1  _2751_
timestamp 1702508443
transform -1 0 6550 0 1 1830
box -12 -8 92 272
use INVX1  _2752_
timestamp 1701862152
transform -1 0 7850 0 1 2350
box -12 -8 52 272
use OAI22X1  _2753_
timestamp 1701862152
transform -1 0 7670 0 1 2350
box -12 -8 112 272
use INVX1  _2754_
timestamp 1701862152
transform 1 0 8930 0 -1 4950
box -12 -8 52 272
use NOR2X1  _2755_
timestamp 1701862152
transform 1 0 9830 0 1 790
box -12 -8 74 272
use NAND2X1  _2756_
timestamp 1702508443
transform -1 0 10110 0 1 790
box -12 -8 72 272
use NOR2X1  _2757_
timestamp 1701862152
transform 1 0 10770 0 -1 2870
box -12 -8 74 272
use NAND2X1  _2758_
timestamp 1702508443
transform -1 0 9310 0 -1 2870
box -12 -8 72 272
use OAI21X1  _2759_
timestamp 1702508443
transform 1 0 9170 0 1 4430
box -12 -8 92 272
use NOR2X1  _2760_
timestamp 1701862152
transform 1 0 10530 0 -1 790
box -12 -8 74 272
use NAND3X1  _2761_
timestamp 1702508443
transform 1 0 10290 0 -1 790
box -12 -8 92 272
use OR2X2  _2762_
timestamp 1702508443
transform -1 0 11030 0 -1 1830
box -12 -8 92 272
use OAI21X1  _2763_
timestamp 1702508443
transform 1 0 6710 0 1 1830
box -12 -8 92 272
use OAI21X1  _2764_
timestamp 1702508443
transform -1 0 7030 0 1 1830
box -12 -8 92 272
use NOR2X1  _2765_
timestamp 1701862152
transform -1 0 10310 0 1 1830
box -12 -8 74 272
use NOR2X1  _2766_
timestamp 1701862152
transform -1 0 10130 0 -1 1830
box -12 -8 74 272
use OAI21X1  _2767_
timestamp 1702508443
transform -1 0 10550 0 -1 1830
box -12 -8 92 272
use OAI21X1  _2768_
timestamp 1702508443
transform -1 0 10550 0 1 1830
box -12 -8 92 272
use NOR2X1  _2769_
timestamp 1701862152
transform -1 0 10990 0 1 2350
box -12 -8 74 272
use OAI21X1  _2770_
timestamp 1702508443
transform -1 0 10790 0 -1 1830
box -12 -8 92 272
use OAI21X1  _2771_
timestamp 1702508443
transform 1 0 11150 0 1 2350
box -12 -8 92 272
use INVX1  _2772_
timestamp 1701862152
transform -1 0 10830 0 1 4950
box -12 -8 52 272
use AOI22X1  _2773_
timestamp 1701862152
transform 1 0 10550 0 -1 3910
box -14 -8 114 272
use NOR2X1  _2774_
timestamp 1701862152
transform -1 0 10870 0 -1 2350
box -12 -8 74 272
use INVX1  _2775_
timestamp 1701862152
transform -1 0 9230 0 -1 1310
box -12 -8 52 272
use INVX1  _2776_
timestamp 1701862152
transform 1 0 10750 0 -1 790
box -12 -8 52 272
use NAND2X1  _2777_
timestamp 1702508443
transform -1 0 8550 0 -1 270
box -12 -8 72 272
use OR2X2  _2778_
timestamp 1702508443
transform 1 0 11050 0 1 270
box -12 -8 92 272
use NOR2X1  _2779_
timestamp 1701862152
transform 1 0 9130 0 -1 1830
box -12 -8 74 272
use AOI21X1  _2780_
timestamp 1702508443
transform -1 0 10210 0 1 1310
box -12 -8 92 272
use OAI21X1  _2781_
timestamp 1702508443
transform 1 0 10270 0 -1 1310
box -12 -8 92 272
use NAND2X1  _2782_
timestamp 1702508443
transform 1 0 8910 0 1 1830
box -12 -8 72 272
use NAND3X1  _2783_
timestamp 1702508443
transform 1 0 8470 0 -1 1310
box -12 -8 92 272
use OAI22X1  _2784_
timestamp 1701862152
transform 1 0 8710 0 -1 1310
box -12 -8 112 272
use INVX1  _2785_
timestamp 1701862152
transform 1 0 8930 0 -1 1830
box -12 -8 52 272
use NAND2X1  _2786_
timestamp 1702508443
transform -1 0 9450 0 -1 1310
box -12 -8 72 272
use OAI21X1  _2787_
timestamp 1702508443
transform -1 0 9670 0 -1 1830
box -12 -8 92 272
use NOR2X1  _2788_
timestamp 1701862152
transform 1 0 10270 0 -1 1830
box -12 -8 74 272
use INVX1  _2789_
timestamp 1701862152
transform 1 0 10370 0 1 1310
box -12 -8 52 272
use NAND2X1  _2790_
timestamp 1702508443
transform -1 0 10210 0 -1 2350
box -12 -8 72 272
use NOR2X1  _2791_
timestamp 1701862152
transform 1 0 9930 0 -1 2350
box -12 -8 74 272
use OAI21X1  _2792_
timestamp 1702508443
transform -1 0 10450 0 -1 2350
box -12 -8 92 272
use NAND2X1  _2793_
timestamp 1702508443
transform -1 0 10670 0 -1 2350
box -12 -8 72 272
use OAI21X1  _2794_
timestamp 1702508443
transform -1 0 11110 0 -1 2350
box -12 -8 92 272
use OAI21X1  _2795_
timestamp 1702508443
transform -1 0 11070 0 -1 2870
box -12 -8 92 272
use INVX1  _2796_
timestamp 1701862152
transform -1 0 10350 0 -1 2870
box -12 -8 52 272
use OAI21X1  _2797_
timestamp 1702508443
transform -1 0 9910 0 -1 1830
box -12 -8 92 272
use NOR2X1  _2798_
timestamp 1701862152
transform -1 0 10770 0 1 2350
box -12 -8 74 272
use AOI22X1  _2799_
timestamp 1701862152
transform 1 0 10510 0 -1 2870
box -14 -8 114 272
use OAI21X1  _2800_
timestamp 1702508443
transform -1 0 10590 0 -1 4430
box -12 -8 92 272
use INVX1  _2801_
timestamp 1701862152
transform -1 0 9510 0 -1 2870
box -12 -8 52 272
use OAI21X1  _2802_
timestamp 1702508443
transform -1 0 7410 0 -1 1830
box -12 -8 92 272
use OAI22X1  _2803_
timestamp 1701862152
transform 1 0 8530 0 -1 2870
box -12 -8 112 272
use OAI21X1  _2804_
timestamp 1702508443
transform -1 0 9670 0 -1 3390
box -12 -8 92 272
use AND2X2  _2805_
timestamp 1701862152
transform -1 0 9970 0 -1 2870
box -12 -8 94 272
use NOR2X1  _2806_
timestamp 1701862152
transform 1 0 9670 0 -1 2870
box -12 -8 74 272
use AOI22X1  _2807_
timestamp 1701862152
transform 1 0 9010 0 -1 2350
box -14 -8 114 272
use OAI21X1  _2808_
timestamp 1702508443
transform 1 0 8770 0 -1 2350
box -12 -8 92 272
use NAND2X1  _2809_
timestamp 1702508443
transform 1 0 10490 0 1 2350
box -12 -8 72 272
use OAI22X1  _2810_
timestamp 1701862152
transform -1 0 10330 0 1 2350
box -12 -8 112 272
use OAI21X1  _2811_
timestamp 1702508443
transform 1 0 5050 0 -1 4430
box -12 -8 92 272
use NAND2X1  _2812_
timestamp 1702508443
transform -1 0 9050 0 1 4950
box -12 -8 72 272
use NOR2X1  _2813_
timestamp 1701862152
transform 1 0 9110 0 1 3390
box -12 -8 74 272
use INVX1  _2814_
timestamp 1701862152
transform -1 0 8950 0 -1 4430
box -12 -8 52 272
use NAND3X1  _2815_
timestamp 1702508443
transform -1 0 8770 0 1 3910
box -12 -8 92 272
use NAND2X1  _2816_
timestamp 1702508443
transform -1 0 8370 0 1 4950
box -12 -8 72 272
use OAI21X1  _2817_
timestamp 1702508443
transform 1 0 8750 0 1 4950
box -12 -8 92 272
use INVX1  _2818_
timestamp 1701862152
transform 1 0 8470 0 -1 4430
box -12 -8 52 272
use OAI21X1  _2819_
timestamp 1702508443
transform 1 0 8670 0 -1 4430
box -12 -8 92 272
use INVX1  _2820_
timestamp 1701862152
transform -1 0 9650 0 1 2350
box -12 -8 52 272
use AOI22X1  _2821_
timestamp 1701862152
transform 1 0 9150 0 1 2350
box -14 -8 114 272
use NAND3X1  _2822_
timestamp 1702508443
transform -1 0 9210 0 1 1830
box -12 -8 92 272
use OAI21X1  _2823_
timestamp 1702508443
transform -1 0 8990 0 1 2350
box -12 -8 92 272
use OAI21X1  _2824_
timestamp 1702508443
transform 1 0 10050 0 -1 3390
box -12 -8 92 272
use OAI21X1  _2825_
timestamp 1702508443
transform -1 0 10810 0 -1 3390
box -12 -8 92 272
use INVX1  _2826_
timestamp 1701862152
transform 1 0 9630 0 1 790
box -12 -8 52 272
use NAND3X1  _2827_
timestamp 1702508443
transform -1 0 9430 0 -1 1830
box -12 -8 92 272
use OAI21X1  _2828_
timestamp 1702508443
transform 1 0 7090 0 -1 1830
box -12 -8 92 272
use INVX1  _2829_
timestamp 1701862152
transform -1 0 10130 0 1 2870
box -12 -8 52 272
use OAI21X1  _2830_
timestamp 1702508443
transform 1 0 8410 0 -1 3390
box -12 -8 92 272
use OAI21X1  _2831_
timestamp 1702508443
transform 1 0 8450 0 1 3910
box -12 -8 92 272
use NOR2X1  _2832_
timestamp 1701862152
transform -1 0 9450 0 1 2350
box -12 -8 74 272
use OAI21X1  _2833_
timestamp 1702508443
transform -1 0 9430 0 -1 3390
box -12 -8 92 272
use OAI21X1  _2834_
timestamp 1702508443
transform -1 0 9190 0 -1 3390
box -12 -8 92 272
use NOR2X1  _2835_
timestamp 1701862152
transform -1 0 9470 0 1 790
box -12 -8 74 272
use OAI21X1  _2836_
timestamp 1702508443
transform 1 0 9010 0 1 1310
box -12 -8 92 272
use AOI21X1  _2837_
timestamp 1702508443
transform -1 0 9750 0 1 1310
box -12 -8 92 272
use OAI21X1  _2838_
timestamp 1702508443
transform -1 0 9870 0 1 3390
box -12 -8 92 272
use OAI21X1  _2839_
timestamp 1702508443
transform -1 0 9890 0 -1 3390
box -12 -8 92 272
use NAND2X1  _2840_
timestamp 1702508443
transform 1 0 9170 0 -1 270
box -12 -8 72 272
use NAND2X1  _2841_
timestamp 1702508443
transform -1 0 9010 0 -1 270
box -12 -8 72 272
use OAI21X1  _2842_
timestamp 1702508443
transform 1 0 9390 0 -1 270
box -12 -8 92 272
use NAND2X1  _2843_
timestamp 1702508443
transform 1 0 9630 0 -1 270
box -12 -8 72 272
use NOR2X1  _2844_
timestamp 1701862152
transform 1 0 9430 0 1 270
box -12 -8 74 272
use AND2X2  _2845_
timestamp 1701862152
transform -1 0 10170 0 1 270
box -12 -8 94 272
use OAI21X1  _2846_
timestamp 1702508443
transform 1 0 9850 0 1 270
box -12 -8 92 272
use NAND2X1  _2847_
timestamp 1702508443
transform -1 0 11270 0 -1 10670
box -12 -8 72 272
use NAND2X1  _2848_
timestamp 1702508443
transform -1 0 10770 0 -1 1310
box -12 -8 72 272
use INVX1  _2849_
timestamp 1701862152
transform -1 0 11090 0 1 1310
box -12 -8 52 272
use OAI21X1  _2850_
timestamp 1702508443
transform -1 0 11270 0 -1 1830
box -12 -8 92 272
use OAI21X1  _2851_
timestamp 1702508443
transform 1 0 10810 0 -1 3910
box -12 -8 92 272
use NAND2X1  _2852_
timestamp 1702508443
transform -1 0 9050 0 1 270
box -12 -8 72 272
use NOR2X1  _2853_
timestamp 1701862152
transform -1 0 9270 0 1 270
box -12 -8 74 272
use INVX1  _2854_
timestamp 1701862152
transform 1 0 10710 0 1 790
box -12 -8 52 272
use NOR2X1  _2855_
timestamp 1701862152
transform -1 0 9970 0 1 1310
box -12 -8 74 272
use NAND3X1  _2856_
timestamp 1702508443
transform -1 0 10650 0 1 1310
box -12 -8 92 272
use NAND3X1  _2857_
timestamp 1702508443
transform -1 0 10890 0 1 1310
box -12 -8 92 272
use OAI21X1  _2858_
timestamp 1702508443
transform -1 0 11250 0 1 1830
box -12 -8 92 272
use OAI21X1  _2859_
timestamp 1702508443
transform 1 0 11050 0 -1 3910
box -12 -8 92 272
use INVX1  _2860_
timestamp 1701862152
transform 1 0 10970 0 -1 3390
box -12 -8 52 272
use NAND2X1  _2861_
timestamp 1702508443
transform 1 0 9830 0 -1 270
box -12 -8 72 272
use OAI21X1  _2862_
timestamp 1702508443
transform 1 0 8710 0 -1 270
box -12 -8 92 272
use OAI22X1  _2863_
timestamp 1701862152
transform -1 0 10430 0 1 270
box -12 -8 112 272
use NAND2X1  _2864_
timestamp 1702508443
transform 1 0 10590 0 1 270
box -12 -8 72 272
use OAI21X1  _2865_
timestamp 1702508443
transform -1 0 10890 0 1 270
box -12 -8 92 272
use OAI21X1  _2866_
timestamp 1702508443
transform -1 0 11270 0 -1 790
box -12 -8 92 272
use OAI21X1  _2867_
timestamp 1702508443
transform 1 0 11170 0 -1 3390
box -12 -8 92 272
use INVX1  _2868_
timestamp 1701862152
transform 1 0 11130 0 1 790
box -12 -8 52 272
use INVX1  _2869_
timestamp 1701862152
transform 1 0 10270 0 1 790
box -12 -8 52 272
use AOI22X1  _2870_
timestamp 1701862152
transform -1 0 10570 0 1 790
box -14 -8 114 272
use NAND3X1  _2871_
timestamp 1702508443
transform -1 0 10990 0 1 790
box -12 -8 92 272
use INVX1  _2872_
timestamp 1701862152
transform -1 0 11290 0 1 1310
box -12 -8 52 272
use OAI21X1  _2873_
timestamp 1702508443
transform -1 0 10110 0 1 3390
box -12 -8 92 272
use OAI21X1  _2874_
timestamp 1702508443
transform -1 0 10350 0 1 3390
box -12 -8 92 272
use INVX1  _2875_
timestamp 1701862152
transform -1 0 10890 0 -1 4950
box -12 -8 52 272
use NAND2X1  _2876_
timestamp 1702508443
transform -1 0 9850 0 1 1830
box -12 -8 72 272
use OAI21X1  _2877_
timestamp 1702508443
transform 1 0 10010 0 1 1830
box -12 -8 92 272
use NOR2X1  _2878_
timestamp 1701862152
transform 1 0 9830 0 -1 1310
box -12 -8 74 272
use NAND3X1  _2879_
timestamp 1702508443
transform -1 0 10130 0 -1 1310
box -12 -8 92 272
use NAND3X1  _2880_
timestamp 1702508443
transform 1 0 9570 0 1 1830
box -12 -8 92 272
use OAI21X1  _2881_
timestamp 1702508443
transform 1 0 10950 0 -1 790
box -12 -8 92 272
use NOR2X1  _2882_
timestamp 1701862152
transform -1 0 9670 0 -1 1310
box -12 -8 74 272
use NAND2X1  _2883_
timestamp 1702508443
transform -1 0 10550 0 -1 1310
box -12 -8 72 272
use NAND3X1  _2884_
timestamp 1702508443
transform 1 0 11170 0 -1 1310
box -12 -8 92 272
use OR2X2  _2885_
timestamp 1702508443
transform -1 0 11010 0 -1 1310
box -12 -8 92 272
use OAI21X1  _2886_
timestamp 1702508443
transform 1 0 10710 0 1 1830
box -12 -8 92 272
use OAI21X1  _2887_
timestamp 1702508443
transform 1 0 10270 0 -1 4430
box -12 -8 92 272
use NOR2X1  _2888_
timestamp 1701862152
transform -1 0 4130 0 1 5470
box -12 -8 74 272
use OAI21X1  _2889_
timestamp 1702508443
transform 1 0 6210 0 1 2350
box -12 -8 92 272
use NOR2X1  _2890_
timestamp 1701862152
transform -1 0 8510 0 1 5990
box -12 -8 74 272
use INVX2  _2891_
timestamp 1701862152
transform -1 0 8310 0 1 5990
box -12 -8 52 272
use OAI21X1  _2892_
timestamp 1702508443
transform 1 0 7510 0 -1 5470
box -12 -8 92 272
use OAI21X1  _2893_
timestamp 1702508443
transform 1 0 7330 0 1 5470
box -12 -8 92 272
use OAI21X1  _2894_
timestamp 1702508443
transform 1 0 6610 0 -1 6510
box -12 -8 92 272
use OAI21X1  _2895_
timestamp 1702508443
transform 1 0 6750 0 1 6510
box -12 -8 92 272
use OAI21X1  _2896_
timestamp 1702508443
transform -1 0 8070 0 -1 5470
box -12 -8 92 272
use OAI21X1  _2897_
timestamp 1702508443
transform 1 0 7790 0 1 5470
box -12 -8 92 272
use OAI21X1  _2898_
timestamp 1702508443
transform 1 0 7330 0 -1 6510
box -12 -8 92 272
use OAI21X1  _2899_
timestamp 1702508443
transform 1 0 6850 0 -1 6510
box -12 -8 92 272
use OAI21X1  _2900_
timestamp 1702508443
transform -1 0 6450 0 -1 6510
box -12 -8 92 272
use OAI21X1  _2901_
timestamp 1702508443
transform 1 0 6130 0 -1 6510
box -12 -8 92 272
use OAI21X1  _2902_
timestamp 1702508443
transform -1 0 8110 0 1 5990
box -12 -8 92 272
use OAI21X1  _2903_
timestamp 1702508443
transform 1 0 7330 0 1 5990
box -12 -8 92 272
use OAI21X1  _2904_
timestamp 1702508443
transform 1 0 8450 0 -1 5470
box -12 -8 92 272
use OAI21X1  _2905_
timestamp 1702508443
transform 1 0 8450 0 1 5470
box -12 -8 92 272
use OAI21X1  _2906_
timestamp 1702508443
transform 1 0 8210 0 -1 5990
box -12 -8 92 272
use OAI21X1  _2907_
timestamp 1702508443
transform -1 0 8050 0 -1 5990
box -12 -8 92 272
use OAI21X1  _2908_
timestamp 1702508443
transform -1 0 8370 0 -1 4950
box -12 -8 92 272
use OAI21X1  _2909_
timestamp 1702508443
transform 1 0 3450 0 -1 4430
box -12 -8 92 272
use AOI21X1  _2910_
timestamp 1702508443
transform -1 0 6670 0 -1 4430
box -12 -8 92 272
use NOR2X1  _2911_
timestamp 1701862152
transform -1 0 6990 0 1 4430
box -12 -8 74 272
use NOR2X1  _2912_
timestamp 1701862152
transform 1 0 8710 0 -1 4950
box -12 -8 74 272
use AOI21X1  _2913_
timestamp 1702508443
transform -1 0 6970 0 -1 4950
box -12 -8 92 272
use INVX1  _2914_
timestamp 1701862152
transform 1 0 7170 0 -1 8070
box -12 -8 52 272
use NAND3X1  _2915_
timestamp 1702508443
transform 1 0 7290 0 -1 5990
box -12 -8 92 272
use OAI21X1  _2916_
timestamp 1702508443
transform 1 0 7050 0 -1 5990
box -12 -8 92 272
use NAND2X1  _2917_
timestamp 1702508443
transform -1 0 6470 0 -1 5990
box -12 -8 72 272
use OAI21X1  _2918_
timestamp 1702508443
transform 1 0 6350 0 1 5470
box -12 -8 92 272
use NAND2X1  _2919_
timestamp 1702508443
transform 1 0 6250 0 1 4950
box -12 -8 72 272
use OAI21X1  _2920_
timestamp 1702508443
transform 1 0 6030 0 1 4950
box -12 -8 92 272
use NOR2X1  _2921_
timestamp 1701862152
transform -1 0 7530 0 -1 3910
box -12 -8 74 272
use NAND2X1  _2922_
timestamp 1702508443
transform -1 0 7570 0 1 3910
box -12 -8 72 272
use OAI21X1  _2923_
timestamp 1702508443
transform -1 0 6910 0 -1 4430
box -12 -8 92 272
use NAND2X1  _2924_
timestamp 1702508443
transform 1 0 6470 0 1 4950
box -12 -8 72 272
use INVX1  _2925_
timestamp 1701862152
transform 1 0 7370 0 1 7550
box -12 -8 52 272
use INVX1  _2926_
timestamp 1701862152
transform -1 0 7630 0 1 4430
box -12 -8 52 272
use OAI21X1  _2927_
timestamp 1702508443
transform 1 0 7370 0 -1 4950
box -12 -8 92 272
use MUX2X1  _2928_
timestamp 1701862152
transform 1 0 7130 0 -1 4950
box -12 -8 114 272
use OAI21X1  _2929_
timestamp 1702508443
transform -1 0 6770 0 1 4950
box -12 -8 92 272
use NOR2X1  _2930_
timestamp 1701862152
transform 1 0 6250 0 1 1830
box -12 -8 74 272
use NAND2X1  _2931_
timestamp 1702508443
transform 1 0 7130 0 -1 2870
box -12 -8 72 272
use INVX1  _2932_
timestamp 1701862152
transform 1 0 5290 0 -1 4430
box -12 -8 52 272
use AOI21X1  _2933_
timestamp 1702508443
transform 1 0 5490 0 -1 4430
box -12 -8 92 272
use OAI21X1  _2934_
timestamp 1702508443
transform 1 0 5710 0 -1 4430
box -12 -8 92 272
use INVX1  _2935_
timestamp 1701862152
transform 1 0 6550 0 1 6510
box -12 -8 52 272
use NOR2X1  _2936_
timestamp 1701862152
transform 1 0 6430 0 -1 4950
box -12 -8 74 272
use OAI21X1  _2937_
timestamp 1702508443
transform 1 0 6650 0 -1 4950
box -12 -8 92 272
use OAI21X1  _2938_
timestamp 1702508443
transform 1 0 5130 0 1 4950
box -12 -8 92 272
use NOR2X1  _2939_
timestamp 1701862152
transform 1 0 4910 0 1 4950
box -12 -8 74 272
use NAND2X1  _2940_
timestamp 1702508443
transform -1 0 6010 0 -1 5470
box -12 -8 72 272
use OAI21X1  _2941_
timestamp 1702508443
transform 1 0 5710 0 -1 5470
box -12 -8 92 272
use OAI21X1  _2942_
timestamp 1702508443
transform -1 0 9490 0 1 4430
box -12 -8 92 272
use INVX1  _2943_
timestamp 1701862152
transform 1 0 6390 0 -1 4430
box -12 -8 52 272
use NOR2X1  _2944_
timestamp 1701862152
transform -1 0 6450 0 1 3910
box -12 -8 74 272
use AOI22X1  _2945_
timestamp 1701862152
transform -1 0 6570 0 1 4430
box -14 -8 114 272
use NOR2X1  _2946_
timestamp 1701862152
transform 1 0 6250 0 1 4430
box -12 -8 74 272
use OAI21X1  _2947_
timestamp 1702508443
transform -1 0 6710 0 -1 5990
box -12 -8 92 272
use OAI21X1  _2948_
timestamp 1702508443
transform 1 0 6170 0 -1 5990
box -12 -8 92 272
use INVX1  _2949_
timestamp 1701862152
transform -1 0 6030 0 -1 5990
box -12 -8 52 272
use OAI21X1  _2950_
timestamp 1702508443
transform 1 0 5870 0 1 5470
box -12 -8 92 272
use OAI21X1  _2951_
timestamp 1702508443
transform -1 0 6190 0 1 5470
box -12 -8 92 272
use AOI21X1  _2952_
timestamp 1702508443
transform -1 0 6270 0 -1 4950
box -12 -8 92 272
use INVX1  _2953_
timestamp 1701862152
transform -1 0 4510 0 1 4950
box -12 -8 52 272
use INVX1  _2954_
timestamp 1701862152
transform -1 0 6770 0 1 4430
box -12 -8 52 272
use AND2X2  _2955_
timestamp 1701862152
transform -1 0 6090 0 1 4430
box -12 -8 94 272
use AOI22X1  _2956_
timestamp 1701862152
transform 1 0 5290 0 1 4430
box -14 -8 114 272
use OAI21X1  _2957_
timestamp 1702508443
transform 1 0 5250 0 -1 4950
box -12 -8 92 272
use NAND2X1  _2958_
timestamp 1702508443
transform -1 0 5610 0 1 4430
box -12 -8 72 272
use INVX1  _2959_
timestamp 1701862152
transform 1 0 7070 0 -1 5470
box -12 -8 52 272
use MUX2X1  _2960_
timestamp 1701862152
transform -1 0 6690 0 1 5470
box -12 -8 114 272
use AOI21X1  _2961_
timestamp 1702508443
transform 1 0 6370 0 -1 5470
box -12 -8 92 272
use OAI21X1  _2962_
timestamp 1702508443
transform -1 0 6690 0 -1 5470
box -12 -8 92 272
use OAI21X1  _2963_
timestamp 1702508443
transform -1 0 6910 0 -1 5470
box -12 -8 92 272
use NAND3X1  _2964_
timestamp 1702508443
transform -1 0 5570 0 -1 4950
box -12 -8 92 272
use OAI21X1  _2965_
timestamp 1702508443
transform 1 0 5010 0 -1 4950
box -12 -8 92 272
use NOR2X1  _2966_
timestamp 1701862152
transform -1 0 6510 0 1 2350
box -12 -8 74 272
use NAND3X1  _2967_
timestamp 1702508443
transform 1 0 7730 0 1 3910
box -12 -8 92 272
use NOR2X1  _2968_
timestamp 1701862152
transform -1 0 7090 0 -1 3910
box -12 -8 74 272
use NAND2X1  _2969_
timestamp 1702508443
transform -1 0 7310 0 -1 3910
box -12 -8 72 272
use OR2X2  _2970_
timestamp 1702508443
transform -1 0 7350 0 1 3910
box -12 -8 92 272
use OAI21X1  _2971_
timestamp 1702508443
transform -1 0 6890 0 1 3910
box -12 -8 92 272
use AOI21X1  _2972_
timestamp 1702508443
transform 1 0 7050 0 1 3910
box -12 -8 92 272
use NAND2X1  _2973_
timestamp 1702508443
transform -1 0 7210 0 1 4430
box -12 -8 72 272
use AOI21X1  _2974_
timestamp 1702508443
transform 1 0 7070 0 -1 4430
box -12 -8 92 272
use NAND2X1  _2975_
timestamp 1702508443
transform -1 0 7870 0 -1 4430
box -12 -8 72 272
use OAI21X1  _2976_
timestamp 1702508443
transform -1 0 7650 0 -1 4430
box -12 -8 92 272
use MUX2X1  _2977_
timestamp 1701862152
transform 1 0 7310 0 -1 4430
box -12 -8 114 272
use OAI21X1  _2978_
timestamp 1702508443
transform 1 0 7350 0 1 4430
box -12 -8 92 272
use INVX1  _2979_
timestamp 1701862152
transform -1 0 3730 0 -1 4950
box -12 -8 52 272
use NAND2X1  _2980_
timestamp 1702508443
transform -1 0 3130 0 1 7550
box -12 -8 72 272
use OAI21X1  _2981_
timestamp 1702508443
transform 1 0 3610 0 1 4950
box -12 -8 92 272
use NAND2X1  _2982_
timestamp 1702508443
transform 1 0 9670 0 1 6510
box -12 -8 72 272
use OAI21X1  _2983_
timestamp 1702508443
transform 1 0 1990 0 1 4430
box -12 -8 92 272
use OAI21X1  _2984_
timestamp 1702508443
transform -1 0 3670 0 -1 3910
box -12 -8 92 272
use OR2X2  _2985_
timestamp 1702508443
transform 1 0 3750 0 1 4430
box -12 -8 92 272
use OAI21X1  _2986_
timestamp 1702508443
transform -1 0 6030 0 -1 4430
box -12 -8 92 272
use OAI21X1  _2987_
timestamp 1702508443
transform -1 0 5850 0 1 4430
box -12 -8 92 272
use NOR2X1  _2988_
timestamp 1701862152
transform 1 0 9450 0 1 6510
box -12 -8 74 272
use OAI21X1  _2989_
timestamp 1702508443
transform 1 0 6070 0 1 6510
box -12 -8 92 272
use OAI21X1  _2990_
timestamp 1702508443
transform -1 0 6390 0 1 6510
box -12 -8 92 272
use INVX1  _2991_
timestamp 1701862152
transform 1 0 7230 0 1 6510
box -12 -8 52 272
use NOR2X1  _2992_
timestamp 1701862152
transform 1 0 9730 0 1 7030
box -12 -8 74 272
use AOI21X1  _2993_
timestamp 1702508443
transform 1 0 9950 0 1 7030
box -12 -8 92 272
use NOR2X1  _2994_
timestamp 1701862152
transform -1 0 10910 0 -1 7550
box -12 -8 74 272
use NAND3X1  _2995_
timestamp 1702508443
transform -1 0 7730 0 -1 7550
box -12 -8 92 272
use NOR2X1  _2996_
timestamp 1701862152
transform 1 0 7570 0 1 7550
box -12 -8 74 272
use NAND2X1  _2997_
timestamp 1702508443
transform -1 0 7490 0 -1 7550
box -12 -8 72 272
use NAND2X1  _2998_
timestamp 1702508443
transform -1 0 6550 0 -1 7550
box -12 -8 72 272
use NAND2X1  _2999_
timestamp 1702508443
transform 1 0 6210 0 1 7550
box -12 -8 72 272
use INVX1  _3000_
timestamp 1701862152
transform -1 0 6090 0 -1 7550
box -12 -8 52 272
use NOR2X1  _3001_
timestamp 1701862152
transform -1 0 5890 0 -1 7550
box -12 -8 74 272
use OAI21X1  _3002_
timestamp 1702508443
transform -1 0 6330 0 -1 7550
box -12 -8 92 272
use OAI21X1  _3003_
timestamp 1702508443
transform -1 0 6510 0 1 7550
box -12 -8 92 272
use INVX1  _3004_
timestamp 1701862152
transform 1 0 8250 0 1 7550
box -12 -8 52 272
use AOI21X1  _3005_
timestamp 1702508443
transform 1 0 11070 0 -1 7550
box -12 -8 92 272
use NOR2X1  _3006_
timestamp 1701862152
transform -1 0 10590 0 1 7550
box -12 -8 74 272
use XNOR2X1  _3007_ ~/ETRI050_DesignKit/devel/Ref_Design/CPU_6502/layout/digital_ETRI
timestamp 1702508443
transform 1 0 7050 0 1 7030
box -12 -8 132 272
use NAND2X1  _3008_
timestamp 1702508443
transform -1 0 6670 0 1 7030
box -12 -8 72 272
use OAI21X1  _3009_
timestamp 1702508443
transform -1 0 6090 0 -1 7030
box -12 -8 92 272
use INVX1  _3010_
timestamp 1701862152
transform 1 0 6250 0 -1 7030
box -12 -8 52 272
use OAI21X1  _3011_
timestamp 1702508443
transform 1 0 6830 0 1 7030
box -12 -8 92 272
use OAI21X1  _3012_
timestamp 1702508443
transform -1 0 8010 0 -1 7030
box -12 -8 92 272
use INVX1  _3013_
timestamp 1701862152
transform 1 0 8390 0 -1 7030
box -12 -8 52 272
use AOI21X1  _3014_
timestamp 1702508443
transform 1 0 10730 0 1 7550
box -12 -8 92 272
use OAI21X1  _3015_
timestamp 1702508443
transform -1 0 6530 0 -1 7030
box -12 -8 92 272
use XOR2X1  _3016_
timestamp 1702508443
transform -1 0 7450 0 1 7030
box -12 -8 132 272
use XOR2X1  _3017_
timestamp 1702508443
transform 1 0 6690 0 -1 7030
box -12 -8 132 272
use OAI21X1  _3018_
timestamp 1702508443
transform -1 0 7050 0 -1 7030
box -12 -8 92 272
use OAI21X1  _3019_
timestamp 1702508443
transform -1 0 7290 0 -1 7030
box -12 -8 92 272
use INVX1  _3020_
timestamp 1701862152
transform 1 0 8390 0 1 7030
box -12 -8 52 272
use NOR2X1  _3021_
timestamp 1701862152
transform -1 0 9470 0 -1 8070
box -12 -8 74 272
use AOI21X1  _3022_
timestamp 1702508443
transform 1 0 9630 0 -1 8070
box -12 -8 92 272
use OAI21X1  _3023_
timestamp 1702508443
transform -1 0 5910 0 1 6510
box -12 -8 92 272
use OAI21X1  _3024_
timestamp 1702508443
transform 1 0 5590 0 1 6510
box -12 -8 92 272
use INVX1  _3025_
timestamp 1701862152
transform -1 0 5630 0 -1 6510
box -12 -8 52 272
use NOR2X1  _3026_
timestamp 1701862152
transform 1 0 11030 0 -1 5990
box -12 -8 74 272
use AOI21X1  _3027_
timestamp 1702508443
transform -1 0 11330 0 -1 5990
box -12 -8 92 272
use NOR2X1  _3028_
timestamp 1701862152
transform -1 0 9910 0 -1 8070
box -12 -8 74 272
use NAND3X1  _3029_
timestamp 1702508443
transform -1 0 7270 0 -1 7550
box -12 -8 92 272
use NOR2X1  _3030_
timestamp 1701862152
transform -1 0 8230 0 -1 7030
box -12 -8 74 272
use NAND2X1  _3031_
timestamp 1702508443
transform 1 0 8170 0 1 7030
box -12 -8 72 272
use NAND2X1  _3032_
timestamp 1702508443
transform 1 0 7790 0 1 7550
box -12 -8 72 272
use INVX1  _3033_
timestamp 1701862152
transform -1 0 6890 0 1 8070
box -12 -8 52 272
use INVX1  _3034_
timestamp 1701862152
transform -1 0 7870 0 -1 8070
box -12 -8 52 272
use OAI21X1  _3035_
timestamp 1702508443
transform 1 0 7590 0 -1 8070
box -12 -8 92 272
use INVX1  _3036_
timestamp 1701862152
transform -1 0 7070 0 1 8070
box -12 -8 52 272
use OAI21X1  _3037_
timestamp 1702508443
transform -1 0 6690 0 1 8070
box -12 -8 92 272
use OAI21X1  _3038_
timestamp 1702508443
transform -1 0 7310 0 1 8070
box -12 -8 92 272
use INVX1  _3039_
timestamp 1701862152
transform 1 0 7470 0 1 8070
box -12 -8 52 272
use AOI21X1  _3040_
timestamp 1702508443
transform 1 0 9810 0 1 7550
box -12 -8 92 272
use NOR2X1  _3041_
timestamp 1701862152
transform -1 0 9710 0 -1 6510
box -12 -8 74 272
use NOR2X1  _3042_
timestamp 1701862152
transform 1 0 7370 0 -1 8070
box -12 -8 74 272
use XNOR2X1  _3043_
timestamp 1702508443
transform -1 0 6770 0 1 7550
box -12 -8 132 272
use AOI21X1  _3044_
timestamp 1702508443
transform -1 0 6790 0 -1 7550
box -12 -8 92 272
use OAI21X1  _3045_
timestamp 1702508443
transform 1 0 6950 0 -1 7550
box -12 -8 92 272
use OAI21X1  _3046_
timestamp 1702508443
transform -1 0 7970 0 1 6510
box -12 -8 92 272
use INVX1  _3047_
timestamp 1701862152
transform 1 0 9250 0 1 6510
box -12 -8 52 272
use AOI21X1  _3048_
timestamp 1702508443
transform 1 0 9870 0 -1 6510
box -12 -8 92 272
use NAND2X1  _3049_
timestamp 1702508443
transform -1 0 6990 0 1 7550
box -12 -8 72 272
use OAI21X1  _3050_
timestamp 1702508443
transform -1 0 7210 0 1 7550
box -12 -8 92 272
use XNOR2X1  _3051_
timestamp 1702508443
transform -1 0 8010 0 1 7030
box -12 -8 132 272
use XOR2X1  _3052_
timestamp 1702508443
transform 1 0 7610 0 1 7030
box -12 -8 132 272
use OAI21X1  _3053_
timestamp 1702508443
transform 1 0 7450 0 -1 7030
box -12 -8 92 272
use OAI21X1  _3054_
timestamp 1702508443
transform -1 0 7770 0 -1 7030
box -12 -8 92 272
use INVX1  _3055_
timestamp 1701862152
transform 1 0 8130 0 1 6510
box -12 -8 52 272
use NOR2X1  _3056_
timestamp 1701862152
transform -1 0 9690 0 1 5470
box -12 -8 74 272
use AOI21X1  _3057_
timestamp 1702508443
transform -1 0 9470 0 1 5470
box -12 -8 92 272
use INVX2  _3058_
timestamp 1701862152
transform 1 0 8810 0 -1 7550
box -12 -8 52 272
use OR2X2  _3059_
timestamp 1702508443
transform -1 0 8770 0 -1 5990
box -12 -8 92 272
use OAI21X1  _3060_
timestamp 1702508443
transform 1 0 9890 0 1 6510
box -12 -8 92 272
use OAI21X1  _3061_
timestamp 1702508443
transform 1 0 10130 0 1 6510
box -12 -8 92 272
use OAI21X1  _3062_
timestamp 1702508443
transform -1 0 9810 0 -1 7550
box -12 -8 92 272
use OAI21X1  _3063_
timestamp 1702508443
transform 1 0 9490 0 -1 7550
box -12 -8 92 272
use OAI21X1  _3064_
timestamp 1702508443
transform -1 0 10510 0 -1 7030
box -12 -8 92 272
use OAI21X1  _3065_
timestamp 1702508443
transform -1 0 10730 0 -1 7030
box -12 -8 92 272
use OAI21X1  _3066_
timestamp 1702508443
transform -1 0 8670 0 -1 7550
box -12 -8 92 272
use OAI21X1  _3067_
timestamp 1702508443
transform 1 0 8350 0 -1 7550
box -12 -8 92 272
use OAI21X1  _3068_
timestamp 1702508443
transform 1 0 10310 0 -1 5990
box -12 -8 92 272
use OAI21X1  _3069_
timestamp 1702508443
transform 1 0 10550 0 -1 5990
box -12 -8 92 272
use OAI21X1  _3070_
timestamp 1702508443
transform 1 0 9010 0 -1 7550
box -12 -8 92 272
use OAI21X1  _3071_
timestamp 1702508443
transform -1 0 9330 0 -1 7550
box -12 -8 92 272
use OAI21X1  _3072_
timestamp 1702508443
transform -1 0 9930 0 1 5990
box -12 -8 92 272
use OAI21X1  _3073_
timestamp 1702508443
transform -1 0 10170 0 1 5990
box -12 -8 92 272
use OAI21X1  _3074_
timestamp 1702508443
transform 1 0 8930 0 1 5990
box -12 -8 92 272
use OAI21X1  _3075_
timestamp 1702508443
transform 1 0 8930 0 -1 5990
box -12 -8 92 272
use INVX1  _3076_
timestamp 1701862152
transform 1 0 10830 0 1 6510
box -12 -8 52 272
use NOR2X1  _3077_
timestamp 1701862152
transform 1 0 11030 0 1 6510
box -12 -8 74 272
use NOR2X1  _3078_
timestamp 1701862152
transform -1 0 8870 0 -1 7030
box -12 -8 74 272
use AOI21X1  _3079_
timestamp 1702508443
transform -1 0 8650 0 -1 7030
box -12 -8 92 272
use NOR2X1  _3080_
timestamp 1701862152
transform 1 0 11090 0 -1 8590
box -12 -8 74 272
use AOI21X1  _3081_
timestamp 1702508443
transform -1 0 11150 0 -1 270
box -12 -8 92 272
use NOR2X1  _3082_
timestamp 1701862152
transform 1 0 10190 0 -1 8590
box -12 -8 74 272
use AOI21X1  _3083_
timestamp 1702508443
transform -1 0 10030 0 -1 8590
box -12 -8 92 272
use NOR2X1  _3084_
timestamp 1701862152
transform -1 0 9190 0 1 7550
box -12 -8 74 272
use AOI21X1  _3085_
timestamp 1702508443
transform 1 0 9050 0 1 7030
box -12 -8 92 272
use NOR2X1  _3086_
timestamp 1701862152
transform -1 0 10850 0 1 5990
box -12 -8 74 272
use AOI21X1  _3087_
timestamp 1702508443
transform 1 0 10990 0 1 5990
box -12 -8 92 272
use NOR2X1  _3088_
timestamp 1701862152
transform 1 0 8370 0 1 8070
box -12 -8 74 272
use AOI21X1  _3089_
timestamp 1702508443
transform -1 0 8210 0 1 8070
box -12 -8 92 272
use NOR2X1  _3090_
timestamp 1701862152
transform -1 0 11290 0 1 4950
box -12 -8 74 272
use AOI21X1  _3091_
timestamp 1702508443
transform 1 0 10990 0 1 4950
box -12 -8 92 272
use NOR2X1  _3092_
timestamp 1701862152
transform 1 0 8910 0 -1 5470
box -12 -8 74 272
use AOI21X1  _3093_
timestamp 1702508443
transform -1 0 9210 0 -1 5470
box -12 -8 92 272
use INVX1  _3094_
timestamp 1701862152
transform -1 0 10350 0 -1 5470
box -12 -8 52 272
use NOR2X1  _3095_
timestamp 1701862152
transform 1 0 10290 0 1 5470
box -12 -8 74 272
use NOR2X1  _3096_
timestamp 1701862152
transform 1 0 9030 0 1 6510
box -12 -8 74 272
use AOI21X1  _3097_
timestamp 1702508443
transform -1 0 8870 0 1 6510
box -12 -8 92 272
use NOR2X1  _3098_
timestamp 1701862152
transform -1 0 10550 0 1 8070
box -12 -8 74 272
use AOI21X1  _3099_
timestamp 1702508443
transform -1 0 11330 0 -1 8070
box -12 -8 92 272
use NOR2X1  _3100_
timestamp 1701862152
transform 1 0 10270 0 1 8070
box -12 -8 74 272
use AOI21X1  _3101_
timestamp 1702508443
transform 1 0 10390 0 -1 8590
box -12 -8 92 272
use NOR2X1  _3102_
timestamp 1701862152
transform 1 0 8490 0 -1 8070
box -12 -8 74 272
use AOI21X1  _3103_
timestamp 1702508443
transform -1 0 8530 0 1 7550
box -12 -8 92 272
use NOR2X1  _3104_
timestamp 1701862152
transform -1 0 11310 0 1 6510
box -12 -8 74 272
use AOI21X1  _3105_
timestamp 1702508443
transform -1 0 11130 0 -1 4950
box -12 -8 92 272
use NOR2X1  _3106_
timestamp 1701862152
transform 1 0 9490 0 -1 8590
box -12 -8 74 272
use AOI21X1  _3107_
timestamp 1702508443
transform -1 0 9790 0 -1 8590
box -12 -8 92 272
use NOR2X1  _3108_
timestamp 1701862152
transform 1 0 10070 0 1 5470
box -12 -8 74 272
use AOI21X1  _3109_
timestamp 1702508443
transform -1 0 9930 0 1 5470
box -12 -8 92 272
use NOR2X1  _3110_
timestamp 1701862152
transform 1 0 8510 0 -1 6510
box -12 -8 74 272
use AOI21X1  _3111_
timestamp 1702508443
transform -1 0 8350 0 -1 6510
box -12 -8 92 272
use OAI21X1  _3112_
timestamp 1702508443
transform 1 0 630 0 -1 2870
box -12 -8 92 272
use OAI21X1  _3113_
timestamp 1702508443
transform 1 0 170 0 -1 2870
box -12 -8 92 272
use NAND2X1  _3114_
timestamp 1702508443
transform -1 0 470 0 -1 2870
box -12 -8 72 272
use OAI21X1  _3115_
timestamp 1702508443
transform -1 0 1370 0 1 2350
box -12 -8 92 272
use NOR2X1  _3116_
timestamp 1701862152
transform 1 0 1050 0 -1 2350
box -12 -8 74 272
use NOR2X1  _3117_
timestamp 1701862152
transform 1 0 2150 0 -1 1310
box -12 -8 74 272
use AOI21X1  _3118_
timestamp 1702508443
transform -1 0 1590 0 -1 2350
box -12 -8 92 272
use AND2X2  _3119_
timestamp 1701862152
transform -1 0 1350 0 -1 2350
box -12 -8 94 272
use NAND3X1  _3120_
timestamp 1702508443
transform -1 0 650 0 1 2350
box -12 -8 92 272
use NOR2X1  _3121_
timestamp 1701862152
transform 1 0 370 0 1 2870
box -12 -8 74 272
use OAI21X1  _3122_
timestamp 1702508443
transform 1 0 2630 0 -1 3390
box -12 -8 92 272
use OAI21X1  _3123_
timestamp 1702508443
transform 1 0 630 0 1 3390
box -12 -8 92 272
use AND2X2  _3124_
timestamp 1701862152
transform -1 0 490 0 1 3390
box -12 -8 94 272
use NAND3X1  _3125_
timestamp 1702508443
transform -1 0 910 0 -1 2350
box -12 -8 92 272
use OAI21X1  _3126_
timestamp 1702508443
transform -1 0 1610 0 1 2350
box -12 -8 92 272
use OR2X2  _3127_
timestamp 1702508443
transform -1 0 1130 0 1 2350
box -12 -8 92 272
use AOI22X1  _3128_
timestamp 1701862152
transform -1 0 2090 0 1 2350
box -14 -8 114 272
use NOR2X1  _3129_
timestamp 1701862152
transform -1 0 1810 0 -1 2350
box -12 -8 74 272
use NAND3X1  _3130_
timestamp 1702508443
transform -1 0 1830 0 1 2350
box -12 -8 92 272
use OAI21X1  _3131_
timestamp 1702508443
transform -1 0 890 0 1 2350
box -12 -8 92 272
use INVX1  _3132_
timestamp 1701862152
transform 1 0 590 0 1 2870
box -12 -8 52 272
use OAI21X1  _3133_
timestamp 1702508443
transform 1 0 650 0 -1 3910
box -12 -8 92 272
use NAND3X1  _3134_
timestamp 1702508443
transform -1 0 1390 0 1 3390
box -12 -8 92 272
use NOR2X1  _3135_
timestamp 1701862152
transform 1 0 1090 0 1 3390
box -12 -8 74 272
use AND2X2  _3136_
timestamp 1701862152
transform -1 0 730 0 -1 3390
box -12 -8 94 272
use AOI22X1  _3137_
timestamp 1701862152
transform 1 0 390 0 -1 3390
box -14 -8 114 272
use AOI21X1  _3138_
timestamp 1702508443
transform -1 0 1830 0 1 4430
box -12 -8 92 272
use OAI21X1  _3139_
timestamp 1702508443
transform -1 0 2050 0 -1 3390
box -12 -8 92 272
use NOR2X1  _3140_
timestamp 1701862152
transform -1 0 450 0 1 3910
box -12 -8 74 272
use AND2X2  _3141_
timestamp 1701862152
transform 1 0 850 0 1 4430
box -12 -8 94 272
use INVX1  _3142_
timestamp 1701862152
transform 1 0 1090 0 1 4430
box -12 -8 52 272
use NOR2X1  _3143_
timestamp 1701862152
transform 1 0 1110 0 -1 4430
box -12 -8 74 272
use OAI21X1  _3144_
timestamp 1702508443
transform -1 0 1410 0 -1 4430
box -12 -8 92 272
use OAI21X1  _3145_
timestamp 1702508443
transform -1 0 670 0 1 3910
box -12 -8 92 272
use INVX1  _3146_
timestamp 1701862152
transform -1 0 870 0 1 3910
box -12 -8 52 272
use AND2X2  _3147_
timestamp 1701862152
transform 1 0 630 0 -1 4430
box -12 -8 94 272
use NAND3X1  _3148_
timestamp 1702508443
transform -1 0 950 0 -1 4430
box -12 -8 92 272
use OAI21X1  _3149_
timestamp 1702508443
transform -1 0 250 0 -1 3910
box -12 -8 92 272
use OAI21X1  _3150_
timestamp 1702508443
transform -1 0 1110 0 1 3910
box -12 -8 92 272
use NOR2X1  _3151_
timestamp 1701862152
transform 1 0 170 0 1 3910
box -12 -8 74 272
use AND2X2  _3152_
timestamp 1701862152
transform 1 0 150 0 -1 4430
box -12 -8 94 272
use NAND3X1  _3153_
timestamp 1702508443
transform -1 0 470 0 -1 4430
box -12 -8 92 272
use OAI21X1  _3154_
timestamp 1702508443
transform -1 0 970 0 -1 3390
box -12 -8 92 272
use INVX1  _3155_
timestamp 1701862152
transform -1 0 210 0 1 2870
box -12 -8 52 272
use NOR2X1  _3156_
timestamp 1701862152
transform 1 0 170 0 -1 3390
box -12 -8 74 272
use NAND3X1  _3157_
timestamp 1702508443
transform -1 0 250 0 1 3390
box -12 -8 92 272
use NOR2X1  _3158_
timestamp 1701862152
transform 1 0 170 0 1 4430
box -12 -8 74 272
use AOI21X1  _3159_
timestamp 1702508443
transform 1 0 370 0 1 4430
box -12 -8 92 272
use OAI21X1  _3160_
timestamp 1702508443
transform -1 0 690 0 1 4430
box -12 -8 92 272
use NAND2X1  _3161_
timestamp 1702508443
transform 1 0 4270 0 -1 7030
box -12 -8 72 272
use OAI21X1  _3162_
timestamp 1702508443
transform -1 0 4570 0 -1 7030
box -12 -8 92 272
use NAND2X1  _3163_
timestamp 1702508443
transform 1 0 4730 0 -1 7030
box -12 -8 72 272
use OAI21X1  _3164_
timestamp 1702508443
transform 1 0 4970 0 1 7030
box -12 -8 92 272
use NAND2X1  _3165_
timestamp 1702508443
transform 1 0 4230 0 1 7550
box -12 -8 72 272
use OAI21X1  _3166_
timestamp 1702508443
transform -1 0 4530 0 1 7550
box -12 -8 92 272
use NAND2X1  _3167_
timestamp 1702508443
transform 1 0 4930 0 -1 10150
box -12 -8 72 272
use OAI21X1  _3168_
timestamp 1702508443
transform 1 0 5150 0 -1 10150
box -12 -8 92 272
use NAND2X1  _3169_
timestamp 1702508443
transform -1 0 3830 0 -1 10670
box -12 -8 72 272
use OAI21X1  _3170_
timestamp 1702508443
transform -1 0 4070 0 -1 10670
box -12 -8 92 272
use NAND2X1  _3171_
timestamp 1702508443
transform 1 0 4430 0 -1 10670
box -12 -8 72 272
use OAI21X1  _3172_
timestamp 1702508443
transform -1 0 4730 0 -1 10670
box -12 -8 92 272
use NAND2X1  _3173_
timestamp 1702508443
transform 1 0 4270 0 1 10150
box -12 -8 72 272
use OAI21X1  _3174_
timestamp 1702508443
transform -1 0 4550 0 1 10150
box -12 -8 92 272
use NAND2X1  _3175_
timestamp 1702508443
transform 1 0 5610 0 1 10150
box -12 -8 72 272
use OAI21X1  _3176_
timestamp 1702508443
transform 1 0 5370 0 1 10150
box -12 -8 92 272
use NOR2X1  _3177_
timestamp 1701862152
transform -1 0 1890 0 -1 5990
box -12 -8 74 272
use AOI21X1  _3178_
timestamp 1702508443
transform 1 0 2290 0 -1 5990
box -12 -8 92 272
use NOR2X1  _3179_
timestamp 1701862152
transform -1 0 1610 0 1 6510
box -12 -8 74 272
use AOI21X1  _3180_
timestamp 1702508443
transform -1 0 1850 0 1 6510
box -12 -8 92 272
use NOR2X1  _3181_
timestamp 1701862152
transform -1 0 670 0 -1 6510
box -12 -8 74 272
use AOI21X1  _3182_
timestamp 1702508443
transform -1 0 1110 0 -1 6510
box -12 -8 92 272
use NOR2X1  _3183_
timestamp 1701862152
transform 1 0 410 0 1 8070
box -12 -8 74 272
use AOI21X1  _3184_
timestamp 1702508443
transform -1 0 710 0 1 8070
box -12 -8 92 272
use NOR2X1  _3185_
timestamp 1701862152
transform -1 0 230 0 -1 8590
box -12 -8 74 272
use AOI21X1  _3186_
timestamp 1702508443
transform -1 0 250 0 1 8070
box -12 -8 92 272
use NOR2X1  _3187_
timestamp 1701862152
transform 1 0 810 0 -1 9110
box -12 -8 74 272
use AOI21X1  _3188_
timestamp 1702508443
transform 1 0 1030 0 -1 9110
box -12 -8 92 272
use NOR2X1  _3189_
timestamp 1701862152
transform 1 0 2190 0 -1 9630
box -12 -8 74 272
use AOI21X1  _3190_
timestamp 1702508443
transform 1 0 2450 0 1 9110
box -12 -8 92 272
use NOR2X1  _3191_
timestamp 1701862152
transform 1 0 1510 0 -1 9110
box -12 -8 74 272
use AOI21X1  _3192_
timestamp 1702508443
transform -1 0 1810 0 -1 9110
box -12 -8 92 272
use DFFSR  _3193_ ~/ETRI050_DesignKit/devel/Ref_Design/CPU_6502/layout/digital_ETRI
timestamp 1701862152
transform -1 0 1770 0 1 270
box -12 -8 474 272
use DFFSR  _3194_
timestamp 1701862152
transform -1 0 1310 0 -1 270
box -12 -8 474 272
use DFFSR  _3195_
timestamp 1701862152
transform -1 0 1770 0 -1 270
box -12 -8 474 272
use DFFSR  _3196_
timestamp 1701862152
transform 1 0 1770 0 -1 270
box -12 -8 474 272
use DFFSR  _3197_
timestamp 1701862152
transform -1 0 5630 0 1 1830
box -12 -8 474 272
use DFFSR  _3198_
timestamp 1701862152
transform -1 0 4910 0 -1 1830
box -12 -8 474 272
use DFFSR  _3199_
timestamp 1701862152
transform -1 0 3430 0 -1 7030
box -12 -8 474 272
use DFFSR  _3200_
timestamp 1701862152
transform -1 0 3090 0 1 8070
box -12 -8 474 272
use DFFSR  _3201_
timestamp 1701862152
transform -1 0 4870 0 1 9110
box -12 -8 474 272
use DFFSR  _3202_
timestamp 1701862152
transform 1 0 2550 0 1 9630
box -12 -8 474 272
use DFFSR  _3203_
timestamp 1701862152
transform -1 0 4190 0 -1 11190
box -12 -8 474 272
use DFFSR  _3204_
timestamp 1701862152
transform 1 0 2990 0 1 10670
box -12 -8 474 272
use DFFSR  _3205_
timestamp 1701862152
transform 1 0 1350 0 -1 10670
box -12 -8 474 272
use DFFSR  _3206_
timestamp 1701862152
transform 1 0 2530 0 -1 11190
box -12 -8 474 272
use DFFSR  _3207_
timestamp 1701862152
transform 1 0 230 0 -1 5990
box -12 -8 474 272
use DFFSR  _3208_
timestamp 1701862152
transform -1 0 1330 0 1 7030
box -12 -8 474 272
use DFFSR  _3209_
timestamp 1701862152
transform -1 0 1170 0 1 6510
box -12 -8 474 272
use DFFSR  _3210_
timestamp 1701862152
transform 1 0 2170 0 -1 7550
box -12 -8 474 272
use DFFSR  _3211_
timestamp 1701862152
transform -1 0 650 0 -1 9110
box -12 -8 474 272
use DFFSR  _3212_
timestamp 1701862152
transform 1 0 730 0 1 9630
box -12 -8 474 272
use DFFSR  _3213_
timestamp 1701862152
transform 1 0 470 0 1 10670
box -12 -8 474 272
use DFFSR  _3214_
timestamp 1701862152
transform 1 0 890 0 -1 10670
box -12 -8 474 272
use DFFSR  _3215_
timestamp 1701862152
transform -1 0 10630 0 1 4950
box -12 -8 474 272
use DFFSR  _3216_
timestamp 1701862152
transform 1 0 4670 0 -1 5470
box -12 -8 474 272
use DFFSR  _3217_
timestamp 1701862152
transform 1 0 6730 0 1 2350
box -12 -8 474 272
use DFFSR  _3218_
timestamp 1701862152
transform -1 0 6910 0 1 3390
box -12 -8 474 272
use DFFSR  _3219_
timestamp 1701862152
transform -1 0 6270 0 1 3390
box -12 -8 474 272
use DFFSR  _3220_
timestamp 1701862152
transform -1 0 8190 0 -1 3910
box -12 -8 474 272
use DFFSR  _3221_
timestamp 1701862152
transform -1 0 5710 0 1 5470
box -12 -8 474 272
use DFFSR  _3222_
timestamp 1701862152
transform -1 0 7890 0 -1 2870
box -12 -8 474 272
use DFFSR  _3223_
timestamp 1701862152
transform -1 0 8850 0 1 2870
box -12 -8 474 272
use DFFSR  _3224_
timestamp 1701862152
transform -1 0 8250 0 -1 3390
box -12 -8 474 272
use DFFSR  _3225_
timestamp 1701862152
transform -1 0 8610 0 -1 2350
box -12 -8 474 272
use DFFSR  _3226_
timestamp 1701862152
transform -1 0 6490 0 -1 1830
box -12 -8 474 272
use DFFSR  _3227_
timestamp 1701862152
transform -1 0 8310 0 1 2350
box -12 -8 474 272
use DFFSR  _3228_
timestamp 1701862152
transform -1 0 9430 0 -1 4950
box -12 -8 474 272
use DFFSR  _3229_
timestamp 1701862152
transform 1 0 6570 0 -1 2350
box -12 -8 474 272
use DFFSR  _3230_
timestamp 1701862152
transform -1 0 10690 0 1 4430
box -12 -8 474 272
use DFFSR  _3231_
timestamp 1701862152
transform 1 0 10590 0 1 2870
box -12 -8 474 272
use DFFSR  _3232_
timestamp 1701862152
transform -1 0 10590 0 -1 3390
box -12 -8 474 272
use DFFSR  _3233_
timestamp 1701862152
transform 1 0 10590 0 -1 4430
box -12 -8 474 272
use DFFSR  _3234_
timestamp 1701862152
transform -1 0 8950 0 1 3390
box -12 -8 474 272
use DFFSR  _3235_
timestamp 1701862152
transform -1 0 9730 0 1 2870
box -12 -8 474 272
use DFFSR  _3236_
timestamp 1701862152
transform 1 0 9110 0 -1 2350
box -12 -8 474 272
use DFFSR  _3237_
timestamp 1701862152
transform -1 0 10590 0 1 2870
box -12 -8 474 272
use DFFSR  _3238_
timestamp 1701862152
transform -1 0 9510 0 1 4950
box -12 -8 474 272
use DFFSR  _3239_
timestamp 1701862152
transform -1 0 8810 0 1 4430
box -12 -8 474 272
use DFFSR  _3240_
timestamp 1701862152
transform 1 0 8630 0 -1 2870
box -12 -8 474 272
use DFFSR  _3241_
timestamp 1701862152
transform -1 0 10810 0 1 3390
box -12 -8 474 272
use DFFSR  _3242_
timestamp 1701862152
transform 1 0 7630 0 -1 1830
box -12 -8 474 272
use DFFSR  _3243_
timestamp 1701862152
transform -1 0 8950 0 -1 3390
box -12 -8 474 272
use DFFSR  _3244_
timestamp 1701862152
transform 1 0 9170 0 1 3390
box -12 -8 474 272
use DFFSR  _3245_
timestamp 1701862152
transform -1 0 10570 0 1 3910
box -12 -8 474 272
use DFFSR  _3246_
timestamp 1701862152
transform -1 0 11030 0 1 3910
box -12 -8 474 272
use DFFSR  _3247_
timestamp 1701862152
transform -1 0 11270 0 1 3390
box -12 -8 474 272
use DFFSR  _3248_
timestamp 1701862152
transform -1 0 10390 0 -1 3910
box -12 -8 474 272
use DFFSR  _3249_
timestamp 1701862152
transform -1 0 10570 0 -1 270
box -12 -8 474 272
use DFFSR  _3250_
timestamp 1701862152
transform 1 0 6230 0 -1 3390
box -12 -8 474 272
use DFFSR  _3251_
timestamp 1701862152
transform -1 0 7010 0 -1 8070
box -12 -8 474 272
use DFFSR  _3252_
timestamp 1701862152
transform -1 0 470 0 1 5470
box -12 -8 474 272
use DFFSR  _3253_
timestamp 1701862152
transform -1 0 470 0 1 10670
box -12 -8 474 272
use DFFSR  _3254_
timestamp 1701862152
transform -1 0 670 0 -1 7030
box -12 -8 474 272
use DFFSR  _3255_
timestamp 1701862152
transform 1 0 430 0 -1 11190
box -12 -8 474 272
use DFFSR  _3256_
timestamp 1701862152
transform 1 0 1130 0 1 10670
box -12 -8 474 272
use DFFSR  _3257_
timestamp 1701862152
transform 1 0 1590 0 1 9110
box -12 -8 474 272
use DFFSR  _3258_
timestamp 1701862152
transform -1 0 4490 0 -1 5990
box -12 -8 474 272
use DFFPOSX1  _3259_ ~/ETRI050_DesignKit/devel/Ref_Design/CPU_6502/layout/digital_ETRI
timestamp 1702508443
transform 1 0 7410 0 1 5470
box -13 -8 253 272
use DFFPOSX1  _3260_
timestamp 1702508443
transform -1 0 7070 0 1 6510
box -13 -8 253 272
use DFFPOSX1  _3261_
timestamp 1702508443
transform 1 0 7590 0 -1 5470
box -13 -8 253 272
use DFFPOSX1  _3262_
timestamp 1702508443
transform 1 0 6930 0 -1 6510
box -13 -8 253 272
use DFFPOSX1  _3263_
timestamp 1702508443
transform 1 0 6090 0 1 5990
box -13 -8 253 272
use DFFPOSX1  _3264_
timestamp 1702508443
transform 1 0 7410 0 1 5990
box -13 -8 253 272
use DFFPOSX1  _3265_
timestamp 1702508443
transform -1 0 8770 0 1 5470
box -13 -8 253 272
use DFFPOSX1  _3266_
timestamp 1702508443
transform -1 0 8530 0 -1 5990
box -13 -8 253 272
use DFFSR  _3267_
timestamp 1701862152
transform -1 0 7690 0 1 4950
box -12 -8 474 272
use DFFSR  _3268_
timestamp 1701862152
transform 1 0 5210 0 1 4950
box -12 -8 474 272
use DFFSR  _3269_
timestamp 1701862152
transform 1 0 6770 0 1 4950
box -12 -8 474 272
use DFFSR  _3270_
timestamp 1701862152
transform -1 0 5850 0 1 5990
box -12 -8 474 272
use DFFSR  _3271_
timestamp 1701862152
transform -1 0 6030 0 -1 4950
box -12 -8 474 272
use DFFSR  _3272_
timestamp 1701862152
transform 1 0 4190 0 -1 4950
box -12 -8 474 272
use DFFSR  _3273_
timestamp 1701862152
transform -1 0 7910 0 -1 4950
box -12 -8 474 272
use DFFSR  _3274_
timestamp 1701862152
transform -1 0 4190 0 -1 4950
box -12 -8 474 272
use DFFSR  _3275_
timestamp 1701862152
transform -1 0 10490 0 1 7030
box -12 -8 474 272
use DFFSR  _3276_
timestamp 1701862152
transform -1 0 11270 0 1 7550
box -12 -8 474 272
use DFFSR  _3277_
timestamp 1701862152
transform -1 0 10950 0 1 7030
box -12 -8 474 272
use DFFSR  _3278_
timestamp 1701862152
transform -1 0 9850 0 1 8070
box -12 -8 474 272
use DFFSR  _3279_
timestamp 1701862152
transform -1 0 11270 0 -1 5470
box -12 -8 474 272
use DFFSR  _3280_
timestamp 1701862152
transform -1 0 10610 0 -1 8070
box -12 -8 474 272
use DFFSR  _3281_
timestamp 1701862152
transform -1 0 10410 0 -1 6510
box -12 -8 474 272
use DFFSR  _3282_
timestamp 1701862152
transform 1 0 9010 0 -1 5990
box -12 -8 474 272
use DFFSR  _3283_
timestamp 1701862152
transform -1 0 10670 0 1 6510
box -12 -8 474 272
use DFFSR  _3284_
timestamp 1701862152
transform 1 0 9810 0 -1 7550
box -12 -8 474 272
use DFFSR  _3285_
timestamp 1701862152
transform 1 0 9810 0 -1 7030
box -12 -8 474 272
use DFFSR  _3286_
timestamp 1701862152
transform 1 0 7730 0 -1 7550
box -12 -8 474 272
use DFFSR  _3287_
timestamp 1701862152
transform -1 0 10810 0 1 5470
box -12 -8 474 272
use DFFSR  _3288_
timestamp 1701862152
transform -1 0 9650 0 1 7550
box -12 -8 474 272
use DFFSR  _3289_
timestamp 1701862152
transform -1 0 10150 0 -1 5990
box -12 -8 474 272
use DFFSR  _3290_
timestamp 1701862152
transform -1 0 9470 0 1 5990
box -12 -8 474 272
use DFFSR  _3291_
timestamp 1701862152
transform 1 0 8430 0 1 7030
box -12 -8 474 272
use DFFSR  _3292_
timestamp 1701862152
transform -1 0 11290 0 1 8590
box -12 -8 474 272
use DFFSR  _3293_
timestamp 1701862152
transform 1 0 9690 0 1 8590
box -12 -8 474 272
use DFFSR  _3294_
timestamp 1701862152
transform -1 0 9590 0 1 7030
box -12 -8 474 272
use DFFSR  _3295_
timestamp 1701862152
transform -1 0 11270 0 1 5470
box -12 -8 474 272
use DFFSR  _3296_
timestamp 1701862152
transform 1 0 7510 0 1 8070
box -12 -8 474 272
use DFFSR  _3297_
timestamp 1701862152
transform -1 0 10810 0 -1 5470
box -12 -8 474 272
use DFFSR  _3298_
timestamp 1701862152
transform -1 0 9230 0 1 5470
box -12 -8 474 272
use DFFSR  _3299_
timestamp 1701862152
transform 1 0 7270 0 1 6510
box -12 -8 474 272
use DFFSR  _3300_
timestamp 1701862152
transform -1 0 8630 0 1 6510
box -12 -8 474 272
use DFFSR  _3301_
timestamp 1701862152
transform -1 0 11270 0 1 8070
box -12 -8 474 272
use DFFSR  _3302_
timestamp 1701862152
transform -1 0 10930 0 -1 8590
box -12 -8 474 272
use DFFSR  _3303_
timestamp 1701862152
transform 1 0 7870 0 -1 8070
box -12 -8 474 272
use DFFSR  _3304_
timestamp 1701862152
transform 1 0 10650 0 -1 6510
box -12 -8 474 272
use DFFSR  _3305_
timestamp 1701862152
transform -1 0 9390 0 1 8070
box -12 -8 474 272
use DFFSR  _3306_
timestamp 1701862152
transform 1 0 9450 0 -1 5470
box -12 -8 474 272
use DFFSR  _3307_
timestamp 1701862152
transform 1 0 7650 0 -1 6510
box -12 -8 474 272
use DFFSR  _3308_
timestamp 1701862152
transform -1 0 4510 0 1 6510
box -12 -8 474 272
use DFFSR  _3309_
timestamp 1701862152
transform -1 0 4810 0 1 7030
box -12 -8 474 272
use DFFSR  _3310_
timestamp 1701862152
transform 1 0 3370 0 1 7550
box -12 -8 474 272
use DFFSR  _3311_
timestamp 1701862152
transform 1 0 4330 0 -1 10150
box -12 -8 474 272
use DFFSR  _3312_
timestamp 1701862152
transform -1 0 4110 0 1 10670
box -12 -8 474 272
use DFFSR  _3313_
timestamp 1701862152
transform -1 0 4570 0 1 10670
box -12 -8 474 272
use DFFSR  _3314_
timestamp 1701862152
transform 1 0 3650 0 1 10150
box -12 -8 474 272
use DFFSR  _3315_
timestamp 1701862152
transform -1 0 5210 0 1 10150
box -12 -8 474 272
use DFFSR  _3316_
timestamp 1701862152
transform 1 0 2110 0 1 5990
box -12 -8 474 272
use DFFSR  _3317_
timestamp 1701862152
transform 1 0 2250 0 1 7030
box -12 -8 474 272
use DFFSR  _3318_
timestamp 1701862152
transform 1 0 1110 0 -1 6510
box -12 -8 474 272
use DFFSR  _3319_
timestamp 1701862152
transform 1 0 470 0 -1 8070
box -12 -8 474 272
use DFFSR  _3320_
timestamp 1701862152
transform 1 0 930 0 -1 8070
box -12 -8 474 272
use DFFSR  _3321_
timestamp 1701862152
transform 1 0 430 0 1 8590
box -12 -8 474 272
use DFFSR  _3322_
timestamp 1701862152
transform 1 0 2930 0 -1 9110
box -12 -8 474 272
use DFFSR  _3323_
timestamp 1701862152
transform 1 0 1290 0 1 8590
box -12 -8 474 272
use OR2X2  _3324_
timestamp 1702508443
transform 1 0 5690 0 1 8070
box -12 -8 92 272
use NOR2X1  _3325_
timestamp 1701862152
transform -1 0 6450 0 1 8070
box -12 -8 74 272
use NOR2X1  _3326_
timestamp 1701862152
transform -1 0 6350 0 -1 8070
box -12 -8 74 272
use NOR2X1  _3327_
timestamp 1701862152
transform -1 0 6290 0 -1 8590
box -12 -8 74 272
use NAND3X1  _3328_
timestamp 1702508443
transform -1 0 6230 0 1 8070
box -12 -8 92 272
use NOR2X1  _3329_
timestamp 1701862152
transform 1 0 5930 0 1 8070
box -12 -8 74 272
use XOR2X1  _3330_
timestamp 1702508443
transform -1 0 7210 0 1 8590
box -12 -8 132 272
use XNOR2X1  _3331_
timestamp 1702508443
transform 1 0 7390 0 -1 8590
box -12 -8 132 272
use XNOR2X1  _3332_
timestamp 1702508443
transform 1 0 7110 0 -1 8590
box -12 -8 132 272
use INVX4  _3333_
timestamp 1701862152
transform 1 0 10310 0 1 8590
box -12 -8 72 272
use INVX4  _3334_
timestamp 1701862152
transform 1 0 9410 0 1 8590
box -12 -8 72 272
use NAND2X1  _3335_
timestamp 1702508443
transform 1 0 7970 0 -1 10150
box -12 -8 72 272
use INVX2  _3336_
timestamp 1701862152
transform -1 0 6830 0 1 9630
box -12 -8 52 272
use NAND2X1  _3337_
timestamp 1702508443
transform -1 0 6370 0 1 9630
box -12 -8 72 272
use INVX2  _3338_
timestamp 1701862152
transform 1 0 7290 0 -1 10150
box -12 -8 52 272
use AND2X2  _3339_
timestamp 1701862152
transform -1 0 8230 0 1 10150
box -12 -8 94 272
use NAND2X1  _3340_
timestamp 1702508443
transform 1 0 7930 0 1 10150
box -12 -8 72 272
use AOI22X1  _3341_
timestamp 1701862152
transform 1 0 7670 0 1 10150
box -14 -8 114 272
use INVX2  _3342_
timestamp 1701862152
transform 1 0 6910 0 -1 11190
box -12 -8 52 272
use OAI21X1  _3343_
timestamp 1702508443
transform -1 0 7570 0 -1 10150
box -12 -8 92 272
use OAI21X1  _3344_
timestamp 1702508443
transform 1 0 7730 0 -1 10150
box -12 -8 92 272
use INVX4  _3345_
timestamp 1701862152
transform -1 0 9150 0 1 9630
box -12 -8 72 272
use OAI21X1  _3346_
timestamp 1702508443
transform 1 0 8630 0 1 10150
box -12 -8 92 272
use AOI21X1  _3347_
timestamp 1702508443
transform -1 0 8470 0 1 10150
box -12 -8 92 272
use NOR2X1  _3348_
timestamp 1701862152
transform 1 0 9230 0 -1 10670
box -12 -8 74 272
use AOI21X1  _3349_
timestamp 1702508443
transform 1 0 7950 0 1 9630
box -12 -8 92 272
use NAND2X1  _3350_
timestamp 1702508443
transform 1 0 7670 0 -1 8590
box -12 -8 72 272
use OAI21X1  _3351_
timestamp 1702508443
transform -1 0 7910 0 1 8590
box -12 -8 92 272
use INVX1  _3352_
timestamp 1701862152
transform -1 0 8330 0 -1 9110
box -12 -8 52 272
use OAI21X1  _3353_
timestamp 1702508443
transform 1 0 8190 0 -1 10150
box -12 -8 92 272
use NAND2X1  _3354_
timestamp 1702508443
transform 1 0 7870 0 -1 10670
box -12 -8 72 272
use AND2X2  _3355_
timestamp 1701862152
transform -1 0 7710 0 -1 10670
box -12 -8 94 272
use NAND2X1  _3356_
timestamp 1702508443
transform 1 0 7410 0 -1 10670
box -12 -8 72 272
use AOI22X1  _3357_
timestamp 1701862152
transform 1 0 7250 0 1 10670
box -14 -8 114 272
use OAI21X1  _3358_
timestamp 1702508443
transform 1 0 7510 0 1 10670
box -12 -8 92 272
use OAI21X1  _3359_
timestamp 1702508443
transform 1 0 7750 0 1 10670
box -12 -8 92 272
use NAND2X1  _3360_
timestamp 1702508443
transform -1 0 8050 0 1 10670
box -12 -8 72 272
use INVX2  _3361_
timestamp 1701862152
transform 1 0 9030 0 -1 10670
box -12 -8 52 272
use OAI21X1  _3362_
timestamp 1702508443
transform 1 0 8090 0 -1 10670
box -12 -8 92 272
use OAI21X1  _3363_
timestamp 1702508443
transform 1 0 8190 0 1 10670
box -12 -8 92 272
use NAND2X1  _3364_
timestamp 1702508443
transform 1 0 8050 0 -1 11190
box -12 -8 72 272
use AND2X2  _3365_
timestamp 1701862152
transform -1 0 7650 0 -1 11190
box -12 -8 94 272
use NAND2X1  _3366_
timestamp 1702508443
transform 1 0 7110 0 -1 11190
box -12 -8 72 272
use AOI22X1  _3367_
timestamp 1701862152
transform 1 0 6990 0 1 10670
box -14 -8 114 272
use OAI21X1  _3368_
timestamp 1702508443
transform 1 0 7330 0 -1 11190
box -12 -8 92 272
use OAI21X1  _3369_
timestamp 1702508443
transform 1 0 7810 0 -1 11190
box -12 -8 92 272
use OAI21X1  _3370_
timestamp 1702508443
transform 1 0 8310 0 -1 10670
box -12 -8 92 272
use OAI21X1  _3371_
timestamp 1702508443
transform 1 0 8430 0 1 10670
box -12 -8 92 272
use NAND2X1  _3372_
timestamp 1702508443
transform 1 0 9610 0 1 10670
box -12 -8 72 272
use NAND2X1  _3373_
timestamp 1702508443
transform -1 0 6750 0 -1 11190
box -12 -8 72 272
use AND2X2  _3374_
timestamp 1701862152
transform 1 0 5810 0 1 10670
box -12 -8 94 272
use NAND2X1  _3375_
timestamp 1702508443
transform -1 0 6110 0 1 10670
box -12 -8 72 272
use AOI22X1  _3376_
timestamp 1701862152
transform -1 0 6370 0 1 10670
box -14 -8 114 272
use OAI21X1  _3377_
timestamp 1702508443
transform 1 0 6530 0 1 10670
box -12 -8 92 272
use OAI21X1  _3378_
timestamp 1702508443
transform 1 0 6450 0 -1 11190
box -12 -8 92 272
use OAI21X1  _3379_
timestamp 1702508443
transform 1 0 8790 0 -1 10670
box -12 -8 92 272
use OAI21X1  _3380_
timestamp 1702508443
transform 1 0 8910 0 1 10670
box -12 -8 92 272
use NAND2X1  _3381_
timestamp 1702508443
transform -1 0 6830 0 1 10670
box -12 -8 72 272
use AND2X2  _3382_
timestamp 1701862152
transform 1 0 6250 0 -1 10670
box -12 -8 94 272
use NAND2X1  _3383_
timestamp 1702508443
transform -1 0 6550 0 -1 10670
box -12 -8 72 272
use AOI22X1  _3384_
timestamp 1701862152
transform -1 0 7030 0 -1 10670
box -14 -8 114 272
use OAI21X1  _3385_
timestamp 1702508443
transform 1 0 6690 0 -1 10670
box -12 -8 92 272
use OAI21X1  _3386_
timestamp 1702508443
transform 1 0 7190 0 -1 10670
box -12 -8 92 272
use OAI21X1  _3387_
timestamp 1702508443
transform 1 0 8550 0 -1 10670
box -12 -8 92 272
use OAI21X1  _3388_
timestamp 1702508443
transform 1 0 8670 0 1 10670
box -12 -8 92 272
use NAND2X1  _3389_
timestamp 1702508443
transform 1 0 10330 0 -1 10670
box -12 -8 72 272
use INVX1  _3390_
timestamp 1701862152
transform 1 0 9890 0 -1 10670
box -12 -8 52 272
use AND2X2  _3391_
timestamp 1701862152
transform 1 0 10090 0 -1 10670
box -12 -8 94 272
use OAI21X1  _3392_
timestamp 1702508443
transform 1 0 10530 0 -1 10670
box -12 -8 92 272
use INVX1  _3393_
timestamp 1701862152
transform -1 0 11310 0 -1 10150
box -12 -8 52 272
use NAND2X1  _3394_
timestamp 1702508443
transform 1 0 7470 0 1 10150
box -12 -8 72 272
use NAND3X1  _3395_
timestamp 1702508443
transform 1 0 6530 0 1 10150
box -12 -8 92 272
use AOI22X1  _3396_
timestamp 1701862152
transform -1 0 6870 0 1 10150
box -14 -8 114 272
use INVX1  _3397_
timestamp 1701862152
transform -1 0 7130 0 -1 10150
box -12 -8 52 272
use INVX1  _3398_
timestamp 1701862152
transform 1 0 6390 0 -1 10150
box -12 -8 52 272
use OAI21X1  _3399_
timestamp 1702508443
transform -1 0 6930 0 -1 10150
box -12 -8 92 272
use NAND2X1  _3400_
timestamp 1702508443
transform -1 0 7070 0 1 10150
box -12 -8 72 272
use OAI21X1  _3401_
timestamp 1702508443
transform 1 0 7230 0 1 10150
box -12 -8 92 272
use NOR2X1  _3402_
timestamp 1701862152
transform -1 0 9210 0 1 10150
box -12 -8 74 272
use XOR2X1  _3403_
timestamp 1702508443
transform 1 0 9610 0 1 10150
box -12 -8 132 272
use NAND3X1  _3404_
timestamp 1702508443
transform -1 0 5930 0 1 9630
box -12 -8 92 272
use AOI22X1  _3405_
timestamp 1701862152
transform -1 0 6230 0 -1 10150
box -14 -8 114 272
use INVX1  _3406_
timestamp 1701862152
transform 1 0 6510 0 -1 9630
box -12 -8 52 272
use NOR2X1  _3407_
timestamp 1701862152
transform -1 0 6750 0 -1 9630
box -12 -8 74 272
use OAI21X1  _3408_
timestamp 1702508443
transform 1 0 6990 0 1 9630
box -12 -8 92 272
use OAI22X1  _3409_
timestamp 1701862152
transform -1 0 6690 0 -1 10150
box -12 -8 112 272
use OAI21X1  _3410_
timestamp 1702508443
transform 1 0 9350 0 -1 10150
box -12 -8 92 272
use AOI21X1  _3411_
timestamp 1702508443
transform 1 0 9370 0 1 10150
box -12 -8 92 272
use OAI21X1  _3412_
timestamp 1702508443
transform 1 0 10090 0 1 10150
box -12 -8 92 272
use NAND2X1  _3413_
timestamp 1702508443
transform -1 0 6150 0 1 9630
box -12 -8 72 272
use NAND2X1  _3414_
timestamp 1702508443
transform 1 0 8230 0 1 9110
box -12 -8 72 272
use AOI22X1  _3415_
timestamp 1701862152
transform 1 0 6530 0 1 9630
box -14 -8 114 272
use INVX1  _3416_
timestamp 1701862152
transform 1 0 7370 0 1 8590
box -12 -8 52 272
use INVX1  _3417_
timestamp 1701862152
transform 1 0 7450 0 -1 9110
box -12 -8 52 272
use OAI21X1  _3418_
timestamp 1702508443
transform -1 0 7650 0 -1 9630
box -12 -8 92 272
use NAND2X1  _3419_
timestamp 1702508443
transform 1 0 7350 0 -1 9630
box -12 -8 72 272
use NAND2X1  _3420_
timestamp 1702508443
transform -1 0 6970 0 -1 9630
box -12 -8 72 272
use OAI21X1  _3421_
timestamp 1702508443
transform -1 0 7190 0 -1 9630
box -12 -8 92 272
use OAI21X1  _3422_
timestamp 1702508443
transform -1 0 7310 0 1 9630
box -12 -8 92 272
use INVX1  _3423_
timestamp 1701862152
transform -1 0 8330 0 -1 9630
box -12 -8 52 272
use OAI21X1  _3424_
timestamp 1702508443
transform -1 0 7890 0 -1 9630
box -12 -8 92 272
use OAI21X1  _3425_
timestamp 1702508443
transform -1 0 7550 0 1 9630
box -12 -8 92 272
use OAI21X1  _3426_
timestamp 1702508443
transform -1 0 9190 0 -1 10150
box -12 -8 92 272
use NOR2X1  _3427_
timestamp 1701862152
transform 1 0 8890 0 -1 10150
box -12 -8 74 272
use MUX2X1  _3428_
timestamp 1701862152
transform 1 0 7570 0 1 8590
box -12 -8 114 272
use NAND2X1  _3429_
timestamp 1702508443
transform 1 0 7630 0 -1 9110
box -12 -8 72 272
use NAND2X1  _3430_
timestamp 1702508443
transform -1 0 7910 0 -1 9110
box -12 -8 72 272
use AOI21X1  _3431_
timestamp 1702508443
transform 1 0 7790 0 1 9110
box -12 -8 92 272
use NAND2X1  _3432_
timestamp 1702508443
transform 1 0 8030 0 1 9110
box -12 -8 72 272
use NAND3X1  _3433_
timestamp 1702508443
transform -1 0 8130 0 -1 9630
box -12 -8 92 272
use AOI22X1  _3434_
timestamp 1701862152
transform 1 0 7710 0 1 9630
box -14 -8 114 272
use NOR2X1  _3435_
timestamp 1701862152
transform 1 0 10330 0 1 10150
box -12 -8 74 272
use OAI21X1  _3436_
timestamp 1702508443
transform -1 0 10370 0 -1 10150
box -12 -8 92 272
use NAND2X1  _3437_
timestamp 1702508443
transform 1 0 10770 0 1 10150
box -12 -8 72 272
use NAND2X1  _3438_
timestamp 1702508443
transform 1 0 10550 0 1 10150
box -12 -8 72 272
use INVX1  _3439_
timestamp 1701862152
transform 1 0 10990 0 1 10150
box -12 -8 52 272
use OAI21X1  _3440_
timestamp 1702508443
transform -1 0 10870 0 -1 10150
box -12 -8 92 272
use INVX1  _3441_
timestamp 1701862152
transform -1 0 10690 0 1 9630
box -12 -8 52 272
use AOI22X1  _3442_
timestamp 1701862152
transform -1 0 10630 0 -1 10150
box -14 -8 114 272
use XOR2X1  _3443_
timestamp 1702508443
transform -1 0 11190 0 1 9630
box -12 -8 132 272
use AOI21X1  _3444_
timestamp 1702508443
transform -1 0 8570 0 -1 9630
box -12 -8 92 272
use OAI21X1  _3445_
timestamp 1702508443
transform -1 0 8270 0 1 9630
box -12 -8 92 272
use INVX1  _3446_
timestamp 1701862152
transform 1 0 8650 0 1 9630
box -12 -8 52 272
use NOR2X1  _3447_
timestamp 1701862152
transform 1 0 8430 0 1 9630
box -12 -8 74 272
use OAI21X1  _3448_
timestamp 1702508443
transform -1 0 8930 0 1 9630
box -12 -8 92 272
use INVX1  _3449_
timestamp 1701862152
transform -1 0 9930 0 1 10150
box -12 -8 52 272
use OAI21X1  _3450_
timestamp 1702508443
transform -1 0 9910 0 -1 10150
box -12 -8 92 272
use MUX2X1  _3451_
timestamp 1701862152
transform 1 0 9590 0 -1 10150
box -12 -8 114 272
use NAND2X1  _3452_
timestamp 1702508443
transform -1 0 9370 0 1 9630
box -12 -8 72 272
use OAI21X1  _3453_
timestamp 1702508443
transform -1 0 10150 0 -1 10150
box -12 -8 92 272
use NAND2X1  _3454_
timestamp 1702508443
transform 1 0 9530 0 1 9630
box -12 -8 72 272
use NAND2X1  _3455_
timestamp 1702508443
transform 1 0 9750 0 1 9630
box -12 -8 72 272
use NAND2X1  _3456_
timestamp 1702508443
transform -1 0 10490 0 1 9630
box -12 -8 72 272
use NAND3X1  _3457_
timestamp 1702508443
transform -1 0 10050 0 1 9630
box -12 -8 92 272
use NAND3X1  _3458_
timestamp 1702508443
transform -1 0 10270 0 1 9630
box -12 -8 92 272
use NAND2X1  _3459_
timestamp 1702508443
transform -1 0 10410 0 -1 9630
box -12 -8 72 272
use OAI21X1  _3460_
timestamp 1702508443
transform 1 0 11030 0 -1 10150
box -12 -8 92 272
use INVX1  _3461_
timestamp 1701862152
transform -1 0 11290 0 -1 9630
box -12 -8 52 272
use OAI21X1  _3462_
timestamp 1702508443
transform -1 0 10870 0 -1 9630
box -12 -8 92 272
use NAND2X1  _3463_
timestamp 1702508443
transform 1 0 10490 0 -1 11190
box -12 -8 72 272
use OAI21X1  _3464_
timestamp 1702508443
transform 1 0 9830 0 -1 11190
box -12 -8 92 272
use INVX1  _3465_
timestamp 1701862152
transform 1 0 10050 0 -1 11190
box -12 -8 52 272
use OAI21X1  _3466_
timestamp 1702508443
transform 1 0 10250 0 -1 11190
box -12 -8 92 272
use INVX1  _3467_
timestamp 1701862152
transform -1 0 11250 0 1 10670
box -12 -8 52 272
use AOI22X1  _3468_
timestamp 1701862152
transform 1 0 10730 0 1 10670
box -14 -8 114 272
use OAI21X1  _3469_
timestamp 1702508443
transform 1 0 9450 0 -1 10670
box -12 -8 92 272
use INVX1  _3470_
timestamp 1701862152
transform 1 0 9690 0 -1 10670
box -12 -8 52 272
use OAI21X1  _3471_
timestamp 1702508443
transform 1 0 9830 0 1 10670
box -12 -8 92 272
use OAI21X1  _3472_
timestamp 1702508443
transform -1 0 10130 0 1 10670
box -12 -8 92 272
use NAND2X1  _3473_
timestamp 1702508443
transform 1 0 8710 0 -1 11190
box -12 -8 72 272
use OAI21X1  _3474_
timestamp 1702508443
transform 1 0 8270 0 -1 11190
box -12 -8 92 272
use INVX1  _3475_
timestamp 1701862152
transform 1 0 8510 0 -1 11190
box -12 -8 52 272
use OAI21X1  _3476_
timestamp 1702508443
transform -1 0 9010 0 -1 11190
box -12 -8 92 272
use INVX1  _3477_
timestamp 1701862152
transform 1 0 9170 0 -1 11190
box -12 -8 52 272
use AOI22X1  _3478_
timestamp 1701862152
transform 1 0 9150 0 1 10670
box -14 -8 114 272
use OAI21X1  _3479_
timestamp 1702508443
transform 1 0 8430 0 -1 10150
box -12 -8 92 272
use OAI21X1  _3480_
timestamp 1702508443
transform -1 0 8730 0 -1 10150
box -12 -8 92 272
use NAND2X1  _3481_
timestamp 1702508443
transform -1 0 8510 0 1 9110
box -12 -8 72 272
use XOR2X1  _3482_
timestamp 1702508443
transform -1 0 8790 0 1 9110
box -12 -8 132 272
use XOR2X1  _3483_
timestamp 1702508443
transform 1 0 8870 0 1 10150
box -12 -8 132 272
use INVX1  _3484_
timestamp 1701862152
transform -1 0 10190 0 -1 9630
box -12 -8 52 272
use XOR2X1  _3485_
timestamp 1702508443
transform 1 0 11190 0 1 10150
box -12 -8 132 272
use XOR2X1  _3486_
timestamp 1702508443
transform 1 0 10530 0 1 9110
box -12 -8 132 272
use AOI21X1  _3487_
timestamp 1702508443
transform 1 0 10550 0 -1 9630
box -12 -8 92 272
use AOI21X1  _3488_
timestamp 1702508443
transform -1 0 10930 0 1 9630
box -12 -8 92 272
use OAI21X1  _3489_
timestamp 1702508443
transform 1 0 10710 0 -1 11190
box -12 -8 92 272
use INVX1  _3490_
timestamp 1701862152
transform 1 0 11170 0 -1 11190
box -12 -8 52 272
use NAND2X1  _3491_
timestamp 1702508443
transform -1 0 11010 0 -1 11190
box -12 -8 72 272
use NAND2X1  _3492_
timestamp 1702508443
transform -1 0 10570 0 1 10670
box -12 -8 72 272
use NAND2X1  _3493_
timestamp 1702508443
transform -1 0 10350 0 1 10670
box -12 -8 72 272
use NAND2X1  _3494_
timestamp 1702508443
transform 1 0 9390 0 1 10670
box -12 -8 72 272
use NAND3X1  _3495_
timestamp 1702508443
transform -1 0 9670 0 -1 11190
box -12 -8 92 272
use NAND2X1  _3496_
timestamp 1702508443
transform 1 0 9370 0 -1 11190
box -12 -8 72 272
use AOI21X1  _3497_
timestamp 1702508443
transform -1 0 9530 0 -1 9630
box -12 -8 92 272
use AOI21X1  _3498_
timestamp 1702508443
transform -1 0 9030 0 1 9110
box -12 -8 92 272
use AOI22X1  _3499_
timestamp 1701862152
transform 1 0 8490 0 -1 9110
box -14 -8 114 272
use NAND2X1  _3500_
timestamp 1702508443
transform 1 0 9870 0 1 9110
box -12 -8 72 272
use OAI21X1  _3501_
timestamp 1702508443
transform -1 0 10150 0 1 9110
box -12 -8 92 272
use NAND2X1  _3502_
timestamp 1702508443
transform -1 0 8410 0 -1 8590
box -12 -8 72 272
use AOI21X1  _3503_
timestamp 1702508443
transform -1 0 8810 0 -1 9630
box -12 -8 92 272
use OAI21X1  _3504_
timestamp 1702508443
transform 1 0 8970 0 -1 9630
box -12 -8 92 272
use OAI21X1  _3505_
timestamp 1702508443
transform -1 0 9290 0 -1 9630
box -12 -8 92 272
use OAI21X1  _3506_
timestamp 1702508443
transform -1 0 8810 0 1 8590
box -12 -8 92 272
use NAND2X1  _3507_
timestamp 1702508443
transform 1 0 10830 0 -1 9110
box -12 -8 72 272
use OAI21X1  _3508_
timestamp 1702508443
transform 1 0 10590 0 -1 9110
box -12 -8 92 272
use NAND2X1  _3509_
timestamp 1702508443
transform 1 0 8510 0 1 8590
box -12 -8 72 272
use OAI21X1  _3510_
timestamp 1702508443
transform -1 0 9050 0 1 8590
box -12 -8 92 272
use NAND2X1  _3511_
timestamp 1702508443
transform 1 0 10050 0 -1 270
box -12 -8 72 272
use OAI21X1  _3512_
timestamp 1702508443
transform 1 0 11050 0 -1 9110
box -12 -8 92 272
use NAND2X1  _3513_
timestamp 1702508443
transform 1 0 11030 0 -1 9630
box -12 -8 72 272
use NOR2X1  _3514_
timestamp 1701862152
transform 1 0 10990 0 1 10670
box -12 -8 74 272
use OAI21X1  _3515_
timestamp 1702508443
transform -1 0 10850 0 -1 10670
box -12 -8 92 272
use OAI21X1  _3516_
timestamp 1702508443
transform 1 0 10990 0 -1 10670
box -12 -8 92 272
use NAND2X1  _3517_
timestamp 1702508443
transform 1 0 9690 0 -1 9630
box -12 -8 72 272
use OAI21X1  _3518_
timestamp 1702508443
transform 1 0 9910 0 -1 9630
box -12 -8 92 272
use NAND2X1  _3519_
timestamp 1702508443
transform 1 0 9190 0 1 9110
box -12 -8 72 272
use OAI21X1  _3520_
timestamp 1702508443
transform -1 0 9490 0 1 9110
box -12 -8 92 272
use INVX1  _3521_
timestamp 1701862152
transform 1 0 6670 0 1 8590
box -12 -8 52 272
use NAND2X1  _3522_
timestamp 1702508443
transform 1 0 8070 0 -1 9110
box -12 -8 72 272
use OAI21X1  _3523_
timestamp 1702508443
transform 1 0 6850 0 1 8590
box -12 -8 92 272
use INVX1  _3524_
timestamp 1701862152
transform 1 0 7590 0 1 9110
box -12 -8 52 272
use NAND2X1  _3525_
timestamp 1702508443
transform 1 0 7130 0 1 9110
box -12 -8 72 272
use OAI21X1  _3526_
timestamp 1702508443
transform -1 0 7430 0 1 9110
box -12 -8 92 272
use DFFSR  _3527_
timestamp 1701862152
transform -1 0 8190 0 -1 8590
box -12 -8 474 272
use DFFSR  _3528_
timestamp 1701862152
transform -1 0 8370 0 1 8590
box -12 -8 474 272
use DFFSR  _3529_
timestamp 1701862152
transform -1 0 9970 0 -1 9110
box -12 -8 474 272
use DFFSR  _3530_
timestamp 1701862152
transform -1 0 8870 0 -1 8590
box -12 -8 474 272
use DFFSR  _3531_
timestamp 1701862152
transform -1 0 10430 0 -1 9110
box -12 -8 474 272
use DFFSR  _3532_
timestamp 1701862152
transform -1 0 9330 0 -1 8590
box -12 -8 474 272
use DFFSR  _3533_
timestamp 1701862152
transform -1 0 10830 0 1 8590
box -12 -8 474 272
use DFFSR  _3534_
timestamp 1701862152
transform -1 0 11110 0 1 9110
box -12 -8 474 272
use DFFSR  _3535_
timestamp 1701862152
transform -1 0 9510 0 -1 9110
box -12 -8 474 272
use DFFSR  _3536_
timestamp 1701862152
transform -1 0 9050 0 -1 9110
box -12 -8 474 272
use DFFSR  _3537_
timestamp 1701862152
transform -1 0 6950 0 -1 8590
box -12 -8 474 272
use DFFSR  _3538_
timestamp 1701862152
transform 1 0 6830 0 -1 9110
box -12 -8 474 272
use BUFX2  _3539_ ~/ETRI050_DesignKit/devel/Ref_Design/CPU_6502/layout/digital_ETRI
timestamp 1702508443
transform 1 0 11230 0 -1 7030
box -12 -8 72 272
use BUFX2  _3540_
timestamp 1702508443
transform 1 0 4730 0 1 10670
box -12 -8 72 272
use BUFX2  _3541_
timestamp 1702508443
transform -1 0 230 0 1 5990
box -12 -8 72 272
use BUFX2  _3542_
timestamp 1702508443
transform -1 0 230 0 -1 8070
box -12 -8 72 272
use BUFX2  _3543_
timestamp 1702508443
transform -1 0 210 0 1 8590
box -12 -8 72 272
use BUFX2  _3544_
timestamp 1702508443
transform -1 0 230 0 1 9110
box -12 -8 72 272
use BUFX2  _3545_
timestamp 1702508443
transform -1 0 2070 0 -1 11190
box -12 -8 72 272
use BUFX2  _3546_
timestamp 1702508443
transform -1 0 690 0 1 9110
box -12 -8 72 272
use BUFX2  _3547_
timestamp 1702508443
transform 1 0 4770 0 -1 11190
box -12 -8 72 272
use BUFX2  _3548_
timestamp 1702508443
transform 1 0 5370 0 1 10670
box -12 -8 72 272
use BUFX2  _3549_
timestamp 1702508443
transform -1 0 4410 0 -1 11190
box -12 -8 72 272
use BUFX2  _3550_
timestamp 1702508443
transform -1 0 5230 0 -1 11190
box -12 -8 72 272
use BUFX2  _3551_
timestamp 1702508443
transform 1 0 5610 0 -1 11190
box -12 -8 72 272
use BUFX2  _3552_
timestamp 1702508443
transform 1 0 5390 0 -1 11190
box -12 -8 72 272
use BUFX2  _3553_
timestamp 1702508443
transform -1 0 230 0 -1 5990
box -12 -8 72 272
use BUFX2  _3554_
timestamp 1702508443
transform -1 0 430 0 1 7030
box -12 -8 72 272
use BUFX2  _3555_
timestamp 1702508443
transform -1 0 5210 0 1 10670
box -12 -8 72 272
use BUFX2  _3556_
timestamp 1702508443
transform 1 0 6310 0 1 10150
box -12 -8 72 272
use BUFX2  _3557_
timestamp 1702508443
transform -1 0 5870 0 -1 11190
box -12 -8 72 272
use BUFX2  _3558_
timestamp 1702508443
transform 1 0 6250 0 -1 11190
box -12 -8 72 272
use BUFX2  _3559_
timestamp 1702508443
transform -1 0 4950 0 -1 10670
box -12 -8 72 272
use BUFX2  _3560_
timestamp 1702508443
transform 1 0 5590 0 1 10670
box -12 -8 72 272
use BUFX2  _3561_
timestamp 1702508443
transform 1 0 6030 0 -1 11190
box -12 -8 72 272
use BUFX2  _3562_
timestamp 1702508443
transform 1 0 5830 0 1 10150
box -12 -8 72 272
use BUFX2  _3563_
timestamp 1702508443
transform 1 0 5290 0 1 3390
box -12 -8 72 272
use BUFX2  BUFX2_insert0
timestamp 1702508443
transform 1 0 5910 0 -1 10150
box -12 -8 72 272
use BUFX2  BUFX2_insert1
timestamp 1702508443
transform 1 0 6670 0 1 2350
box -12 -8 72 272
use BUFX2  BUFX2_insert2
timestamp 1702508443
transform 1 0 5510 0 -1 1830
box -12 -8 72 272
use BUFX2  BUFX2_insert3
timestamp 1702508443
transform -1 0 690 0 -1 5470
box -12 -8 72 272
use BUFX2  BUFX2_insert4
timestamp 1702508443
transform 1 0 3390 0 1 4950
box -12 -8 72 272
use BUFX2  BUFX2_insert5
timestamp 1702508443
transform 1 0 1450 0 -1 1830
box -12 -8 72 272
use BUFX2  BUFX2_insert6
timestamp 1702508443
transform -1 0 210 0 -1 11190
box -12 -8 72 272
use BUFX2  BUFX2_insert7
timestamp 1702508443
transform 1 0 1750 0 1 10670
box -12 -8 72 272
use BUFX2  BUFX2_insert8
timestamp 1702508443
transform 1 0 1710 0 1 1830
box -12 -8 72 272
use BUFX2  BUFX2_insert9
timestamp 1702508443
transform 1 0 2010 0 -1 3910
box -12 -8 72 272
use BUFX2  BUFX2_insert10
timestamp 1702508443
transform 1 0 1830 0 -1 4430
box -12 -8 72 272
use BUFX2  BUFX2_insert11
timestamp 1702508443
transform -1 0 1850 0 -1 3910
box -12 -8 72 272
use BUFX2  BUFX2_insert12
timestamp 1702508443
transform -1 0 1630 0 -1 3910
box -12 -8 72 272
use BUFX2  BUFX2_insert13
timestamp 1702508443
transform -1 0 1530 0 -1 1310
box -12 -8 72 272
use BUFX2  BUFX2_insert14
timestamp 1702508443
transform -1 0 3750 0 1 3390
box -12 -8 72 272
use BUFX2  BUFX2_insert15
timestamp 1702508443
transform 1 0 4610 0 -1 5470
box -12 -8 72 272
use BUFX2  BUFX2_insert16
timestamp 1702508443
transform 1 0 1410 0 -1 4950
box -12 -8 72 272
use BUFX2  BUFX2_insert17
timestamp 1702508443
transform 1 0 3690 0 1 1310
box -12 -8 72 272
use BUFX2  BUFX2_insert18
timestamp 1702508443
transform -1 0 9870 0 1 2350
box -12 -8 72 272
use BUFX2  BUFX2_insert19
timestamp 1702508443
transform -1 0 8610 0 -1 790
box -12 -8 72 272
use BUFX2  BUFX2_insert20
timestamp 1702508443
transform 1 0 10030 0 1 2350
box -12 -8 72 272
use BUFX2  BUFX2_insert21
timestamp 1702508443
transform -1 0 7890 0 -1 1310
box -12 -8 72 272
use BUFX2  BUFX2_insert22
timestamp 1702508443
transform -1 0 3310 0 -1 2870
box -12 -8 72 272
use BUFX2  BUFX2_insert23
timestamp 1702508443
transform -1 0 2850 0 -1 4950
box -12 -8 72 272
use BUFX2  BUFX2_insert24
timestamp 1702508443
transform -1 0 3750 0 -1 4430
box -12 -8 72 272
use BUFX2  BUFX2_insert25
timestamp 1702508443
transform 1 0 4450 0 1 4430
box -12 -8 72 272
use BUFX2  BUFX2_insert26
timestamp 1702508443
transform 1 0 4270 0 1 2870
box -12 -8 72 272
use BUFX2  BUFX2_insert27
timestamp 1702508443
transform 1 0 9670 0 1 4950
box -12 -8 72 272
use BUFX2  BUFX2_insert28
timestamp 1702508443
transform -1 0 7570 0 -1 5990
box -12 -8 72 272
use BUFX2  BUFX2_insert29
timestamp 1702508443
transform -1 0 1390 0 1 6510
box -12 -8 72 272
use BUFX2  BUFX2_insert30
timestamp 1702508443
transform -1 0 8890 0 -1 3910
box -12 -8 72 272
use BUFX2  BUFX2_insert31
timestamp 1702508443
transform -1 0 9670 0 1 3910
box -12 -8 72 272
use BUFX2  BUFX2_insert32
timestamp 1702508443
transform 1 0 5930 0 -1 3910
box -12 -8 72 272
use BUFX2  BUFX2_insert33
timestamp 1702508443
transform -1 0 9650 0 -1 4950
box -12 -8 72 272
use BUFX2  BUFX2_insert34
timestamp 1702508443
transform 1 0 5270 0 1 8590
box -12 -8 72 272
use BUFX2  BUFX2_insert35
timestamp 1702508443
transform -1 0 6070 0 1 7550
box -12 -8 72 272
use BUFX2  BUFX2_insert36
timestamp 1702508443
transform -1 0 1290 0 1 8590
box -12 -8 72 272
use BUFX2  BUFX2_insert37
timestamp 1702508443
transform -1 0 9690 0 1 8590
box -12 -8 72 272
use BUFX2  BUFX2_insert49
timestamp 1702508443
transform -1 0 3150 0 1 6510
box -12 -8 72 272
use BUFX2  BUFX2_insert50
timestamp 1702508443
transform 1 0 2390 0 -1 8590
box -12 -8 72 272
use BUFX2  BUFX2_insert51
timestamp 1702508443
transform 1 0 3270 0 -1 8590
box -12 -8 72 272
use BUFX2  BUFX2_insert52
timestamp 1702508443
transform 1 0 3450 0 1 5470
box -12 -8 72 272
use BUFX2  BUFX2_insert53
timestamp 1702508443
transform -1 0 11330 0 1 9110
box -12 -8 72 272
use BUFX2  BUFX2_insert54
timestamp 1702508443
transform -1 0 9270 0 1 8590
box -12 -8 72 272
use BUFX2  BUFX2_insert55
timestamp 1702508443
transform -1 0 9710 0 1 9110
box -12 -8 72 272
use BUFX2  BUFX2_insert56
timestamp 1702508443
transform -1 0 10370 0 1 9110
box -12 -8 72 272
use BUFX2  BUFX2_insert57
timestamp 1702508443
transform -1 0 11310 0 -1 2350
box -12 -8 72 272
use BUFX2  BUFX2_insert58
timestamp 1702508443
transform -1 0 9070 0 1 2870
box -12 -8 72 272
use BUFX2  BUFX2_insert59
timestamp 1702508443
transform -1 0 7650 0 1 1830
box -12 -8 72 272
use BUFX2  BUFX2_insert60
timestamp 1702508443
transform 1 0 10950 0 1 1830
box -12 -8 72 272
use BUFX2  BUFX2_insert61
timestamp 1702508443
transform -1 0 11270 0 1 2870
box -12 -8 72 272
use BUFX2  BUFX2_insert62
timestamp 1702508443
transform 1 0 2270 0 1 3910
box -12 -8 72 272
use BUFX2  BUFX2_insert63
timestamp 1702508443
transform 1 0 2190 0 1 3390
box -12 -8 72 272
use BUFX2  BUFX2_insert64
timestamp 1702508443
transform -1 0 1890 0 1 3910
box -12 -8 72 272
use BUFX2  BUFX2_insert65
timestamp 1702508443
transform -1 0 1810 0 1 3390
box -12 -8 72 272
use BUFX2  BUFX2_insert66
timestamp 1702508443
transform -1 0 4410 0 1 1310
box -12 -8 72 272
use BUFX2  BUFX2_insert67
timestamp 1702508443
transform -1 0 3710 0 -1 10150
box -12 -8 72 272
use BUFX2  BUFX2_insert68
timestamp 1702508443
transform -1 0 7270 0 1 2870
box -12 -8 72 272
use BUFX2  BUFX2_insert69
timestamp 1702508443
transform -1 0 5750 0 -1 3390
box -12 -8 72 272
use BUFX2  BUFX2_insert70
timestamp 1702508443
transform -1 0 3770 0 -1 1830
box -12 -8 72 272
use BUFX2  BUFX2_insert71
timestamp 1702508443
transform -1 0 7410 0 1 2350
box -12 -8 72 272
use BUFX2  BUFX2_insert72
timestamp 1702508443
transform -1 0 6570 0 1 1310
box -12 -8 72 272
use BUFX2  BUFX2_insert73
timestamp 1702508443
transform 1 0 3670 0 1 5470
box -12 -8 72 272
use BUFX2  BUFX2_insert74
timestamp 1702508443
transform 1 0 7630 0 -1 2350
box -12 -8 72 272
use BUFX2  BUFX2_insert75
timestamp 1702508443
transform 1 0 7650 0 1 2870
box -12 -8 72 272
use BUFX2  BUFX2_insert76
timestamp 1702508443
transform 1 0 7430 0 1 2870
box -12 -8 72 272
use BUFX2  BUFX2_insert77
timestamp 1702508443
transform -1 0 3530 0 -1 2870
box -12 -8 72 272
use BUFX2  BUFX2_insert78
timestamp 1702508443
transform 1 0 1990 0 -1 2870
box -12 -8 72 272
use BUFX2  BUFX2_insert79
timestamp 1702508443
transform -1 0 2250 0 -1 2870
box -12 -8 72 272
use BUFX2  BUFX2_insert80
timestamp 1702508443
transform 1 0 2470 0 1 4430
box -12 -8 72 272
use BUFX2  BUFX2_insert81
timestamp 1702508443
transform -1 0 2110 0 1 3910
box -12 -8 72 272
use BUFX2  BUFX2_insert82
timestamp 1702508443
transform -1 0 430 0 1 8590
box -12 -8 72 272
use BUFX2  BUFX2_insert83
timestamp 1702508443
transform 1 0 4270 0 -1 10150
box -12 -8 72 272
use BUFX2  BUFX2_insert84
timestamp 1702508443
transform 1 0 4230 0 -1 7550
box -12 -8 72 272
use BUFX2  BUFX2_insert85
timestamp 1702508443
transform -1 0 230 0 -1 6510
box -12 -8 72 272
use BUFX2  BUFX2_insert86
timestamp 1702508443
transform 1 0 1990 0 -1 10150
box -12 -8 72 272
use CLKBUF1  CLKBUF1_insert38 ~/ETRI050_DesignKit/devel/Ref_Design/CPU_6502/layout/digital_ETRI
timestamp 1701862152
transform 1 0 2990 0 -1 7550
box -12 -8 192 272
use CLKBUF1  CLKBUF1_insert39
timestamp 1701862152
transform -1 0 4950 0 -1 6510
box -12 -8 192 272
use CLKBUF1  CLKBUF1_insert40
timestamp 1701862152
transform -1 0 1250 0 -1 4950
box -12 -8 192 272
use CLKBUF1  CLKBUF1_insert41
timestamp 1701862152
transform -1 0 10910 0 -1 270
box -12 -8 192 272
use CLKBUF1  CLKBUF1_insert42
timestamp 1701862152
transform 1 0 9810 0 -1 4950
box -12 -8 192 272
use CLKBUF1  CLKBUF1_insert43
timestamp 1701862152
transform -1 0 11270 0 1 7030
box -12 -8 192 272
use CLKBUF1  CLKBUF1_insert44
timestamp 1701862152
transform -1 0 11030 0 1 4430
box -12 -8 192 272
use CLKBUF1  CLKBUF1_insert45
timestamp 1701862152
transform 1 0 5790 0 -1 6510
box -12 -8 192 272
use CLKBUF1  CLKBUF1_insert46
timestamp 1701862152
transform 1 0 4110 0 1 5990
box -12 -8 192 272
use CLKBUF1  CLKBUF1_insert47
timestamp 1701862152
transform -1 0 2390 0 1 7550
box -12 -8 192 272
use CLKBUF1  CLKBUF1_insert48
timestamp 1701862152
transform -1 0 11070 0 -1 7030
box -12 -8 192 272
use FILL  FILL166650x93750 ~/ETRI050_DesignKit/devel/Ref_Design/CPU_6502/layout/digital_ETRI
timestamp 1701859473
transform -1 0 11130 0 -1 6510
box -12 -8 32 272
use FILL  FILL166950x4050
timestamp 1701859473
transform 1 0 11130 0 1 270
box -12 -8 32 272
use FILL  FILL166950x54750
timestamp 1701859473
transform -1 0 11150 0 -1 3910
box -12 -8 32 272
use FILL  FILL166950x70350
timestamp 1701859473
transform -1 0 11150 0 -1 4950
box -12 -8 32 272
use FILL  FILL166950x93750
timestamp 1701859473
transform -1 0 11150 0 -1 6510
box -12 -8 32 272
use FILL  FILL166950x132750
timestamp 1701859473
transform -1 0 11150 0 -1 9110
box -12 -8 32 272
use FILL  FILL167250x150
timestamp 1701859473
transform -1 0 11170 0 -1 270
box -12 -8 32 272
use FILL  FILL167250x4050
timestamp 1701859473
transform 1 0 11150 0 1 270
box -12 -8 32 272
use FILL  FILL167250x54750
timestamp 1701859473
transform -1 0 11170 0 -1 3910
box -12 -8 32 272
use FILL  FILL167250x70350
timestamp 1701859473
transform -1 0 11170 0 -1 4950
box -12 -8 32 272
use FILL  FILL167250x93750
timestamp 1701859473
transform -1 0 11170 0 -1 6510
box -12 -8 32 272
use FILL  FILL167250x109350
timestamp 1701859473
transform -1 0 11170 0 -1 7550
box -12 -8 32 272
use FILL  FILL167250x124950
timestamp 1701859473
transform -1 0 11170 0 -1 8590
box -12 -8 32 272
use FILL  FILL167250x132750
timestamp 1701859473
transform -1 0 11170 0 -1 9110
box -12 -8 32 272
use FILL  FILL167550x150
timestamp 1701859473
transform -1 0 11190 0 -1 270
box -12 -8 32 272
use FILL  FILL167550x4050
timestamp 1701859473
transform 1 0 11170 0 1 270
box -12 -8 32 272
use FILL  FILL167550x11850
timestamp 1701859473
transform 1 0 11170 0 1 790
box -12 -8 32 272
use FILL  FILL167550x54750
timestamp 1701859473
transform -1 0 11190 0 -1 3910
box -12 -8 32 272
use FILL  FILL167550x70350
timestamp 1701859473
transform -1 0 11190 0 -1 4950
box -12 -8 32 272
use FILL  FILL167550x93750
timestamp 1701859473
transform -1 0 11190 0 -1 6510
box -12 -8 32 272
use FILL  FILL167550x109350
timestamp 1701859473
transform -1 0 11190 0 -1 7550
box -12 -8 32 272
use FILL  FILL167550x124950
timestamp 1701859473
transform -1 0 11190 0 -1 8590
box -12 -8 32 272
use FILL  FILL167550x132750
timestamp 1701859473
transform -1 0 11190 0 -1 9110
box -12 -8 32 272
use FILL  FILL167850x150
timestamp 1701859473
transform -1 0 11210 0 -1 270
box -12 -8 32 272
use FILL  FILL167850x4050
timestamp 1701859473
transform 1 0 11190 0 1 270
box -12 -8 32 272
use FILL  FILL167850x11850
timestamp 1701859473
transform 1 0 11190 0 1 790
box -12 -8 32 272
use FILL  FILL167850x54750
timestamp 1701859473
transform -1 0 11210 0 -1 3910
box -12 -8 32 272
use FILL  FILL167850x70350
timestamp 1701859473
transform -1 0 11210 0 -1 4950
box -12 -8 32 272
use FILL  FILL167850x93750
timestamp 1701859473
transform -1 0 11210 0 -1 6510
box -12 -8 32 272
use FILL  FILL167850x109350
timestamp 1701859473
transform -1 0 11210 0 -1 7550
box -12 -8 32 272
use FILL  FILL167850x124950
timestamp 1701859473
transform -1 0 11210 0 -1 8590
box -12 -8 32 272
use FILL  FILL167850x132750
timestamp 1701859473
transform -1 0 11210 0 -1 9110
box -12 -8 32 272
use FILL  FILL167850x144450
timestamp 1701859473
transform 1 0 11190 0 1 9630
box -12 -8 32 272
use FILL  FILL168150x150
timestamp 1701859473
transform -1 0 11230 0 -1 270
box -12 -8 32 272
use FILL  FILL168150x4050
timestamp 1701859473
transform 1 0 11210 0 1 270
box -12 -8 32 272
use FILL  FILL168150x11850
timestamp 1701859473
transform 1 0 11210 0 1 790
box -12 -8 32 272
use FILL  FILL168150x54750
timestamp 1701859473
transform -1 0 11230 0 -1 3910
box -12 -8 32 272
use FILL  FILL168150x58650
timestamp 1701859473
transform 1 0 11210 0 1 3910
box -12 -8 32 272
use FILL  FILL168150x70350
timestamp 1701859473
transform -1 0 11230 0 -1 4950
box -12 -8 32 272
use FILL  FILL168150x93750
timestamp 1701859473
transform -1 0 11230 0 -1 6510
box -12 -8 32 272
use FILL  FILL168150x109350
timestamp 1701859473
transform -1 0 11230 0 -1 7550
box -12 -8 32 272
use FILL  FILL168150x124950
timestamp 1701859473
transform -1 0 11230 0 -1 8590
box -12 -8 32 272
use FILL  FILL168150x132750
timestamp 1701859473
transform -1 0 11230 0 -1 9110
box -12 -8 32 272
use FILL  FILL168150x144450
timestamp 1701859473
transform 1 0 11210 0 1 9630
box -12 -8 32 272
use FILL  FILL168150x163950
timestamp 1701859473
transform -1 0 11230 0 -1 11190
box -12 -8 32 272
use FILL  FILL168450x150
timestamp 1701859473
transform -1 0 11250 0 -1 270
box -12 -8 32 272
use FILL  FILL168450x4050
timestamp 1701859473
transform 1 0 11230 0 1 270
box -12 -8 32 272
use FILL  FILL168450x11850
timestamp 1701859473
transform 1 0 11230 0 1 790
box -12 -8 32 272
use FILL  FILL168450x35250
timestamp 1701859473
transform 1 0 11230 0 1 2350
box -12 -8 32 272
use FILL  FILL168450x54750
timestamp 1701859473
transform -1 0 11250 0 -1 3910
box -12 -8 32 272
use FILL  FILL168450x58650
timestamp 1701859473
transform 1 0 11230 0 1 3910
box -12 -8 32 272
use FILL  FILL168450x66450
timestamp 1701859473
transform 1 0 11230 0 1 4430
box -12 -8 32 272
use FILL  FILL168450x70350
timestamp 1701859473
transform -1 0 11250 0 -1 4950
box -12 -8 32 272
use FILL  FILL168450x93750
timestamp 1701859473
transform -1 0 11250 0 -1 6510
box -12 -8 32 272
use FILL  FILL168450x109350
timestamp 1701859473
transform -1 0 11250 0 -1 7550
box -12 -8 32 272
use FILL  FILL168450x124950
timestamp 1701859473
transform -1 0 11250 0 -1 8590
box -12 -8 32 272
use FILL  FILL168450x132750
timestamp 1701859473
transform -1 0 11250 0 -1 9110
box -12 -8 32 272
use FILL  FILL168450x144450
timestamp 1701859473
transform 1 0 11230 0 1 9630
box -12 -8 32 272
use FILL  FILL168450x163950
timestamp 1701859473
transform -1 0 11250 0 -1 11190
box -12 -8 32 272
use FILL  FILL168750x150
timestamp 1701859473
transform -1 0 11270 0 -1 270
box -12 -8 32 272
use FILL  FILL168750x4050
timestamp 1701859473
transform 1 0 11250 0 1 270
box -12 -8 32 272
use FILL  FILL168750x11850
timestamp 1701859473
transform 1 0 11250 0 1 790
box -12 -8 32 272
use FILL  FILL168750x15750
timestamp 1701859473
transform -1 0 11270 0 -1 1310
box -12 -8 32 272
use FILL  FILL168750x27450
timestamp 1701859473
transform 1 0 11250 0 1 1830
box -12 -8 32 272
use FILL  FILL168750x35250
timestamp 1701859473
transform 1 0 11250 0 1 2350
box -12 -8 32 272
use FILL  FILL168750x46950
timestamp 1701859473
transform -1 0 11270 0 -1 3390
box -12 -8 32 272
use FILL  FILL168750x54750
timestamp 1701859473
transform -1 0 11270 0 -1 3910
box -12 -8 32 272
use FILL  FILL168750x58650
timestamp 1701859473
transform 1 0 11250 0 1 3910
box -12 -8 32 272
use FILL  FILL168750x62550
timestamp 1701859473
transform -1 0 11270 0 -1 4430
box -12 -8 32 272
use FILL  FILL168750x66450
timestamp 1701859473
transform 1 0 11250 0 1 4430
box -12 -8 32 272
use FILL  FILL168750x70350
timestamp 1701859473
transform -1 0 11270 0 -1 4950
box -12 -8 32 272
use FILL  FILL168750x93750
timestamp 1701859473
transform -1 0 11270 0 -1 6510
box -12 -8 32 272
use FILL  FILL168750x109350
timestamp 1701859473
transform -1 0 11270 0 -1 7550
box -12 -8 32 272
use FILL  FILL168750x124950
timestamp 1701859473
transform -1 0 11270 0 -1 8590
box -12 -8 32 272
use FILL  FILL168750x132750
timestamp 1701859473
transform -1 0 11270 0 -1 9110
box -12 -8 32 272
use FILL  FILL168750x144450
timestamp 1701859473
transform 1 0 11250 0 1 9630
box -12 -8 32 272
use FILL  FILL168750x160050
timestamp 1701859473
transform 1 0 11250 0 1 10670
box -12 -8 32 272
use FILL  FILL168750x163950
timestamp 1701859473
transform -1 0 11270 0 -1 11190
box -12 -8 32 272
use FILL  FILL169050x150
timestamp 1701859473
transform -1 0 11290 0 -1 270
box -12 -8 32 272
use FILL  FILL169050x4050
timestamp 1701859473
transform 1 0 11270 0 1 270
box -12 -8 32 272
use FILL  FILL169050x7950
timestamp 1701859473
transform -1 0 11290 0 -1 790
box -12 -8 32 272
use FILL  FILL169050x11850
timestamp 1701859473
transform 1 0 11270 0 1 790
box -12 -8 32 272
use FILL  FILL169050x15750
timestamp 1701859473
transform -1 0 11290 0 -1 1310
box -12 -8 32 272
use FILL  FILL169050x23550
timestamp 1701859473
transform -1 0 11290 0 -1 1830
box -12 -8 32 272
use FILL  FILL169050x27450
timestamp 1701859473
transform 1 0 11270 0 1 1830
box -12 -8 32 272
use FILL  FILL169050x35250
timestamp 1701859473
transform 1 0 11270 0 1 2350
box -12 -8 32 272
use FILL  FILL169050x39150
timestamp 1701859473
transform -1 0 11290 0 -1 2870
box -12 -8 32 272
use FILL  FILL169050x43050
timestamp 1701859473
transform 1 0 11270 0 1 2870
box -12 -8 32 272
use FILL  FILL169050x46950
timestamp 1701859473
transform -1 0 11290 0 -1 3390
box -12 -8 32 272
use FILL  FILL169050x50850
timestamp 1701859473
transform 1 0 11270 0 1 3390
box -12 -8 32 272
use FILL  FILL169050x54750
timestamp 1701859473
transform -1 0 11290 0 -1 3910
box -12 -8 32 272
use FILL  FILL169050x58650
timestamp 1701859473
transform 1 0 11270 0 1 3910
box -12 -8 32 272
use FILL  FILL169050x62550
timestamp 1701859473
transform -1 0 11290 0 -1 4430
box -12 -8 32 272
use FILL  FILL169050x66450
timestamp 1701859473
transform 1 0 11270 0 1 4430
box -12 -8 32 272
use FILL  FILL169050x70350
timestamp 1701859473
transform -1 0 11290 0 -1 4950
box -12 -8 32 272
use FILL  FILL169050x78150
timestamp 1701859473
transform -1 0 11290 0 -1 5470
box -12 -8 32 272
use FILL  FILL169050x82050
timestamp 1701859473
transform 1 0 11270 0 1 5470
box -12 -8 32 272
use FILL  FILL169050x89850
timestamp 1701859473
transform 1 0 11270 0 1 5990
box -12 -8 32 272
use FILL  FILL169050x93750
timestamp 1701859473
transform -1 0 11290 0 -1 6510
box -12 -8 32 272
use FILL  FILL169050x105450
timestamp 1701859473
transform 1 0 11270 0 1 7030
box -12 -8 32 272
use FILL  FILL169050x109350
timestamp 1701859473
transform -1 0 11290 0 -1 7550
box -12 -8 32 272
use FILL  FILL169050x113250
timestamp 1701859473
transform 1 0 11270 0 1 7550
box -12 -8 32 272
use FILL  FILL169050x121050
timestamp 1701859473
transform 1 0 11270 0 1 8070
box -12 -8 32 272
use FILL  FILL169050x124950
timestamp 1701859473
transform -1 0 11290 0 -1 8590
box -12 -8 32 272
use FILL  FILL169050x132750
timestamp 1701859473
transform -1 0 11290 0 -1 9110
box -12 -8 32 272
use FILL  FILL169050x144450
timestamp 1701859473
transform 1 0 11270 0 1 9630
box -12 -8 32 272
use FILL  FILL169050x156150
timestamp 1701859473
transform -1 0 11290 0 -1 10670
box -12 -8 32 272
use FILL  FILL169050x160050
timestamp 1701859473
transform 1 0 11270 0 1 10670
box -12 -8 32 272
use FILL  FILL169050x163950
timestamp 1701859473
transform -1 0 11290 0 -1 11190
box -12 -8 32 272
use FILL  FILL169350x150
timestamp 1701859473
transform -1 0 11310 0 -1 270
box -12 -8 32 272
use FILL  FILL169350x4050
timestamp 1701859473
transform 1 0 11290 0 1 270
box -12 -8 32 272
use FILL  FILL169350x7950
timestamp 1701859473
transform -1 0 11310 0 -1 790
box -12 -8 32 272
use FILL  FILL169350x11850
timestamp 1701859473
transform 1 0 11290 0 1 790
box -12 -8 32 272
use FILL  FILL169350x15750
timestamp 1701859473
transform -1 0 11310 0 -1 1310
box -12 -8 32 272
use FILL  FILL169350x19650
timestamp 1701859473
transform 1 0 11290 0 1 1310
box -12 -8 32 272
use FILL  FILL169350x23550
timestamp 1701859473
transform -1 0 11310 0 -1 1830
box -12 -8 32 272
use FILL  FILL169350x27450
timestamp 1701859473
transform 1 0 11290 0 1 1830
box -12 -8 32 272
use FILL  FILL169350x35250
timestamp 1701859473
transform 1 0 11290 0 1 2350
box -12 -8 32 272
use FILL  FILL169350x39150
timestamp 1701859473
transform -1 0 11310 0 -1 2870
box -12 -8 32 272
use FILL  FILL169350x43050
timestamp 1701859473
transform 1 0 11290 0 1 2870
box -12 -8 32 272
use FILL  FILL169350x46950
timestamp 1701859473
transform -1 0 11310 0 -1 3390
box -12 -8 32 272
use FILL  FILL169350x50850
timestamp 1701859473
transform 1 0 11290 0 1 3390
box -12 -8 32 272
use FILL  FILL169350x54750
timestamp 1701859473
transform -1 0 11310 0 -1 3910
box -12 -8 32 272
use FILL  FILL169350x58650
timestamp 1701859473
transform 1 0 11290 0 1 3910
box -12 -8 32 272
use FILL  FILL169350x62550
timestamp 1701859473
transform -1 0 11310 0 -1 4430
box -12 -8 32 272
use FILL  FILL169350x66450
timestamp 1701859473
transform 1 0 11290 0 1 4430
box -12 -8 32 272
use FILL  FILL169350x70350
timestamp 1701859473
transform -1 0 11310 0 -1 4950
box -12 -8 32 272
use FILL  FILL169350x74250
timestamp 1701859473
transform 1 0 11290 0 1 4950
box -12 -8 32 272
use FILL  FILL169350x78150
timestamp 1701859473
transform -1 0 11310 0 -1 5470
box -12 -8 32 272
use FILL  FILL169350x82050
timestamp 1701859473
transform 1 0 11290 0 1 5470
box -12 -8 32 272
use FILL  FILL169350x89850
timestamp 1701859473
transform 1 0 11290 0 1 5990
box -12 -8 32 272
use FILL  FILL169350x93750
timestamp 1701859473
transform -1 0 11310 0 -1 6510
box -12 -8 32 272
use FILL  FILL169350x101550
timestamp 1701859473
transform -1 0 11310 0 -1 7030
box -12 -8 32 272
use FILL  FILL169350x105450
timestamp 1701859473
transform 1 0 11290 0 1 7030
box -12 -8 32 272
use FILL  FILL169350x109350
timestamp 1701859473
transform -1 0 11310 0 -1 7550
box -12 -8 32 272
use FILL  FILL169350x113250
timestamp 1701859473
transform 1 0 11290 0 1 7550
box -12 -8 32 272
use FILL  FILL169350x121050
timestamp 1701859473
transform 1 0 11290 0 1 8070
box -12 -8 32 272
use FILL  FILL169350x124950
timestamp 1701859473
transform -1 0 11310 0 -1 8590
box -12 -8 32 272
use FILL  FILL169350x128850
timestamp 1701859473
transform 1 0 11290 0 1 8590
box -12 -8 32 272
use FILL  FILL169350x132750
timestamp 1701859473
transform -1 0 11310 0 -1 9110
box -12 -8 32 272
use FILL  FILL169350x140550
timestamp 1701859473
transform -1 0 11310 0 -1 9630
box -12 -8 32 272
use FILL  FILL169350x144450
timestamp 1701859473
transform 1 0 11290 0 1 9630
box -12 -8 32 272
use FILL  FILL169350x156150
timestamp 1701859473
transform -1 0 11310 0 -1 10670
box -12 -8 32 272
use FILL  FILL169350x160050
timestamp 1701859473
transform 1 0 11290 0 1 10670
box -12 -8 32 272
use FILL  FILL169350x163950
timestamp 1701859473
transform -1 0 11310 0 -1 11190
box -12 -8 32 272
use FILL  FILL169650x150
timestamp 1701859473
transform -1 0 11330 0 -1 270
box -12 -8 32 272
use FILL  FILL169650x4050
timestamp 1701859473
transform 1 0 11310 0 1 270
box -12 -8 32 272
use FILL  FILL169650x7950
timestamp 1701859473
transform -1 0 11330 0 -1 790
box -12 -8 32 272
use FILL  FILL169650x11850
timestamp 1701859473
transform 1 0 11310 0 1 790
box -12 -8 32 272
use FILL  FILL169650x15750
timestamp 1701859473
transform -1 0 11330 0 -1 1310
box -12 -8 32 272
use FILL  FILL169650x19650
timestamp 1701859473
transform 1 0 11310 0 1 1310
box -12 -8 32 272
use FILL  FILL169650x23550
timestamp 1701859473
transform -1 0 11330 0 -1 1830
box -12 -8 32 272
use FILL  FILL169650x27450
timestamp 1701859473
transform 1 0 11310 0 1 1830
box -12 -8 32 272
use FILL  FILL169650x31350
timestamp 1701859473
transform -1 0 11330 0 -1 2350
box -12 -8 32 272
use FILL  FILL169650x35250
timestamp 1701859473
transform 1 0 11310 0 1 2350
box -12 -8 32 272
use FILL  FILL169650x39150
timestamp 1701859473
transform -1 0 11330 0 -1 2870
box -12 -8 32 272
use FILL  FILL169650x43050
timestamp 1701859473
transform 1 0 11310 0 1 2870
box -12 -8 32 272
use FILL  FILL169650x46950
timestamp 1701859473
transform -1 0 11330 0 -1 3390
box -12 -8 32 272
use FILL  FILL169650x50850
timestamp 1701859473
transform 1 0 11310 0 1 3390
box -12 -8 32 272
use FILL  FILL169650x54750
timestamp 1701859473
transform -1 0 11330 0 -1 3910
box -12 -8 32 272
use FILL  FILL169650x58650
timestamp 1701859473
transform 1 0 11310 0 1 3910
box -12 -8 32 272
use FILL  FILL169650x62550
timestamp 1701859473
transform -1 0 11330 0 -1 4430
box -12 -8 32 272
use FILL  FILL169650x66450
timestamp 1701859473
transform 1 0 11310 0 1 4430
box -12 -8 32 272
use FILL  FILL169650x70350
timestamp 1701859473
transform -1 0 11330 0 -1 4950
box -12 -8 32 272
use FILL  FILL169650x74250
timestamp 1701859473
transform 1 0 11310 0 1 4950
box -12 -8 32 272
use FILL  FILL169650x78150
timestamp 1701859473
transform -1 0 11330 0 -1 5470
box -12 -8 32 272
use FILL  FILL169650x82050
timestamp 1701859473
transform 1 0 11310 0 1 5470
box -12 -8 32 272
use FILL  FILL169650x89850
timestamp 1701859473
transform 1 0 11310 0 1 5990
box -12 -8 32 272
use FILL  FILL169650x93750
timestamp 1701859473
transform -1 0 11330 0 -1 6510
box -12 -8 32 272
use FILL  FILL169650x97650
timestamp 1701859473
transform 1 0 11310 0 1 6510
box -12 -8 32 272
use FILL  FILL169650x101550
timestamp 1701859473
transform -1 0 11330 0 -1 7030
box -12 -8 32 272
use FILL  FILL169650x105450
timestamp 1701859473
transform 1 0 11310 0 1 7030
box -12 -8 32 272
use FILL  FILL169650x109350
timestamp 1701859473
transform -1 0 11330 0 -1 7550
box -12 -8 32 272
use FILL  FILL169650x113250
timestamp 1701859473
transform 1 0 11310 0 1 7550
box -12 -8 32 272
use FILL  FILL169650x121050
timestamp 1701859473
transform 1 0 11310 0 1 8070
box -12 -8 32 272
use FILL  FILL169650x124950
timestamp 1701859473
transform -1 0 11330 0 -1 8590
box -12 -8 32 272
use FILL  FILL169650x128850
timestamp 1701859473
transform 1 0 11310 0 1 8590
box -12 -8 32 272
use FILL  FILL169650x132750
timestamp 1701859473
transform -1 0 11330 0 -1 9110
box -12 -8 32 272
use FILL  FILL169650x140550
timestamp 1701859473
transform -1 0 11330 0 -1 9630
box -12 -8 32 272
use FILL  FILL169650x144450
timestamp 1701859473
transform 1 0 11310 0 1 9630
box -12 -8 32 272
use FILL  FILL169650x148350
timestamp 1701859473
transform -1 0 11330 0 -1 10150
box -12 -8 32 272
use FILL  FILL169650x152250
timestamp 1701859473
transform 1 0 11310 0 1 10150
box -12 -8 32 272
use FILL  FILL169650x156150
timestamp 1701859473
transform -1 0 11330 0 -1 10670
box -12 -8 32 272
use FILL  FILL169650x160050
timestamp 1701859473
transform 1 0 11310 0 1 10670
box -12 -8 32 272
use FILL  FILL169650x163950
timestamp 1701859473
transform -1 0 11330 0 -1 11190
box -12 -8 32 272
use FILL  FILL_0__1668_
timestamp 1701859473
transform 1 0 6690 0 -1 3390
box -12 -8 32 272
use FILL  FILL_0__1669_
timestamp 1701859473
transform -1 0 6730 0 -1 790
box -12 -8 32 272
use FILL  FILL_0__1670_
timestamp 1701859473
transform 1 0 6510 0 -1 2870
box -12 -8 32 272
use FILL  FILL_0__1671_
timestamp 1701859473
transform -1 0 6310 0 -1 8590
box -12 -8 32 272
use FILL  FILL_0__1672_
timestamp 1701859473
transform 1 0 5870 0 -1 10670
box -12 -8 32 272
use FILL  FILL_0__1673_
timestamp 1701859473
transform 1 0 6270 0 1 8590
box -12 -8 32 272
use FILL  FILL_0__1674_
timestamp 1701859473
transform -1 0 6350 0 -1 9110
box -12 -8 32 272
use FILL  FILL_0__1675_
timestamp 1701859473
transform 1 0 10 0 -1 5470
box -12 -8 32 272
use FILL  FILL_0__1676_
timestamp 1701859473
transform -1 0 250 0 -1 5470
box -12 -8 32 272
use FILL  FILL_0__1677_
timestamp 1701859473
transform -1 0 490 0 1 5470
box -12 -8 32 272
use FILL  FILL_0__1678_
timestamp 1701859473
transform 1 0 10 0 -1 10670
box -12 -8 32 272
use FILL  FILL_0__1679_
timestamp 1701859473
transform -1 0 230 0 -1 11190
box -12 -8 32 272
use FILL  FILL_0__1680_
timestamp 1701859473
transform 1 0 210 0 -1 10670
box -12 -8 32 272
use FILL  FILL_0__1681_
timestamp 1701859473
transform -1 0 30 0 -1 7030
box -12 -8 32 272
use FILL  FILL_0__1682_
timestamp 1701859473
transform -1 0 30 0 1 7030
box -12 -8 32 272
use FILL  FILL_0__1683_
timestamp 1701859473
transform 1 0 10 0 1 6510
box -12 -8 32 272
use FILL  FILL_0__1684_
timestamp 1701859473
transform 1 0 890 0 -1 11190
box -12 -8 32 272
use FILL  FILL_0__1685_
timestamp 1701859473
transform -1 0 1150 0 -1 11190
box -12 -8 32 272
use FILL  FILL_0__1686_
timestamp 1701859473
transform -1 0 950 0 1 10670
box -12 -8 32 272
use FILL  FILL_0__1687_
timestamp 1701859473
transform 1 0 1370 0 -1 11190
box -12 -8 32 272
use FILL  FILL_0__1688_
timestamp 1701859473
transform -1 0 1630 0 -1 11190
box -12 -8 32 272
use FILL  FILL_0__1689_
timestamp 1701859473
transform -1 0 1890 0 1 10150
box -12 -8 32 272
use FILL  FILL_0__1690_
timestamp 1701859473
transform 1 0 2050 0 1 9110
box -12 -8 32 272
use FILL  FILL_0__1691_
timestamp 1701859473
transform -1 0 2070 0 -1 9110
box -12 -8 32 272
use FILL  FILL_0__1692_
timestamp 1701859473
transform 1 0 10 0 1 790
box -12 -8 32 272
use FILL  FILL_0__1693_
timestamp 1701859473
transform 1 0 10 0 -1 1310
box -12 -8 32 272
use FILL  FILL_0__1694_
timestamp 1701859473
transform 1 0 430 0 -1 270
box -12 -8 32 272
use FILL  FILL_0__1695_
timestamp 1701859473
transform -1 0 650 0 -1 270
box -12 -8 32 272
use FILL  FILL_0__1696_
timestamp 1701859473
transform 1 0 1070 0 1 2870
box -12 -8 32 272
use FILL  FILL_0__1697_
timestamp 1701859473
transform -1 0 2730 0 -1 2870
box -12 -8 32 272
use FILL  FILL_0__1698_
timestamp 1701859473
transform -1 0 1830 0 1 3390
box -12 -8 32 272
use FILL  FILL_0__1699_
timestamp 1701859473
transform 1 0 3750 0 1 3390
box -12 -8 32 272
use FILL  FILL_0__1700_
timestamp 1701859473
transform -1 0 2550 0 -1 3910
box -12 -8 32 272
use FILL  FILL_0__1701_
timestamp 1701859473
transform -1 0 1090 0 1 270
box -12 -8 32 272
use FILL  FILL_0__1702_
timestamp 1701859473
transform 1 0 850 0 1 270
box -12 -8 32 272
use FILL  FILL_0__1703_
timestamp 1701859473
transform -1 0 1330 0 1 1830
box -12 -8 32 272
use FILL  FILL_0__1704_
timestamp 1701859473
transform -1 0 9090 0 1 2870
box -12 -8 32 272
use FILL  FILL_0__1705_
timestamp 1701859473
transform 1 0 9710 0 -1 790
box -12 -8 32 272
use FILL  FILL_0__1706_
timestamp 1701859473
transform -1 0 7930 0 -1 4950
box -12 -8 32 272
use FILL  FILL_0__1707_
timestamp 1701859473
transform 1 0 8370 0 -1 4950
box -12 -8 32 272
use FILL  FILL_0__1708_
timestamp 1701859473
transform 1 0 4990 0 -1 5990
box -12 -8 32 272
use FILL  FILL_0__1709_
timestamp 1701859473
transform -1 0 11090 0 1 5990
box -12 -8 32 272
use FILL  FILL_0__1710_
timestamp 1701859473
transform 1 0 5370 0 -1 5470
box -12 -8 32 272
use FILL  FILL_0__1711_
timestamp 1701859473
transform -1 0 5210 0 -1 5990
box -12 -8 32 272
use FILL  FILL_0__1712_
timestamp 1701859473
transform -1 0 5030 0 1 5470
box -12 -8 32 272
use FILL  FILL_0__1713_
timestamp 1701859473
transform 1 0 7890 0 1 4430
box -12 -8 32 272
use FILL  FILL_0__1714_
timestamp 1701859473
transform 1 0 7690 0 1 4950
box -12 -8 32 272
use FILL  FILL_0__1715_
timestamp 1701859473
transform -1 0 7930 0 1 4950
box -12 -8 32 272
use FILL  FILL_0__1716_
timestamp 1701859473
transform -1 0 8150 0 1 4430
box -12 -8 32 272
use FILL  FILL_0__1717_
timestamp 1701859473
transform -1 0 7930 0 1 1310
box -12 -8 32 272
use FILL  FILL_0__1718_
timestamp 1701859473
transform -1 0 5870 0 1 5990
box -12 -8 32 272
use FILL  FILL_0__1719_
timestamp 1701859473
transform -1 0 6730 0 -1 5990
box -12 -8 32 272
use FILL  FILL_0__1720_
timestamp 1701859473
transform -1 0 6710 0 1 5470
box -12 -8 32 272
use FILL  FILL_0__1721_
timestamp 1701859473
transform -1 0 6950 0 1 5470
box -12 -8 32 272
use FILL  FILL_0__1722_
timestamp 1701859473
transform -1 0 7650 0 1 4430
box -12 -8 32 272
use FILL  FILL_0__1723_
timestamp 1701859473
transform 1 0 7870 0 1 1830
box -12 -8 32 272
use FILL  FILL_0__1724_
timestamp 1701859473
transform -1 0 7910 0 -1 1310
box -12 -8 32 272
use FILL  FILL_0__1725_
timestamp 1701859473
transform 1 0 6510 0 1 5990
box -12 -8 32 272
use FILL  FILL_0__1726_
timestamp 1701859473
transform 1 0 6710 0 1 5990
box -12 -8 32 272
use FILL  FILL_0__1727_
timestamp 1701859473
transform -1 0 6950 0 1 5990
box -12 -8 32 272
use FILL  FILL_0__1728_
timestamp 1701859473
transform 1 0 7650 0 1 5990
box -12 -8 32 272
use FILL  FILL_0__1729_
timestamp 1701859473
transform -1 0 7590 0 -1 5990
box -12 -8 32 272
use FILL  FILL_0__1730_
timestamp 1701859473
transform -1 0 8070 0 1 3390
box -12 -8 32 272
use FILL  FILL_0__1731_
timestamp 1701859473
transform -1 0 7930 0 -1 270
box -12 -8 32 272
use FILL  FILL_0__1732_
timestamp 1701859473
transform -1 0 7890 0 1 5470
box -12 -8 32 272
use FILL  FILL_0__1733_
timestamp 1701859473
transform -1 0 8110 0 1 5470
box -12 -8 32 272
use FILL  FILL_0__1734_
timestamp 1701859473
transform 1 0 8070 0 -1 5470
box -12 -8 32 272
use FILL  FILL_0__1735_
timestamp 1701859473
transform 1 0 8530 0 -1 5470
box -12 -8 32 272
use FILL  FILL_0__1736_
timestamp 1701859473
transform 1 0 8370 0 1 4950
box -12 -8 32 272
use FILL  FILL_0__1737_
timestamp 1701859473
transform -1 0 8450 0 -1 3910
box -12 -8 32 272
use FILL  FILL_0__1738_
timestamp 1701859473
transform 1 0 8850 0 1 790
box -12 -8 32 272
use FILL  FILL_0__1739_
timestamp 1701859473
transform -1 0 9070 0 -1 790
box -12 -8 32 272
use FILL  FILL_0__1740_
timestamp 1701859473
transform 1 0 6430 0 1 270
box -12 -8 32 272
use FILL  FILL_0__1741_
timestamp 1701859473
transform 1 0 6330 0 1 790
box -12 -8 32 272
use FILL  FILL_0__1742_
timestamp 1701859473
transform -1 0 6270 0 -1 790
box -12 -8 32 272
use FILL  FILL_0__1743_
timestamp 1701859473
transform -1 0 2270 0 -1 3390
box -12 -8 32 272
use FILL  FILL_0__1744_
timestamp 1701859473
transform 1 0 250 0 -1 4950
box -12 -8 32 272
use FILL  FILL_0__1745_
timestamp 1701859473
transform 1 0 2070 0 -1 3910
box -12 -8 32 272
use FILL  FILL_0__1746_
timestamp 1701859473
transform -1 0 5090 0 -1 3390
box -12 -8 32 272
use FILL  FILL_0__1747_
timestamp 1701859473
transform -1 0 250 0 -1 270
box -12 -8 32 272
use FILL  FILL_0__1748_
timestamp 1701859473
transform -1 0 450 0 1 270
box -12 -8 32 272
use FILL  FILL_0__1749_
timestamp 1701859473
transform -1 0 890 0 1 1310
box -12 -8 32 272
use FILL  FILL_0__1750_
timestamp 1701859473
transform -1 0 1110 0 1 1310
box -12 -8 32 272
use FILL  FILL_0__1751_
timestamp 1701859473
transform -1 0 4470 0 -1 2870
box -12 -8 32 272
use FILL  FILL_0__1752_
timestamp 1701859473
transform 1 0 4670 0 -1 2870
box -12 -8 32 272
use FILL  FILL_0__1753_
timestamp 1701859473
transform -1 0 4290 0 1 790
box -12 -8 32 272
use FILL  FILL_0__1754_
timestamp 1701859473
transform 1 0 230 0 -1 790
box -12 -8 32 272
use FILL  FILL_0__1755_
timestamp 1701859473
transform -1 0 450 0 -1 790
box -12 -8 32 272
use FILL  FILL_0__1756_
timestamp 1701859473
transform -1 0 30 0 -1 270
box -12 -8 32 272
use FILL  FILL_0__1757_
timestamp 1701859473
transform 1 0 630 0 -1 790
box -12 -8 32 272
use FILL  FILL_0__1758_
timestamp 1701859473
transform 1 0 10 0 1 2350
box -12 -8 32 272
use FILL  FILL_0__1759_
timestamp 1701859473
transform -1 0 2510 0 -1 2870
box -12 -8 32 272
use FILL  FILL_0__1760_
timestamp 1701859473
transform 1 0 2890 0 -1 2870
box -12 -8 32 272
use FILL  FILL_0__1761_
timestamp 1701859473
transform -1 0 3210 0 -1 3390
box -12 -8 32 272
use FILL  FILL_0__1762_
timestamp 1701859473
transform -1 0 30 0 1 270
box -12 -8 32 272
use FILL  FILL_0__1763_
timestamp 1701859473
transform 1 0 10 0 -1 790
box -12 -8 32 272
use FILL  FILL_0__1764_
timestamp 1701859473
transform 1 0 450 0 1 1310
box -12 -8 32 272
use FILL  FILL_0__1765_
timestamp 1701859473
transform 1 0 1310 0 1 1310
box -12 -8 32 272
use FILL  FILL_0__1766_
timestamp 1701859473
transform -1 0 3110 0 -1 1830
box -12 -8 32 272
use FILL  FILL_0__1767_
timestamp 1701859473
transform 1 0 1410 0 -1 4430
box -12 -8 32 272
use FILL  FILL_0__1768_
timestamp 1701859473
transform 1 0 230 0 -1 1310
box -12 -8 32 272
use FILL  FILL_0__1769_
timestamp 1701859473
transform -1 0 450 0 1 1830
box -12 -8 32 272
use FILL  FILL_0__1770_
timestamp 1701859473
transform 1 0 2050 0 -1 3390
box -12 -8 32 272
use FILL  FILL_0__1771_
timestamp 1701859473
transform -1 0 2310 0 -1 3910
box -12 -8 32 272
use FILL  FILL_0__1772_
timestamp 1701859473
transform -1 0 2970 0 -1 3910
box -12 -8 32 272
use FILL  FILL_0__1773_
timestamp 1701859473
transform 1 0 3870 0 1 2870
box -12 -8 32 272
use FILL  FILL_0__1774_
timestamp 1701859473
transform -1 0 5250 0 -1 2350
box -12 -8 32 272
use FILL  FILL_0__1775_
timestamp 1701859473
transform 1 0 210 0 1 790
box -12 -8 32 272
use FILL  FILL_0__1776_
timestamp 1701859473
transform -1 0 250 0 1 1310
box -12 -8 32 272
use FILL  FILL_0__1777_
timestamp 1701859473
transform 1 0 670 0 -1 1830
box -12 -8 32 272
use FILL  FILL_0__1778_
timestamp 1701859473
transform -1 0 4390 0 1 5470
box -12 -8 32 272
use FILL  FILL_0__1779_
timestamp 1701859473
transform -1 0 6030 0 -1 5470
box -12 -8 32 272
use FILL  FILL_0__1780_
timestamp 1701859473
transform 1 0 4750 0 1 2870
box -12 -8 32 272
use FILL  FILL_0__1781_
timestamp 1701859473
transform 1 0 4330 0 1 2870
box -12 -8 32 272
use FILL  FILL_0__1782_
timestamp 1701859473
transform -1 0 30 0 1 1310
box -12 -8 32 272
use FILL  FILL_0__1783_
timestamp 1701859473
transform -1 0 1310 0 1 2870
box -12 -8 32 272
use FILL  FILL_0__1784_
timestamp 1701859473
transform -1 0 5010 0 1 2870
box -12 -8 32 272
use FILL  FILL_0__1785_
timestamp 1701859473
transform 1 0 4930 0 -1 2870
box -12 -8 32 272
use FILL  FILL_0__1786_
timestamp 1701859473
transform -1 0 5010 0 -1 2350
box -12 -8 32 272
use FILL  FILL_0__1787_
timestamp 1701859473
transform 1 0 4990 0 1 2350
box -12 -8 32 272
use FILL  FILL_0__1788_
timestamp 1701859473
transform -1 0 4790 0 -1 2350
box -12 -8 32 272
use FILL  FILL_0__1789_
timestamp 1701859473
transform 1 0 10 0 1 1830
box -12 -8 32 272
use FILL  FILL_0__1790_
timestamp 1701859473
transform -1 0 250 0 -1 2350
box -12 -8 32 272
use FILL  FILL_0__1791_
timestamp 1701859473
transform -1 0 2050 0 -1 2350
box -12 -8 32 272
use FILL  FILL_0__1792_
timestamp 1701859473
transform -1 0 3430 0 -1 2350
box -12 -8 32 272
use FILL  FILL_0__1793_
timestamp 1701859473
transform -1 0 4530 0 1 1830
box -12 -8 32 272
use FILL  FILL_0__1794_
timestamp 1701859473
transform 1 0 850 0 1 1830
box -12 -8 32 272
use FILL  FILL_0__1795_
timestamp 1701859473
transform -1 0 2110 0 1 2350
box -12 -8 32 272
use FILL  FILL_0__1796_
timestamp 1701859473
transform -1 0 1730 0 -1 1830
box -12 -8 32 272
use FILL  FILL_0__1797_
timestamp 1701859473
transform 1 0 1950 0 -1 1830
box -12 -8 32 272
use FILL  FILL_0__1798_
timestamp 1701859473
transform 1 0 870 0 -1 1310
box -12 -8 32 272
use FILL  FILL_0__1799_
timestamp 1701859473
transform 1 0 3690 0 1 3910
box -12 -8 32 272
use FILL  FILL_0__1800_
timestamp 1701859473
transform 1 0 3370 0 1 1830
box -12 -8 32 272
use FILL  FILL_0__1801_
timestamp 1701859473
transform -1 0 1110 0 1 1830
box -12 -8 32 272
use FILL  FILL_0__1802_
timestamp 1701859473
transform -1 0 3650 0 1 2350
box -12 -8 32 272
use FILL  FILL_0__1803_
timestamp 1701859473
transform -1 0 3870 0 1 2350
box -12 -8 32 272
use FILL  FILL_0__1804_
timestamp 1701859473
transform -1 0 4110 0 1 2350
box -12 -8 32 272
use FILL  FILL_0__1805_
timestamp 1701859473
transform 1 0 5410 0 1 2350
box -12 -8 32 272
use FILL  FILL_0__1806_
timestamp 1701859473
transform -1 0 4810 0 1 2350
box -12 -8 32 272
use FILL  FILL_0__1807_
timestamp 1701859473
transform -1 0 5210 0 1 2350
box -12 -8 32 272
use FILL  FILL_0__1808_
timestamp 1701859473
transform 1 0 4730 0 1 1830
box -12 -8 32 272
use FILL  FILL_0__1809_
timestamp 1701859473
transform -1 0 7090 0 -1 270
box -12 -8 32 272
use FILL  FILL_0__1810_
timestamp 1701859473
transform -1 0 7070 0 1 1310
box -12 -8 32 272
use FILL  FILL_0__1811_
timestamp 1701859473
transform 1 0 7410 0 -1 1830
box -12 -8 32 272
use FILL  FILL_0__1812_
timestamp 1701859473
transform -1 0 7490 0 -1 1310
box -12 -8 32 272
use FILL  FILL_0__1813_
timestamp 1701859473
transform 1 0 9070 0 1 790
box -12 -8 32 272
use FILL  FILL_0__1814_
timestamp 1701859473
transform -1 0 8110 0 -1 1830
box -12 -8 32 272
use FILL  FILL_0__1815_
timestamp 1701859473
transform 1 0 8310 0 1 2350
box -12 -8 32 272
use FILL  FILL_0__1816_
timestamp 1701859473
transform -1 0 9590 0 -1 2350
box -12 -8 32 272
use FILL  FILL_0__1817_
timestamp 1701859473
transform -1 0 9310 0 1 1310
box -12 -8 32 272
use FILL  FILL_0__1818_
timestamp 1701859473
transform -1 0 9510 0 1 270
box -12 -8 32 272
use FILL  FILL_0__1819_
timestamp 1701859473
transform -1 0 8330 0 -1 1830
box -12 -8 32 272
use FILL  FILL_0__1820_
timestamp 1701859473
transform -1 0 8410 0 1 1310
box -12 -8 32 272
use FILL  FILL_0__1821_
timestamp 1701859473
transform -1 0 4850 0 1 1310
box -12 -8 32 272
use FILL  FILL_0__1822_
timestamp 1701859473
transform -1 0 4650 0 -1 790
box -12 -8 32 272
use FILL  FILL_0__1823_
timestamp 1701859473
transform -1 0 4190 0 -1 790
box -12 -8 32 272
use FILL  FILL_0__1824_
timestamp 1701859473
transform 1 0 4570 0 1 2350
box -12 -8 32 272
use FILL  FILL_0__1825_
timestamp 1701859473
transform 1 0 5630 0 1 1830
box -12 -8 32 272
use FILL  FILL_0__1826_
timestamp 1701859473
transform 1 0 8130 0 -1 270
box -12 -8 32 272
use FILL  FILL_0__1827_
timestamp 1701859473
transform 1 0 9270 0 -1 790
box -12 -8 32 272
use FILL  FILL_0__1828_
timestamp 1701859473
transform 1 0 8430 0 1 270
box -12 -8 32 272
use FILL  FILL_0__1829_
timestamp 1701859473
transform 1 0 5730 0 1 270
box -12 -8 32 272
use FILL  FILL_0__1830_
timestamp 1701859473
transform 1 0 3170 0 1 4430
box -12 -8 32 272
use FILL  FILL_0__1831_
timestamp 1701859473
transform -1 0 7950 0 -1 790
box -12 -8 32 272
use FILL  FILL_0__1832_
timestamp 1701859473
transform 1 0 6450 0 -1 790
box -12 -8 32 272
use FILL  FILL_0__1833_
timestamp 1701859473
transform -1 0 650 0 1 270
box -12 -8 32 272
use FILL  FILL_0__1834_
timestamp 1701859473
transform 1 0 1090 0 -1 1310
box -12 -8 32 272
use FILL  FILL_0__1835_
timestamp 1701859473
transform -1 0 2470 0 -1 1310
box -12 -8 32 272
use FILL  FILL_0__1836_
timestamp 1701859473
transform 1 0 1030 0 1 790
box -12 -8 32 272
use FILL  FILL_0__1837_
timestamp 1701859473
transform -1 0 2430 0 1 790
box -12 -8 32 272
use FILL  FILL_0__1838_
timestamp 1701859473
transform 1 0 2170 0 1 790
box -12 -8 32 272
use FILL  FILL_0__1839_
timestamp 1701859473
transform -1 0 230 0 1 270
box -12 -8 32 272
use FILL  FILL_0__1840_
timestamp 1701859473
transform -1 0 870 0 1 2870
box -12 -8 32 272
use FILL  FILL_0__1841_
timestamp 1701859473
transform 1 0 3650 0 1 2870
box -12 -8 32 272
use FILL  FILL_0__1842_
timestamp 1701859473
transform -1 0 2910 0 -1 1830
box -12 -8 32 272
use FILL  FILL_0__1843_
timestamp 1701859473
transform -1 0 3870 0 -1 2350
box -12 -8 32 272
use FILL  FILL_0__1844_
timestamp 1701859473
transform 1 0 3770 0 -1 2870
box -12 -8 32 272
use FILL  FILL_0__1845_
timestamp 1701859473
transform -1 0 1710 0 -1 4950
box -12 -8 32 272
use FILL  FILL_0__1846_
timestamp 1701859473
transform 1 0 4070 0 1 4430
box -12 -8 32 272
use FILL  FILL_0__1847_
timestamp 1701859473
transform 1 0 3390 0 1 4430
box -12 -8 32 272
use FILL  FILL_0__1848_
timestamp 1701859473
transform 1 0 3830 0 1 4430
box -12 -8 32 272
use FILL  FILL_0__1849_
timestamp 1701859473
transform -1 0 4030 0 -1 2870
box -12 -8 32 272
use FILL  FILL_0__1850_
timestamp 1701859473
transform -1 0 850 0 1 790
box -12 -8 32 272
use FILL  FILL_0__1851_
timestamp 1701859473
transform 1 0 1510 0 -1 1830
box -12 -8 32 272
use FILL  FILL_0__1852_
timestamp 1701859473
transform -1 0 2330 0 1 2350
box -12 -8 32 272
use FILL  FILL_0__1853_
timestamp 1701859473
transform 1 0 10 0 -1 2350
box -12 -8 32 272
use FILL  FILL_0__1854_
timestamp 1701859473
transform 1 0 2250 0 -1 2350
box -12 -8 32 272
use FILL  FILL_0__1855_
timestamp 1701859473
transform -1 0 2510 0 -1 2350
box -12 -8 32 272
use FILL  FILL_0__1856_
timestamp 1701859473
transform 1 0 1410 0 -1 790
box -12 -8 32 272
use FILL  FILL_0__1857_
timestamp 1701859473
transform -1 0 2610 0 -1 790
box -12 -8 32 272
use FILL  FILL_0__1858_
timestamp 1701859473
transform 1 0 2350 0 -1 790
box -12 -8 32 272
use FILL  FILL_0__1859_
timestamp 1701859473
transform 1 0 2130 0 -1 790
box -12 -8 32 272
use FILL  FILL_0__1860_
timestamp 1701859473
transform -1 0 1670 0 -1 790
box -12 -8 32 272
use FILL  FILL_0__1861_
timestamp 1701859473
transform -1 0 1910 0 -1 790
box -12 -8 32 272
use FILL  FILL_0__1862_
timestamp 1701859473
transform -1 0 1990 0 1 270
box -12 -8 32 272
use FILL  FILL_0__1863_
timestamp 1701859473
transform 1 0 2210 0 1 270
box -12 -8 32 272
use FILL  FILL_0__1864_
timestamp 1701859473
transform 1 0 3450 0 1 270
box -12 -8 32 272
use FILL  FILL_0__1865_
timestamp 1701859473
transform 1 0 7250 0 -1 1310
box -12 -8 32 272
use FILL  FILL_0__1866_
timestamp 1701859473
transform 1 0 3610 0 -1 1310
box -12 -8 32 272
use FILL  FILL_0__1867_
timestamp 1701859473
transform 1 0 1070 0 -1 1830
box -12 -8 32 272
use FILL  FILL_0__1868_
timestamp 1701859473
transform 1 0 1510 0 1 1310
box -12 -8 32 272
use FILL  FILL_0__1869_
timestamp 1701859473
transform 1 0 1930 0 1 1310
box -12 -8 32 272
use FILL  FILL_0__1870_
timestamp 1701859473
transform -1 0 1550 0 -1 1310
box -12 -8 32 272
use FILL  FILL_0__1871_
timestamp 1701859473
transform -1 0 2670 0 -1 1310
box -12 -8 32 272
use FILL  FILL_0__1872_
timestamp 1701859473
transform -1 0 450 0 1 790
box -12 -8 32 272
use FILL  FILL_0__1873_
timestamp 1701859473
transform 1 0 630 0 1 790
box -12 -8 32 272
use FILL  FILL_0__1874_
timestamp 1701859473
transform -1 0 1270 0 1 790
box -12 -8 32 272
use FILL  FILL_0__1875_
timestamp 1701859473
transform 1 0 850 0 -1 790
box -12 -8 32 272
use FILL  FILL_0__1876_
timestamp 1701859473
transform 1 0 1170 0 -1 790
box -12 -8 32 272
use FILL  FILL_0__1877_
timestamp 1701859473
transform 1 0 2110 0 1 4950
box -12 -8 32 272
use FILL  FILL_0__1878_
timestamp 1701859473
transform 1 0 450 0 -1 1310
box -12 -8 32 272
use FILL  FILL_0__1879_
timestamp 1701859473
transform 1 0 670 0 1 1310
box -12 -8 32 272
use FILL  FILL_0__1880_
timestamp 1701859473
transform -1 0 1930 0 -1 4950
box -12 -8 32 272
use FILL  FILL_0__1881_
timestamp 1701859473
transform -1 0 2170 0 -1 4950
box -12 -8 32 272
use FILL  FILL_0__1882_
timestamp 1701859473
transform 1 0 1490 0 -1 3390
box -12 -8 32 272
use FILL  FILL_0__1883_
timestamp 1701859473
transform 1 0 970 0 -1 3390
box -12 -8 32 272
use FILL  FILL_0__1884_
timestamp 1701859473
transform -1 0 3990 0 1 3390
box -12 -8 32 272
use FILL  FILL_0__1885_
timestamp 1701859473
transform -1 0 3710 0 -1 3390
box -12 -8 32 272
use FILL  FILL_0__1886_
timestamp 1701859473
transform 1 0 3450 0 -1 3390
box -12 -8 32 272
use FILL  FILL_0__1887_
timestamp 1701859473
transform -1 0 3430 0 1 2870
box -12 -8 32 272
use FILL  FILL_0__1888_
timestamp 1701859473
transform -1 0 2470 0 1 270
box -12 -8 32 272
use FILL  FILL_0__1889_
timestamp 1701859473
transform 1 0 1610 0 -1 2870
box -12 -8 32 272
use FILL  FILL_0__1890_
timestamp 1701859473
transform -1 0 250 0 -1 1830
box -12 -8 32 272
use FILL  FILL_0__1891_
timestamp 1701859473
transform 1 0 10 0 -1 1830
box -12 -8 32 272
use FILL  FILL_0__1892_
timestamp 1701859473
transform 1 0 4850 0 -1 3390
box -12 -8 32 272
use FILL  FILL_0__1893_
timestamp 1701859473
transform 1 0 3850 0 1 1830
box -12 -8 32 272
use FILL  FILL_0__1894_
timestamp 1701859473
transform 1 0 4050 0 1 1830
box -12 -8 32 272
use FILL  FILL_0__1895_
timestamp 1701859473
transform -1 0 1790 0 1 1830
box -12 -8 32 272
use FILL  FILL_0__1896_
timestamp 1701859473
transform 1 0 1810 0 -1 2350
box -12 -8 32 272
use FILL  FILL_0__1897_
timestamp 1701859473
transform 1 0 3430 0 1 2350
box -12 -8 32 272
use FILL  FILL_0__1898_
timestamp 1701859473
transform 1 0 3210 0 1 2350
box -12 -8 32 272
use FILL  FILL_0__1899_
timestamp 1701859473
transform -1 0 3190 0 -1 2350
box -12 -8 32 272
use FILL  FILL_0__1900_
timestamp 1701859473
transform -1 0 4030 0 -1 1830
box -12 -8 32 272
use FILL  FILL_0__1901_
timestamp 1701859473
transform -1 0 670 0 1 1830
box -12 -8 32 272
use FILL  FILL_0__1902_
timestamp 1701859473
transform 1 0 4970 0 1 1830
box -12 -8 32 272
use FILL  FILL_0__1903_
timestamp 1701859473
transform 1 0 3290 0 1 1310
box -12 -8 32 272
use FILL  FILL_0__1904_
timestamp 1701859473
transform -1 0 3390 0 -1 1310
box -12 -8 32 272
use FILL  FILL_0__1905_
timestamp 1701859473
transform 1 0 2930 0 1 270
box -12 -8 32 272
use FILL  FILL_0__1906_
timestamp 1701859473
transform 1 0 210 0 1 2350
box -12 -8 32 272
use FILL  FILL_0__1907_
timestamp 1701859473
transform -1 0 2970 0 -1 2350
box -12 -8 32 272
use FILL  FILL_0__1908_
timestamp 1701859473
transform 1 0 6390 0 -1 2350
box -12 -8 32 272
use FILL  FILL_0__1909_
timestamp 1701859473
transform -1 0 5990 0 -1 2350
box -12 -8 32 272
use FILL  FILL_0__1910_
timestamp 1701859473
transform -1 0 5490 0 -1 2350
box -12 -8 32 272
use FILL  FILL_0__1911_
timestamp 1701859473
transform -1 0 650 0 1 2870
box -12 -8 32 272
use FILL  FILL_0__1912_
timestamp 1701859473
transform -1 0 3250 0 1 3910
box -12 -8 32 272
use FILL  FILL_0__1913_
timestamp 1701859473
transform -1 0 970 0 -1 2870
box -12 -8 32 272
use FILL  FILL_0__1914_
timestamp 1701859473
transform -1 0 1410 0 1 3390
box -12 -8 32 272
use FILL  FILL_0__1915_
timestamp 1701859473
transform 1 0 2490 0 1 3390
box -12 -8 32 272
use FILL  FILL_0__1916_
timestamp 1701859473
transform -1 0 3350 0 1 3390
box -12 -8 32 272
use FILL  FILL_0__1917_
timestamp 1701859473
transform -1 0 4630 0 -1 3390
box -12 -8 32 272
use FILL  FILL_0__1918_
timestamp 1701859473
transform 1 0 1670 0 1 4950
box -12 -8 32 272
use FILL  FILL_0__1919_
timestamp 1701859473
transform -1 0 1190 0 -1 2870
box -12 -8 32 272
use FILL  FILL_0__1920_
timestamp 1701859473
transform -1 0 4970 0 1 4430
box -12 -8 32 272
use FILL  FILL_0__1921_
timestamp 1701859473
transform 1 0 4730 0 1 4430
box -12 -8 32 272
use FILL  FILL_0__1922_
timestamp 1701859473
transform -1 0 4530 0 1 4430
box -12 -8 32 272
use FILL  FILL_0__1923_
timestamp 1701859473
transform 1 0 4390 0 -1 3390
box -12 -8 32 272
use FILL  FILL_0__1924_
timestamp 1701859473
transform 1 0 1890 0 1 4950
box -12 -8 32 272
use FILL  FILL_0__1925_
timestamp 1701859473
transform 1 0 6030 0 -1 4430
box -12 -8 32 272
use FILL  FILL_0__1926_
timestamp 1701859473
transform 1 0 650 0 -1 1310
box -12 -8 32 272
use FILL  FILL_0__1927_
timestamp 1701859473
transform 1 0 2890 0 -1 1310
box -12 -8 32 272
use FILL  FILL_0__1928_
timestamp 1701859473
transform -1 0 3150 0 -1 1310
box -12 -8 32 272
use FILL  FILL_0__1929_
timestamp 1701859473
transform 1 0 3330 0 1 790
box -12 -8 32 272
use FILL  FILL_0__1930_
timestamp 1701859473
transform 1 0 3150 0 1 270
box -12 -8 32 272
use FILL  FILL_0__1931_
timestamp 1701859473
transform 1 0 3750 0 1 270
box -12 -8 32 272
use FILL  FILL_0__1932_
timestamp 1701859473
transform -1 0 3990 0 1 270
box -12 -8 32 272
use FILL  FILL_0__1933_
timestamp 1701859473
transform -1 0 1790 0 1 270
box -12 -8 32 272
use FILL  FILL_0__1934_
timestamp 1701859473
transform -1 0 5410 0 1 790
box -12 -8 32 272
use FILL  FILL_0__1935_
timestamp 1701859473
transform 1 0 5530 0 -1 270
box -12 -8 32 272
use FILL  FILL_0__1936_
timestamp 1701859473
transform -1 0 8290 0 1 3390
box -12 -8 32 272
use FILL  FILL_0__1937_
timestamp 1701859473
transform -1 0 7510 0 -1 270
box -12 -8 32 272
use FILL  FILL_0__1938_
timestamp 1701859473
transform -1 0 7710 0 -1 270
box -12 -8 32 272
use FILL  FILL_0__1939_
timestamp 1701859473
transform -1 0 6630 0 -1 270
box -12 -8 32 272
use FILL  FILL_0__1940_
timestamp 1701859473
transform -1 0 5750 0 -1 270
box -12 -8 32 272
use FILL  FILL_0__1941_
timestamp 1701859473
transform 1 0 5770 0 -1 790
box -12 -8 32 272
use FILL  FILL_0__1942_
timestamp 1701859473
transform 1 0 4750 0 -1 1310
box -12 -8 32 272
use FILL  FILL_0__1943_
timestamp 1701859473
transform 1 0 8010 0 1 270
box -12 -8 32 272
use FILL  FILL_0__1944_
timestamp 1701859473
transform -1 0 8250 0 1 270
box -12 -8 32 272
use FILL  FILL_0__1945_
timestamp 1701859473
transform 1 0 7790 0 1 270
box -12 -8 32 272
use FILL  FILL_0__1946_
timestamp 1701859473
transform -1 0 5990 0 1 270
box -12 -8 32 272
use FILL  FILL_0__1947_
timestamp 1701859473
transform -1 0 6010 0 -1 790
box -12 -8 32 272
use FILL  FILL_0__1948_
timestamp 1701859473
transform 1 0 5290 0 -1 790
box -12 -8 32 272
use FILL  FILL_0__1949_
timestamp 1701859473
transform 1 0 4530 0 -1 1310
box -12 -8 32 272
use FILL  FILL_0__1950_
timestamp 1701859473
transform -1 0 8170 0 -1 790
box -12 -8 32 272
use FILL  FILL_0__1951_
timestamp 1701859473
transform 1 0 450 0 -1 2350
box -12 -8 32 272
use FILL  FILL_0__1952_
timestamp 1701859473
transform -1 0 5630 0 1 2350
box -12 -8 32 272
use FILL  FILL_0__1953_
timestamp 1701859473
transform 1 0 5730 0 -1 2350
box -12 -8 32 272
use FILL  FILL_0__1954_
timestamp 1701859473
transform 1 0 8110 0 -1 1310
box -12 -8 32 272
use FILL  FILL_0__1955_
timestamp 1701859473
transform -1 0 8650 0 1 1310
box -12 -8 32 272
use FILL  FILL_0__1956_
timestamp 1701859473
transform -1 0 6190 0 -1 1310
box -12 -8 32 272
use FILL  FILL_0__1957_
timestamp 1701859473
transform -1 0 5950 0 -1 1310
box -12 -8 32 272
use FILL  FILL_0__1958_
timestamp 1701859473
transform 1 0 5210 0 -1 1310
box -12 -8 32 272
use FILL  FILL_0__1959_
timestamp 1701859473
transform 1 0 5650 0 -1 2870
box -12 -8 32 272
use FILL  FILL_0__1960_
timestamp 1701859473
transform -1 0 6090 0 -1 2870
box -12 -8 32 272
use FILL  FILL_0__1961_
timestamp 1701859473
transform -1 0 4350 0 1 2350
box -12 -8 32 272
use FILL  FILL_0__1962_
timestamp 1701859473
transform 1 0 5810 0 1 2350
box -12 -8 32 272
use FILL  FILL_0__1963_
timestamp 1701859473
transform 1 0 5270 0 1 1310
box -12 -8 32 272
use FILL  FILL_0__1964_
timestamp 1701859473
transform 1 0 9090 0 1 1310
box -12 -8 32 272
use FILL  FILL_0__1965_
timestamp 1701859473
transform 1 0 7490 0 1 790
box -12 -8 32 272
use FILL  FILL_0__1966_
timestamp 1701859473
transform -1 0 7610 0 1 270
box -12 -8 32 272
use FILL  FILL_0__1967_
timestamp 1701859473
transform -1 0 6670 0 1 270
box -12 -8 32 272
use FILL  FILL_0__1968_
timestamp 1701859473
transform 1 0 5450 0 -1 1310
box -12 -8 32 272
use FILL  FILL_0__1969_
timestamp 1701859473
transform 1 0 5650 0 1 2870
box -12 -8 32 272
use FILL  FILL_0__1970_
timestamp 1701859473
transform 1 0 5290 0 -1 3390
box -12 -8 32 272
use FILL  FILL_0__1971_
timestamp 1701859473
transform 1 0 5730 0 1 3910
box -12 -8 32 272
use FILL  FILL_0__1972_
timestamp 1701859473
transform 1 0 5670 0 1 4950
box -12 -8 32 272
use FILL  FILL_0__1973_
timestamp 1701859473
transform -1 0 6010 0 -1 3910
box -12 -8 32 272
use FILL  FILL_0__1974_
timestamp 1701859473
transform 1 0 6190 0 -1 3910
box -12 -8 32 272
use FILL  FILL_0__1975_
timestamp 1701859473
transform -1 0 5990 0 1 3910
box -12 -8 32 272
use FILL  FILL_0__1976_
timestamp 1701859473
transform -1 0 6450 0 -1 3910
box -12 -8 32 272
use FILL  FILL_0__1977_
timestamp 1701859473
transform 1 0 6770 0 1 2870
box -12 -8 32 272
use FILL  FILL_0__1978_
timestamp 1701859473
transform -1 0 6310 0 -1 2870
box -12 -8 32 272
use FILL  FILL_0__1979_
timestamp 1701859473
transform 1 0 6350 0 1 2870
box -12 -8 32 272
use FILL  FILL_0__1980_
timestamp 1701859473
transform 1 0 6550 0 1 2870
box -12 -8 32 272
use FILL  FILL_0__1981_
timestamp 1701859473
transform 1 0 6130 0 1 2870
box -12 -8 32 272
use FILL  FILL_0__1982_
timestamp 1701859473
transform -1 0 5590 0 -1 1830
box -12 -8 32 272
use FILL  FILL_0__1983_
timestamp 1701859473
transform -1 0 4690 0 -1 270
box -12 -8 32 272
use FILL  FILL_0__1984_
timestamp 1701859473
transform -1 0 6390 0 -1 1310
box -12 -8 32 272
use FILL  FILL_0__1985_
timestamp 1701859473
transform 1 0 4950 0 -1 1310
box -12 -8 32 272
use FILL  FILL_0__1986_
timestamp 1701859473
transform 1 0 8150 0 1 790
box -12 -8 32 272
use FILL  FILL_0__1987_
timestamp 1701859473
transform 1 0 6830 0 1 1310
box -12 -8 32 272
use FILL  FILL_0__1988_
timestamp 1701859473
transform -1 0 7290 0 1 1310
box -12 -8 32 272
use FILL  FILL_0__1989_
timestamp 1701859473
transform 1 0 2650 0 -1 5470
box -12 -8 32 272
use FILL  FILL_0__1990_
timestamp 1701859473
transform 1 0 1970 0 1 1830
box -12 -8 32 272
use FILL  FILL_0__1991_
timestamp 1701859473
transform -1 0 2690 0 1 1830
box -12 -8 32 272
use FILL  FILL_0__1992_
timestamp 1701859473
transform -1 0 4090 0 -1 2350
box -12 -8 32 272
use FILL  FILL_0__1993_
timestamp 1701859473
transform -1 0 4330 0 -1 2350
box -12 -8 32 272
use FILL  FILL_0__1994_
timestamp 1701859473
transform 1 0 2430 0 1 1830
box -12 -8 32 272
use FILL  FILL_0__1995_
timestamp 1701859473
transform 1 0 2910 0 1 1830
box -12 -8 32 272
use FILL  FILL_0__1996_
timestamp 1701859473
transform -1 0 6590 0 1 790
box -12 -8 32 272
use FILL  FILL_0__1997_
timestamp 1701859473
transform -1 0 4930 0 1 790
box -12 -8 32 272
use FILL  FILL_0__1998_
timestamp 1701859473
transform 1 0 4190 0 1 270
box -12 -8 32 272
use FILL  FILL_0__1999_
timestamp 1701859473
transform -1 0 3790 0 -1 270
box -12 -8 32 272
use FILL  FILL_0__2000_
timestamp 1701859473
transform -1 0 4470 0 -1 270
box -12 -8 32 272
use FILL  FILL_0__2001_
timestamp 1701859473
transform -1 0 5850 0 -1 2870
box -12 -8 32 272
use FILL  FILL_0__2002_
timestamp 1701859473
transform -1 0 1790 0 1 2870
box -12 -8 32 272
use FILL  FILL_0__2003_
timestamp 1701859473
transform 1 0 1290 0 -1 3390
box -12 -8 32 272
use FILL  FILL_0__2004_
timestamp 1701859473
transform 1 0 2710 0 -1 3390
box -12 -8 32 272
use FILL  FILL_0__2005_
timestamp 1701859473
transform -1 0 2990 0 1 2870
box -12 -8 32 272
use FILL  FILL_0__2006_
timestamp 1701859473
transform 1 0 2730 0 1 2870
box -12 -8 32 272
use FILL  FILL_0__2007_
timestamp 1701859473
transform 1 0 6750 0 -1 2870
box -12 -8 32 272
use FILL  FILL_0__2008_
timestamp 1701859473
transform 1 0 430 0 -1 1830
box -12 -8 32 272
use FILL  FILL_0__2009_
timestamp 1701859473
transform -1 0 3950 0 -1 3390
box -12 -8 32 272
use FILL  FILL_0__2010_
timestamp 1701859473
transform -1 0 4250 0 -1 2870
box -12 -8 32 272
use FILL  FILL_0__2011_
timestamp 1701859473
transform -1 0 1990 0 1 790
box -12 -8 32 272
use FILL  FILL_0__2012_
timestamp 1701859473
transform 1 0 1490 0 1 790
box -12 -8 32 272
use FILL  FILL_0__2013_
timestamp 1701859473
transform -1 0 1750 0 1 790
box -12 -8 32 272
use FILL  FILL_0__2014_
timestamp 1701859473
transform 1 0 4410 0 1 1310
box -12 -8 32 272
use FILL  FILL_0__2015_
timestamp 1701859473
transform 1 0 3130 0 1 1830
box -12 -8 32 272
use FILL  FILL_0__2016_
timestamp 1701859473
transform -1 0 3630 0 1 1830
box -12 -8 32 272
use FILL  FILL_0__2017_
timestamp 1701859473
transform -1 0 5150 0 -1 1830
box -12 -8 32 272
use FILL  FILL_0__2018_
timestamp 1701859473
transform 1 0 4910 0 -1 1830
box -12 -8 32 272
use FILL  FILL_0__2019_
timestamp 1701859473
transform -1 0 5430 0 -1 2870
box -12 -8 32 272
use FILL  FILL_0__2020_
timestamp 1701859473
transform -1 0 5190 0 -1 2870
box -12 -8 32 272
use FILL  FILL_0__2021_
timestamp 1701859473
transform -1 0 6830 0 -1 1310
box -12 -8 32 272
use FILL  FILL_0__2022_
timestamp 1701859473
transform -1 0 7070 0 1 790
box -12 -8 32 272
use FILL  FILL_0__2023_
timestamp 1701859473
transform 1 0 8110 0 1 1830
box -12 -8 32 272
use FILL  FILL_0__2024_
timestamp 1701859473
transform -1 0 8330 0 1 1830
box -12 -8 32 272
use FILL  FILL_0__2025_
timestamp 1701859473
transform 1 0 9490 0 -1 790
box -12 -8 32 272
use FILL  FILL_0__2026_
timestamp 1701859473
transform -1 0 8630 0 1 790
box -12 -8 32 272
use FILL  FILL_0__2027_
timestamp 1701859473
transform -1 0 6830 0 1 790
box -12 -8 32 272
use FILL  FILL_0__2028_
timestamp 1701859473
transform 1 0 6930 0 -1 790
box -12 -8 32 272
use FILL  FILL_0__2029_
timestamp 1701859473
transform 1 0 7370 0 1 270
box -12 -8 32 272
use FILL  FILL_0__2030_
timestamp 1701859473
transform -1 0 7050 0 -1 1310
box -12 -8 32 272
use FILL  FILL_0__2031_
timestamp 1701859473
transform 1 0 7370 0 -1 790
box -12 -8 32 272
use FILL  FILL_0__2032_
timestamp 1701859473
transform -1 0 8670 0 1 270
box -12 -8 32 272
use FILL  FILL_0__2033_
timestamp 1701859473
transform 1 0 8150 0 1 1310
box -12 -8 32 272
use FILL  FILL_0__2034_
timestamp 1701859473
transform -1 0 8830 0 -1 1310
box -12 -8 32 272
use FILL  FILL_0__2035_
timestamp 1701859473
transform -1 0 8410 0 1 790
box -12 -8 32 272
use FILL  FILL_0__2036_
timestamp 1701859473
transform -1 0 8570 0 -1 1830
box -12 -8 32 272
use FILL  FILL_0__2037_
timestamp 1701859473
transform -1 0 8630 0 -1 790
box -12 -8 32 272
use FILL  FILL_0__2038_
timestamp 1701859473
transform 1 0 7930 0 1 790
box -12 -8 32 272
use FILL  FILL_0__2039_
timestamp 1701859473
transform 1 0 7710 0 1 790
box -12 -8 32 272
use FILL  FILL_0__2040_
timestamp 1701859473
transform -1 0 7630 0 -1 790
box -12 -8 32 272
use FILL  FILL_0__2041_
timestamp 1701859473
transform -1 0 6850 0 -1 270
box -12 -8 32 272
use FILL  FILL_0__2042_
timestamp 1701859473
transform 1 0 8830 0 -1 790
box -12 -8 32 272
use FILL  FILL_0__2043_
timestamp 1701859473
transform 1 0 7150 0 1 270
box -12 -8 32 272
use FILL  FILL_0__2044_
timestamp 1701859473
transform 1 0 6890 0 1 270
box -12 -8 32 272
use FILL  FILL_0__2045_
timestamp 1701859473
transform -1 0 6210 0 1 270
box -12 -8 32 272
use FILL  FILL_0__2046_
timestamp 1701859473
transform 1 0 6390 0 -1 270
box -12 -8 32 272
use FILL  FILL_0__2047_
timestamp 1701859473
transform -1 0 6170 0 -1 270
box -12 -8 32 272
use FILL  FILL_0__2048_
timestamp 1701859473
transform -1 0 5970 0 -1 270
box -12 -8 32 272
use FILL  FILL_0__2049_
timestamp 1701859473
transform -1 0 7150 0 -1 790
box -12 -8 32 272
use FILL  FILL_0__2050_
timestamp 1701859473
transform 1 0 1390 0 -1 2870
box -12 -8 32 272
use FILL  FILL_0__2051_
timestamp 1701859473
transform 1 0 6190 0 -1 2350
box -12 -8 32 272
use FILL  FILL_0__2052_
timestamp 1701859473
transform -1 0 6090 0 1 790
box -12 -8 32 272
use FILL  FILL_0__2053_
timestamp 1701859473
transform -1 0 4310 0 1 1830
box -12 -8 32 272
use FILL  FILL_0__2054_
timestamp 1701859473
transform 1 0 2810 0 1 1310
box -12 -8 32 272
use FILL  FILL_0__2055_
timestamp 1701859473
transform -1 0 3070 0 1 1310
box -12 -8 32 272
use FILL  FILL_0__2056_
timestamp 1701859473
transform -1 0 1790 0 -1 1310
box -12 -8 32 272
use FILL  FILL_0__2057_
timestamp 1701859473
transform 1 0 2650 0 1 790
box -12 -8 32 272
use FILL  FILL_0__2058_
timestamp 1701859473
transform 1 0 3570 0 1 790
box -12 -8 32 272
use FILL  FILL_0__2059_
timestamp 1701859473
transform 1 0 3810 0 1 790
box -12 -8 32 272
use FILL  FILL_0__2060_
timestamp 1701859473
transform -1 0 4050 0 1 790
box -12 -8 32 272
use FILL  FILL_0__2061_
timestamp 1701859473
transform -1 0 2910 0 -1 270
box -12 -8 32 272
use FILL  FILL_0__2062_
timestamp 1701859473
transform 1 0 2690 0 1 270
box -12 -8 32 272
use FILL  FILL_0__2063_
timestamp 1701859473
transform 1 0 3070 0 -1 270
box -12 -8 32 272
use FILL  FILL_0__2064_
timestamp 1701859473
transform 1 0 3310 0 -1 270
box -12 -8 32 272
use FILL  FILL_0__2065_
timestamp 1701859473
transform -1 0 3550 0 -1 270
box -12 -8 32 272
use FILL  FILL_0__2066_
timestamp 1701859473
transform -1 0 5330 0 -1 270
box -12 -8 32 272
use FILL  FILL_0__2067_
timestamp 1701859473
transform 1 0 7270 0 1 790
box -12 -8 32 272
use FILL  FILL_0__2068_
timestamp 1701859473
transform 1 0 5830 0 1 790
box -12 -8 32 272
use FILL  FILL_0__2069_
timestamp 1701859473
transform 1 0 3310 0 -1 1830
box -12 -8 32 272
use FILL  FILL_0__2070_
timestamp 1701859473
transform -1 0 3790 0 -1 1830
box -12 -8 32 272
use FILL  FILL_0__2071_
timestamp 1701859473
transform -1 0 5630 0 1 790
box -12 -8 32 272
use FILL  FILL_0__2072_
timestamp 1701859473
transform -1 0 7690 0 1 1310
box -12 -8 32 272
use FILL  FILL_0__2073_
timestamp 1701859473
transform 1 0 6570 0 1 1310
box -12 -8 32 272
use FILL  FILL_0__2074_
timestamp 1701859473
transform 1 0 1710 0 1 1310
box -12 -8 32 272
use FILL  FILL_0__2075_
timestamp 1701859473
transform -1 0 2190 0 1 1310
box -12 -8 32 272
use FILL  FILL_0__2076_
timestamp 1701859473
transform -1 0 2230 0 -1 1310
box -12 -8 32 272
use FILL  FILL_0__2077_
timestamp 1701859473
transform 1 0 4090 0 -1 1310
box -12 -8 32 272
use FILL  FILL_0__2078_
timestamp 1701859473
transform -1 0 2230 0 1 1830
box -12 -8 32 272
use FILL  FILL_0__2079_
timestamp 1701859473
transform -1 0 870 0 -1 1830
box -12 -8 32 272
use FILL  FILL_0__2080_
timestamp 1701859473
transform 1 0 2190 0 -1 1830
box -12 -8 32 272
use FILL  FILL_0__2081_
timestamp 1701859473
transform 1 0 2430 0 -1 1830
box -12 -8 32 272
use FILL  FILL_0__2082_
timestamp 1701859473
transform -1 0 2650 0 -1 1830
box -12 -8 32 272
use FILL  FILL_0__2083_
timestamp 1701859473
transform 1 0 4330 0 -1 1310
box -12 -8 32 272
use FILL  FILL_0__2084_
timestamp 1701859473
transform -1 0 5170 0 1 790
box -12 -8 32 272
use FILL  FILL_0__2085_
timestamp 1701859473
transform -1 0 5010 0 -1 270
box -12 -8 32 272
use FILL  FILL_0__2086_
timestamp 1701859473
transform -1 0 4230 0 -1 270
box -12 -8 32 272
use FILL  FILL_0__2087_
timestamp 1701859473
transform -1 0 4710 0 1 790
box -12 -8 32 272
use FILL  FILL_0__2088_
timestamp 1701859473
transform -1 0 5550 0 1 270
box -12 -8 32 272
use FILL  FILL_0__2089_
timestamp 1701859473
transform 1 0 5310 0 1 270
box -12 -8 32 272
use FILL  FILL_0__2090_
timestamp 1701859473
transform -1 0 4890 0 -1 790
box -12 -8 32 272
use FILL  FILL_0__2091_
timestamp 1701859473
transform 1 0 3110 0 1 790
box -12 -8 32 272
use FILL  FILL_0__2092_
timestamp 1701859473
transform 1 0 2670 0 -1 270
box -12 -8 32 272
use FILL  FILL_0__2093_
timestamp 1701859473
transform -1 0 2830 0 -1 790
box -12 -8 32 272
use FILL  FILL_0__2094_
timestamp 1701859473
transform 1 0 2230 0 -1 270
box -12 -8 32 272
use FILL  FILL_0__2095_
timestamp 1701859473
transform 1 0 2430 0 -1 270
box -12 -8 32 272
use FILL  FILL_0__2096_
timestamp 1701859473
transform -1 0 4890 0 1 270
box -12 -8 32 272
use FILL  FILL_0__2097_
timestamp 1701859473
transform -1 0 5110 0 1 270
box -12 -8 32 272
use FILL  FILL_0__2098_
timestamp 1701859473
transform 1 0 4650 0 1 270
box -12 -8 32 272
use FILL  FILL_0__2099_
timestamp 1701859473
transform 1 0 3970 0 -1 270
box -12 -8 32 272
use FILL  FILL_0__2100_
timestamp 1701859473
transform -1 0 5830 0 -1 1830
box -12 -8 32 272
use FILL  FILL_0__2101_
timestamp 1701859473
transform -1 0 5750 0 1 1310
box -12 -8 32 272
use FILL  FILL_0__2102_
timestamp 1701859473
transform -1 0 6150 0 1 1310
box -12 -8 32 272
use FILL  FILL_0__2103_
timestamp 1701859473
transform 1 0 5710 0 -1 1310
box -12 -8 32 272
use FILL  FILL_0__2104_
timestamp 1701859473
transform -1 0 5950 0 1 1310
box -12 -8 32 272
use FILL  FILL_0__2105_
timestamp 1701859473
transform -1 0 4250 0 -1 1830
box -12 -8 32 272
use FILL  FILL_0__2106_
timestamp 1701859473
transform 1 0 3930 0 -1 790
box -12 -8 32 272
use FILL  FILL_0__2107_
timestamp 1701859473
transform -1 0 3510 0 -1 790
box -12 -8 32 272
use FILL  FILL_0__2108_
timestamp 1701859473
transform 1 0 2870 0 1 790
box -12 -8 32 272
use FILL  FILL_0__2109_
timestamp 1701859473
transform -1 0 3290 0 -1 790
box -12 -8 32 272
use FILL  FILL_0__2110_
timestamp 1701859473
transform 1 0 3050 0 -1 790
box -12 -8 32 272
use FILL  FILL_0__2111_
timestamp 1701859473
transform -1 0 3730 0 -1 790
box -12 -8 32 272
use FILL  FILL_0__2112_
timestamp 1701859473
transform -1 0 5090 0 -1 790
box -12 -8 32 272
use FILL  FILL_0__2113_
timestamp 1701859473
transform -1 0 5070 0 1 1310
box -12 -8 32 272
use FILL  FILL_0__2114_
timestamp 1701859473
transform -1 0 5510 0 1 1310
box -12 -8 32 272
use FILL  FILL_0__2115_
timestamp 1701859473
transform -1 0 5550 0 -1 790
box -12 -8 32 272
use FILL  FILL_0__2116_
timestamp 1701859473
transform 1 0 2370 0 1 1310
box -12 -8 32 272
use FILL  FILL_0__2117_
timestamp 1701859473
transform 1 0 2570 0 1 1310
box -12 -8 32 272
use FILL  FILL_0__2118_
timestamp 1701859473
transform 1 0 3750 0 1 1310
box -12 -8 32 272
use FILL  FILL_0__2119_
timestamp 1701859473
transform -1 0 4010 0 1 1310
box -12 -8 32 272
use FILL  FILL_0__2120_
timestamp 1701859473
transform 1 0 3870 0 -1 1310
box -12 -8 32 272
use FILL  FILL_0__2121_
timestamp 1701859473
transform -1 0 4450 0 1 270
box -12 -8 32 272
use FILL  FILL_0__2122_
timestamp 1701859473
transform -1 0 2790 0 1 2350
box -12 -8 32 272
use FILL  FILL_0__2123_
timestamp 1701859473
transform 1 0 2730 0 -1 2350
box -12 -8 32 272
use FILL  FILL_0__2124_
timestamp 1701859473
transform -1 0 3630 0 -1 2350
box -12 -8 32 272
use FILL  FILL_0__2125_
timestamp 1701859473
transform 1 0 5750 0 -1 3390
box -12 -8 32 272
use FILL  FILL_0__2126_
timestamp 1701859473
transform 1 0 5430 0 1 2870
box -12 -8 32 272
use FILL  FILL_0__2127_
timestamp 1701859473
transform -1 0 5910 0 1 2870
box -12 -8 32 272
use FILL  FILL_0__2128_
timestamp 1701859473
transform 1 0 4530 0 1 2870
box -12 -8 32 272
use FILL  FILL_0__2129_
timestamp 1701859473
transform 1 0 5210 0 1 2870
box -12 -8 32 272
use FILL  FILL_0__2130_
timestamp 1701859473
transform -1 0 4570 0 -1 2350
box -12 -8 32 272
use FILL  FILL_0__2131_
timestamp 1701859473
transform 1 0 4610 0 1 1310
box -12 -8 32 272
use FILL  FILL_0__2132_
timestamp 1701859473
transform -1 0 4490 0 1 790
box -12 -8 32 272
use FILL  FILL_0__2133_
timestamp 1701859473
transform 1 0 4410 0 -1 790
box -12 -8 32 272
use FILL  FILL_0__2134_
timestamp 1701859473
transform 1 0 3530 0 -1 2870
box -12 -8 32 272
use FILL  FILL_0__2135_
timestamp 1701859473
transform 1 0 4150 0 -1 3390
box -12 -8 32 272
use FILL  FILL_0__2136_
timestamp 1701859473
transform -1 0 2690 0 1 3390
box -12 -8 32 272
use FILL  FILL_0__2137_
timestamp 1701859473
transform 1 0 2250 0 1 3390
box -12 -8 32 272
use FILL  FILL_0__2138_
timestamp 1701859473
transform 1 0 3050 0 -1 4430
box -12 -8 32 272
use FILL  FILL_0__2139_
timestamp 1701859473
transform -1 0 2830 0 -1 4430
box -12 -8 32 272
use FILL  FILL_0__2140_
timestamp 1701859473
transform 1 0 2750 0 1 4430
box -12 -8 32 272
use FILL  FILL_0__2141_
timestamp 1701859473
transform -1 0 2990 0 1 4430
box -12 -8 32 272
use FILL  FILL_0__2142_
timestamp 1701859473
transform 1 0 2870 0 1 3390
box -12 -8 32 272
use FILL  FILL_0__2143_
timestamp 1701859473
transform -1 0 7370 0 -1 3390
box -12 -8 32 272
use FILL  FILL_0__2144_
timestamp 1701859473
transform 1 0 2010 0 1 2870
box -12 -8 32 272
use FILL  FILL_0__2145_
timestamp 1701859473
transform -1 0 9990 0 -1 2870
box -12 -8 32 272
use FILL  FILL_0__2146_
timestamp 1701859473
transform -1 0 7570 0 -1 3390
box -12 -8 32 272
use FILL  FILL_0__2147_
timestamp 1701859473
transform 1 0 7530 0 -1 3910
box -12 -8 32 272
use FILL  FILL_0__2148_
timestamp 1701859473
transform 1 0 7370 0 1 3390
box -12 -8 32 272
use FILL  FILL_0__2149_
timestamp 1701859473
transform 1 0 7570 0 1 3390
box -12 -8 32 272
use FILL  FILL_0__2150_
timestamp 1701859473
transform -1 0 7830 0 1 3390
box -12 -8 32 272
use FILL  FILL_0__2151_
timestamp 1701859473
transform 1 0 7110 0 -1 3390
box -12 -8 32 272
use FILL  FILL_0__2152_
timestamp 1701859473
transform 1 0 6870 0 -1 3390
box -12 -8 32 272
use FILL  FILL_0__2153_
timestamp 1701859473
transform -1 0 6010 0 -1 3390
box -12 -8 32 272
use FILL  FILL_0__2154_
timestamp 1701859473
transform 1 0 2770 0 -1 7030
box -12 -8 32 272
use FILL  FILL_0__2155_
timestamp 1701859473
transform 1 0 6330 0 1 5990
box -12 -8 32 272
use FILL  FILL_0__2156_
timestamp 1701859473
transform -1 0 4550 0 1 3910
box -12 -8 32 272
use FILL  FILL_0__2157_
timestamp 1701859473
transform -1 0 4690 0 -1 4430
box -12 -8 32 272
use FILL  FILL_0__2158_
timestamp 1701859473
transform -1 0 2550 0 1 2350
box -12 -8 32 272
use FILL  FILL_0__2159_
timestamp 1701859473
transform 1 0 3450 0 1 3910
box -12 -8 32 272
use FILL  FILL_0__2160_
timestamp 1701859473
transform -1 0 3770 0 -1 4430
box -12 -8 32 272
use FILL  FILL_0__2161_
timestamp 1701859473
transform -1 0 3910 0 1 3910
box -12 -8 32 272
use FILL  FILL_0__2162_
timestamp 1701859473
transform -1 0 4350 0 1 3910
box -12 -8 32 272
use FILL  FILL_0__2163_
timestamp 1701859473
transform 1 0 3670 0 -1 3910
box -12 -8 32 272
use FILL  FILL_0__2164_
timestamp 1701859473
transform -1 0 490 0 -1 4950
box -12 -8 32 272
use FILL  FILL_0__2165_
timestamp 1701859473
transform -1 0 3190 0 -1 3910
box -12 -8 32 272
use FILL  FILL_0__2166_
timestamp 1701859473
transform 1 0 3890 0 -1 3910
box -12 -8 32 272
use FILL  FILL_0__2167_
timestamp 1701859473
transform 1 0 4090 0 1 3910
box -12 -8 32 272
use FILL  FILL_0__2168_
timestamp 1701859473
transform 1 0 3010 0 1 3910
box -12 -8 32 272
use FILL  FILL_0__2169_
timestamp 1701859473
transform 1 0 2370 0 -1 4430
box -12 -8 32 272
use FILL  FILL_0__2170_
timestamp 1701859473
transform -1 0 2630 0 -1 4430
box -12 -8 32 272
use FILL  FILL_0__2171_
timestamp 1701859473
transform 1 0 3970 0 -1 4430
box -12 -8 32 272
use FILL  FILL_0__2172_
timestamp 1701859473
transform 1 0 4210 0 -1 4430
box -12 -8 32 272
use FILL  FILL_0__2173_
timestamp 1701859473
transform -1 0 4450 0 -1 4430
box -12 -8 32 272
use FILL  FILL_0__2174_
timestamp 1701859473
transform 1 0 5950 0 1 7030
box -12 -8 32 272
use FILL  FILL_0__2175_
timestamp 1701859473
transform -1 0 2450 0 1 8070
box -12 -8 32 272
use FILL  FILL_0__2176_
timestamp 1701859473
transform -1 0 6370 0 -1 8070
box -12 -8 32 272
use FILL  FILL_0__2177_
timestamp 1701859473
transform 1 0 4890 0 1 8070
box -12 -8 32 272
use FILL  FILL_0__2178_
timestamp 1701859473
transform -1 0 4070 0 -1 8590
box -12 -8 32 272
use FILL  FILL_0__2179_
timestamp 1701859473
transform -1 0 5890 0 -1 8070
box -12 -8 32 272
use FILL  FILL_0__2180_
timestamp 1701859473
transform -1 0 2910 0 -1 9630
box -12 -8 32 272
use FILL  FILL_0__2181_
timestamp 1701859473
transform 1 0 4970 0 1 7550
box -12 -8 32 272
use FILL  FILL_0__2182_
timestamp 1701859473
transform 1 0 5490 0 -1 10150
box -12 -8 32 272
use FILL  FILL_0__2183_
timestamp 1701859473
transform -1 0 3470 0 1 10150
box -12 -8 32 272
use FILL  FILL_0__2184_
timestamp 1701859473
transform 1 0 4290 0 1 8070
box -12 -8 32 272
use FILL  FILL_0__2185_
timestamp 1701859473
transform 1 0 5890 0 1 10150
box -12 -8 32 272
use FILL  FILL_0__2186_
timestamp 1701859473
transform 1 0 3450 0 1 10670
box -12 -8 32 272
use FILL  FILL_0__2187_
timestamp 1701859473
transform -1 0 5370 0 -1 10670
box -12 -8 32 272
use FILL  FILL_0__2188_
timestamp 1701859473
transform 1 0 2050 0 -1 10670
box -12 -8 32 272
use FILL  FILL_0__2189_
timestamp 1701859473
transform 1 0 5610 0 -1 10670
box -12 -8 32 272
use FILL  FILL_0__2190_
timestamp 1701859473
transform -1 0 2770 0 1 10150
box -12 -8 32 272
use FILL  FILL_0__2191_
timestamp 1701859473
transform -1 0 5250 0 -1 10150
box -12 -8 32 272
use FILL  FILL_0__2192_
timestamp 1701859473
transform -1 0 11050 0 1 3910
box -12 -8 32 272
use FILL  FILL_0__2193_
timestamp 1701859473
transform 1 0 1170 0 -1 3910
box -12 -8 32 272
use FILL  FILL_0__2194_
timestamp 1701859473
transform 1 0 970 0 -1 3910
box -12 -8 32 272
use FILL  FILL_0__2195_
timestamp 1701859473
transform 1 0 2550 0 1 3910
box -12 -8 32 272
use FILL  FILL_0__2196_
timestamp 1701859473
transform 1 0 2790 0 1 3910
box -12 -8 32 272
use FILL  FILL_0__2197_
timestamp 1701859473
transform 1 0 5270 0 1 3910
box -12 -8 32 272
use FILL  FILL_0__2198_
timestamp 1701859473
transform 1 0 210 0 1 1830
box -12 -8 32 272
use FILL  FILL_0__2199_
timestamp 1701859473
transform -1 0 2770 0 -1 3910
box -12 -8 32 272
use FILL  FILL_0__2200_
timestamp 1701859473
transform 1 0 5290 0 -1 3910
box -12 -8 32 272
use FILL  FILL_0__2201_
timestamp 1701859473
transform -1 0 5530 0 1 3910
box -12 -8 32 272
use FILL  FILL_0__2202_
timestamp 1701859473
transform -1 0 8110 0 -1 4430
box -12 -8 32 272
use FILL  FILL_0__2203_
timestamp 1701859473
transform -1 0 4830 0 -1 3910
box -12 -8 32 272
use FILL  FILL_0__2204_
timestamp 1701859473
transform 1 0 5050 0 -1 3910
box -12 -8 32 272
use FILL  FILL_0__2205_
timestamp 1701859473
transform -1 0 8910 0 -1 3910
box -12 -8 32 272
use FILL  FILL_0__2206_
timestamp 1701859473
transform 1 0 8990 0 1 3910
box -12 -8 32 272
use FILL  FILL_0__2207_
timestamp 1701859473
transform 1 0 9450 0 -1 3910
box -12 -8 32 272
use FILL  FILL_0__2208_
timestamp 1701859473
transform -1 0 9710 0 -1 3910
box -12 -8 32 272
use FILL  FILL_0__2209_
timestamp 1701859473
transform -1 0 9510 0 1 4430
box -12 -8 32 272
use FILL  FILL_0__2210_
timestamp 1701859473
transform -1 0 10510 0 -1 4950
box -12 -8 32 272
use FILL  FILL_0__2211_
timestamp 1701859473
transform 1 0 9210 0 -1 3910
box -12 -8 32 272
use FILL  FILL_0__2212_
timestamp 1701859473
transform -1 0 8790 0 1 3910
box -12 -8 32 272
use FILL  FILL_0__2213_
timestamp 1701859473
transform -1 0 9230 0 1 3910
box -12 -8 32 272
use FILL  FILL_0__2214_
timestamp 1701859473
transform -1 0 9430 0 -1 4430
box -12 -8 32 272
use FILL  FILL_0__2215_
timestamp 1701859473
transform 1 0 9630 0 -1 4430
box -12 -8 32 272
use FILL  FILL_0__2216_
timestamp 1701859473
transform -1 0 9390 0 -1 7030
box -12 -8 32 272
use FILL  FILL_0__2217_
timestamp 1701859473
transform 1 0 9170 0 -1 4430
box -12 -8 32 272
use FILL  FILL_0__2218_
timestamp 1701859473
transform -1 0 9690 0 1 3910
box -12 -8 32 272
use FILL  FILL_0__2219_
timestamp 1701859473
transform 1 0 9870 0 1 3910
box -12 -8 32 272
use FILL  FILL_0__2220_
timestamp 1701859473
transform 1 0 10250 0 -1 4950
box -12 -8 32 272
use FILL  FILL_0__2221_
timestamp 1701859473
transform -1 0 9630 0 -1 7030
box -12 -8 32 272
use FILL  FILL_0__2222_
timestamp 1701859473
transform 1 0 9990 0 1 4430
box -12 -8 32 272
use FILL  FILL_0__2223_
timestamp 1701859473
transform -1 0 9890 0 -1 4430
box -12 -8 32 272
use FILL  FILL_0__2224_
timestamp 1701859473
transform -1 0 9750 0 1 4430
box -12 -8 32 272
use FILL  FILL_0__2225_
timestamp 1701859473
transform 1 0 9990 0 -1 4950
box -12 -8 32 272
use FILL  FILL_0__2226_
timestamp 1701859473
transform 1 0 8870 0 -1 7030
box -12 -8 32 272
use FILL  FILL_0__2227_
timestamp 1701859473
transform -1 0 9150 0 -1 7030
box -12 -8 32 272
use FILL  FILL_0__2228_
timestamp 1701859473
transform -1 0 5690 0 -1 7030
box -12 -8 32 272
use FILL  FILL_0__2229_
timestamp 1701859473
transform 1 0 4250 0 1 3390
box -12 -8 32 272
use FILL  FILL_0__2230_
timestamp 1701859473
transform -1 0 4350 0 -1 3910
box -12 -8 32 272
use FILL  FILL_0__2231_
timestamp 1701859473
transform -1 0 4130 0 -1 3910
box -12 -8 32 272
use FILL  FILL_0__2232_
timestamp 1701859473
transform 1 0 1530 0 1 2870
box -12 -8 32 272
use FILL  FILL_0__2233_
timestamp 1701859473
transform 1 0 2250 0 1 2870
box -12 -8 32 272
use FILL  FILL_0__2234_
timestamp 1701859473
transform -1 0 2510 0 1 2870
box -12 -8 32 272
use FILL  FILL_0__2235_
timestamp 1701859473
transform 1 0 6270 0 1 3390
box -12 -8 32 272
use FILL  FILL_0__2236_
timestamp 1701859473
transform -1 0 5550 0 -1 3910
box -12 -8 32 272
use FILL  FILL_0__2237_
timestamp 1701859473
transform -1 0 4590 0 -1 3910
box -12 -8 32 272
use FILL  FILL_0__2238_
timestamp 1701859473
transform 1 0 4650 0 -1 4950
box -12 -8 32 272
use FILL  FILL_0__2239_
timestamp 1701859473
transform 1 0 2770 0 1 4950
box -12 -8 32 272
use FILL  FILL_0__2240_
timestamp 1701859473
transform 1 0 2330 0 1 3910
box -12 -8 32 272
use FILL  FILL_0__2241_
timestamp 1701859473
transform -1 0 2350 0 1 4950
box -12 -8 32 272
use FILL  FILL_0__2242_
timestamp 1701859473
transform 1 0 2390 0 -1 4950
box -12 -8 32 272
use FILL  FILL_0__2243_
timestamp 1701859473
transform 1 0 2570 0 1 4950
box -12 -8 32 272
use FILL  FILL_0__2244_
timestamp 1701859473
transform 1 0 2990 0 1 4950
box -12 -8 32 272
use FILL  FILL_0__2245_
timestamp 1701859473
transform 1 0 2830 0 1 5990
box -12 -8 32 272
use FILL  FILL_0__2246_
timestamp 1701859473
transform 1 0 2850 0 -1 4950
box -12 -8 32 272
use FILL  FILL_0__2247_
timestamp 1701859473
transform -1 0 2970 0 -1 6510
box -12 -8 32 272
use FILL  FILL_0__2248_
timestamp 1701859473
transform 1 0 3430 0 -1 7030
box -12 -8 32 272
use FILL  FILL_0__2249_
timestamp 1701859473
transform 1 0 6210 0 1 7030
box -12 -8 32 272
use FILL  FILL_0__2250_
timestamp 1701859473
transform -1 0 10510 0 -1 7550
box -12 -8 32 272
use FILL  FILL_0__2251_
timestamp 1701859473
transform -1 0 10570 0 1 8070
box -12 -8 32 272
use FILL  FILL_0__2252_
timestamp 1701859473
transform -1 0 10870 0 -1 8070
box -12 -8 32 272
use FILL  FILL_0__2253_
timestamp 1701859473
transform -1 0 10630 0 -1 8070
box -12 -8 32 272
use FILL  FILL_0__2254_
timestamp 1701859473
transform 1 0 5330 0 1 8070
box -12 -8 32 272
use FILL  FILL_0__2255_
timestamp 1701859473
transform 1 0 2950 0 1 7030
box -12 -8 32 272
use FILL  FILL_0__2256_
timestamp 1701859473
transform -1 0 5070 0 1 7030
box -12 -8 32 272
use FILL  FILL_0__2257_
timestamp 1701859473
transform 1 0 5010 0 -1 7550
box -12 -8 32 272
use FILL  FILL_0__2258_
timestamp 1701859473
transform 1 0 5650 0 -1 8590
box -12 -8 32 272
use FILL  FILL_0__2259_
timestamp 1701859473
transform 1 0 10270 0 -1 7550
box -12 -8 32 272
use FILL  FILL_0__2260_
timestamp 1701859473
transform 1 0 9850 0 1 8070
box -12 -8 32 272
use FILL  FILL_0__2261_
timestamp 1701859473
transform -1 0 10150 0 1 7550
box -12 -8 32 272
use FILL  FILL_0__2262_
timestamp 1701859473
transform -1 0 9910 0 1 7550
box -12 -8 32 272
use FILL  FILL_0__2263_
timestamp 1701859473
transform 1 0 5410 0 1 7550
box -12 -8 32 272
use FILL  FILL_0__2264_
timestamp 1701859473
transform 1 0 1570 0 -1 6510
box -12 -8 32 272
use FILL  FILL_0__2265_
timestamp 1701859473
transform 1 0 1750 0 -1 6510
box -12 -8 32 272
use FILL  FILL_0__2266_
timestamp 1701859473
transform 1 0 3850 0 1 6510
box -12 -8 32 272
use FILL  FILL_0__2267_
timestamp 1701859473
transform -1 0 3610 0 -1 7550
box -12 -8 32 272
use FILL  FILL_0__2268_
timestamp 1701859473
transform 1 0 4290 0 -1 7550
box -12 -8 32 272
use FILL  FILL_0__2269_
timestamp 1701859473
transform 1 0 5610 0 1 7550
box -12 -8 32 272
use FILL  FILL_0__2270_
timestamp 1701859473
transform 1 0 8530 0 1 7550
box -12 -8 32 272
use FILL  FILL_0__2271_
timestamp 1701859473
transform -1 0 8810 0 -1 8070
box -12 -8 32 272
use FILL  FILL_0__2272_
timestamp 1701859473
transform -1 0 9070 0 -1 8070
box -12 -8 32 272
use FILL  FILL_0__2273_
timestamp 1701859473
transform -1 0 8570 0 -1 8070
box -12 -8 32 272
use FILL  FILL_0__2274_
timestamp 1701859473
transform -1 0 5930 0 -1 9630
box -12 -8 32 272
use FILL  FILL_0__2275_
timestamp 1701859473
transform -1 0 2230 0 1 8070
box -12 -8 32 272
use FILL  FILL_0__2276_
timestamp 1701859473
transform -1 0 3110 0 1 8070
box -12 -8 32 272
use FILL  FILL_0__2277_
timestamp 1701859473
transform -1 0 3590 0 -1 8590
box -12 -8 32 272
use FILL  FILL_0__2278_
timestamp 1701859473
transform 1 0 6490 0 1 9110
box -12 -8 32 272
use FILL  FILL_0__2279_
timestamp 1701859473
transform -1 0 10190 0 1 5990
box -12 -8 32 272
use FILL  FILL_0__2280_
timestamp 1701859473
transform 1 0 10370 0 1 5990
box -12 -8 32 272
use FILL  FILL_0__2281_
timestamp 1701859473
transform -1 0 10650 0 -1 5990
box -12 -8 32 272
use FILL  FILL_0__2282_
timestamp 1701859473
transform -1 0 10430 0 -1 6510
box -12 -8 32 272
use FILL  FILL_0__2283_
timestamp 1701859473
transform 1 0 5890 0 -1 8590
box -12 -8 32 272
use FILL  FILL_0__2284_
timestamp 1701859473
transform -1 0 2010 0 1 8070
box -12 -8 32 272
use FILL  FILL_0__2285_
timestamp 1701859473
transform -1 0 4070 0 1 8070
box -12 -8 32 272
use FILL  FILL_0__2286_
timestamp 1701859473
transform 1 0 4970 0 -1 8590
box -12 -8 32 272
use FILL  FILL_0__2287_
timestamp 1701859473
transform -1 0 6050 0 1 8590
box -12 -8 32 272
use FILL  FILL_0__2288_
timestamp 1701859473
transform -1 0 8770 0 1 7550
box -12 -8 32 272
use FILL  FILL_0__2289_
timestamp 1701859473
transform 1 0 8430 0 1 8070
box -12 -8 32 272
use FILL  FILL_0__2290_
timestamp 1701859473
transform -1 0 9930 0 -1 8070
box -12 -8 32 272
use FILL  FILL_0__2291_
timestamp 1701859473
transform -1 0 8710 0 1 8070
box -12 -8 32 272
use FILL  FILL_0__2292_
timestamp 1701859473
transform -1 0 6150 0 -1 9110
box -12 -8 32 272
use FILL  FILL_0__2293_
timestamp 1701859473
transform -1 0 2470 0 -1 8590
box -12 -8 32 272
use FILL  FILL_0__2294_
timestamp 1701859473
transform -1 0 3950 0 1 8590
box -12 -8 32 272
use FILL  FILL_0__2295_
timestamp 1701859473
transform 1 0 4870 0 1 8590
box -12 -8 32 272
use FILL  FILL_0__2296_
timestamp 1701859473
transform 1 0 6590 0 -1 9110
box -12 -8 32 272
use FILL  FILL_0__2297_
timestamp 1701859473
transform -1 0 9490 0 -1 5990
box -12 -8 32 272
use FILL  FILL_0__2298_
timestamp 1701859473
transform -1 0 9930 0 -1 5470
box -12 -8 32 272
use FILL  FILL_0__2299_
timestamp 1701859473
transform -1 0 9270 0 -1 6510
box -12 -8 32 272
use FILL  FILL_0__2300_
timestamp 1701859473
transform 1 0 9470 0 1 5990
box -12 -8 32 272
use FILL  FILL_0__2301_
timestamp 1701859473
transform 1 0 5510 0 1 9630
box -12 -8 32 272
use FILL  FILL_0__2302_
timestamp 1701859473
transform -1 0 3410 0 -1 9110
box -12 -8 32 272
use FILL  FILL_0__2303_
timestamp 1701859473
transform 1 0 2530 0 1 9110
box -12 -8 32 272
use FILL  FILL_0__2304_
timestamp 1701859473
transform 1 0 2730 0 -1 9110
box -12 -8 32 272
use FILL  FILL_0__2305_
timestamp 1701859473
transform -1 0 3710 0 1 8590
box -12 -8 32 272
use FILL  FILL_0__2306_
timestamp 1701859473
transform 1 0 4390 0 1 8590
box -12 -8 32 272
use FILL  FILL_0__2307_
timestamp 1701859473
transform 1 0 6250 0 1 9110
box -12 -8 32 272
use FILL  FILL_0__2308_
timestamp 1701859473
transform -1 0 8830 0 -1 6510
box -12 -8 32 272
use FILL  FILL_0__2309_
timestamp 1701859473
transform -1 0 8530 0 1 5990
box -12 -8 32 272
use FILL  FILL_0__2310_
timestamp 1701859473
transform -1 0 9030 0 -1 6510
box -12 -8 32 272
use FILL  FILL_0__2311_
timestamp 1701859473
transform -1 0 8590 0 -1 6510
box -12 -8 32 272
use FILL  FILL_0__2312_
timestamp 1701859473
transform -1 0 5490 0 -1 9630
box -12 -8 32 272
use FILL  FILL_0__2313_
timestamp 1701859473
transform -1 0 1770 0 1 8590
box -12 -8 32 272
use FILL  FILL_0__2314_
timestamp 1701859473
transform 1 0 1370 0 -1 8590
box -12 -8 32 272
use FILL  FILL_0__2315_
timestamp 1701859473
transform 1 0 1810 0 -1 8590
box -12 -8 32 272
use FILL  FILL_0__2316_
timestamp 1701859473
transform -1 0 4170 0 1 8590
box -12 -8 32 272
use FILL  FILL_0__2317_
timestamp 1701859473
transform 1 0 4630 0 1 8590
box -12 -8 32 272
use FILL  FILL_0__2318_
timestamp 1701859473
transform 1 0 6730 0 1 9110
box -12 -8 32 272
use FILL  FILL_0__2319_
timestamp 1701859473
transform -1 0 11050 0 1 4430
box -12 -8 32 272
use FILL  FILL_0__2320_
timestamp 1701859473
transform 1 0 5030 0 1 3910
box -12 -8 32 272
use FILL  FILL_0__2321_
timestamp 1701859473
transform 1 0 6450 0 1 3910
box -12 -8 32 272
use FILL  FILL_0__2322_
timestamp 1701859473
transform -1 0 7830 0 1 3910
box -12 -8 32 272
use FILL  FILL_0__2323_
timestamp 1701859473
transform 1 0 7870 0 -1 4430
box -12 -8 32 272
use FILL  FILL_0__2324_
timestamp 1701859473
transform -1 0 11090 0 -1 2870
box -12 -8 32 272
use FILL  FILL_0__2325_
timestamp 1701859473
transform -1 0 8070 0 1 3910
box -12 -8 32 272
use FILL  FILL_0__2326_
timestamp 1701859473
transform -1 0 3110 0 -1 4950
box -12 -8 32 272
use FILL  FILL_0__2327_
timestamp 1701859473
transform -1 0 3310 0 -1 4950
box -12 -8 32 272
use FILL  FILL_0__2328_
timestamp 1701859473
transform 1 0 3790 0 -1 5470
box -12 -8 32 272
use FILL  FILL_0__2329_
timestamp 1701859473
transform 1 0 3550 0 -1 5470
box -12 -8 32 272
use FILL  FILL_0__2330_
timestamp 1701859473
transform 1 0 3690 0 1 4950
box -12 -8 32 272
use FILL  FILL_0__2331_
timestamp 1701859473
transform 1 0 4770 0 1 3910
box -12 -8 32 272
use FILL  FILL_0__2332_
timestamp 1701859473
transform -1 0 4110 0 1 4950
box -12 -8 32 272
use FILL  FILL_0__2333_
timestamp 1701859473
transform -1 0 11070 0 -1 4430
box -12 -8 32 272
use FILL  FILL_0__2334_
timestamp 1701859473
transform 1 0 8950 0 -1 4430
box -12 -8 32 272
use FILL  FILL_0__2335_
timestamp 1701859473
transform 1 0 5130 0 -1 5470
box -12 -8 32 272
use FILL  FILL_0__2336_
timestamp 1701859473
transform -1 0 4990 0 1 5990
box -12 -8 32 272
use FILL  FILL_0__2337_
timestamp 1701859473
transform 1 0 4490 0 1 3390
box -12 -8 32 272
use FILL  FILL_0__2338_
timestamp 1701859473
transform 1 0 3090 0 1 3390
box -12 -8 32 272
use FILL  FILL_0__2339_
timestamp 1701859473
transform 1 0 4670 0 1 3390
box -12 -8 32 272
use FILL  FILL_0__2340_
timestamp 1701859473
transform 1 0 4910 0 1 3390
box -12 -8 32 272
use FILL  FILL_0__2341_
timestamp 1701859473
transform -1 0 490 0 1 5990
box -12 -8 32 272
use FILL  FILL_0__2342_
timestamp 1701859473
transform 1 0 2590 0 1 5470
box -12 -8 32 272
use FILL  FILL_0__2343_
timestamp 1701859473
transform -1 0 4530 0 1 6510
box -12 -8 32 272
use FILL  FILL_0__2344_
timestamp 1701859473
transform -1 0 4810 0 1 5470
box -12 -8 32 272
use FILL  FILL_0__2345_
timestamp 1701859473
transform -1 0 4610 0 1 5470
box -12 -8 32 272
use FILL  FILL_0__2346_
timestamp 1701859473
transform -1 0 4770 0 -1 5990
box -12 -8 32 272
use FILL  FILL_0__2347_
timestamp 1701859473
transform -1 0 5630 0 -1 5990
box -12 -8 32 272
use FILL  FILL_0__2348_
timestamp 1701859473
transform 1 0 5190 0 -1 6510
box -12 -8 32 272
use FILL  FILL_0__2349_
timestamp 1701859473
transform -1 0 4970 0 -1 6510
box -12 -8 32 272
use FILL  FILL_0__2350_
timestamp 1701859473
transform -1 0 4390 0 -1 6510
box -12 -8 32 272
use FILL  FILL_0__2351_
timestamp 1701859473
transform 1 0 5530 0 1 7030
box -12 -8 32 272
use FILL  FILL_0__2352_
timestamp 1701859473
transform -1 0 5750 0 1 7030
box -12 -8 32 272
use FILL  FILL_0__2353_
timestamp 1701859473
transform -1 0 690 0 1 7030
box -12 -8 32 272
use FILL  FILL_0__2354_
timestamp 1701859473
transform 1 0 5390 0 -1 5990
box -12 -8 32 272
use FILL  FILL_0__2355_
timestamp 1701859473
transform 1 0 5290 0 1 7030
box -12 -8 32 272
use FILL  FILL_0__2356_
timestamp 1701859473
transform -1 0 4790 0 -1 7550
box -12 -8 32 272
use FILL  FILL_0__2357_
timestamp 1701859473
transform 1 0 4650 0 1 8070
box -12 -8 32 272
use FILL  FILL_0__2358_
timestamp 1701859473
transform 1 0 5130 0 1 8070
box -12 -8 32 272
use FILL  FILL_0__2359_
timestamp 1701859473
transform -1 0 5450 0 -1 8590
box -12 -8 32 272
use FILL  FILL_0__2360_
timestamp 1701859473
transform -1 0 690 0 -1 6510
box -12 -8 32 272
use FILL  FILL_0__2361_
timestamp 1701859473
transform -1 0 5190 0 1 5990
box -12 -8 32 272
use FILL  FILL_0__2362_
timestamp 1701859473
transform 1 0 5190 0 1 6510
box -12 -8 32 272
use FILL  FILL_0__2363_
timestamp 1701859473
transform 1 0 5210 0 -1 7030
box -12 -8 32 272
use FILL  FILL_0__2364_
timestamp 1701859473
transform 1 0 5210 0 -1 8070
box -12 -8 32 272
use FILL  FILL_0__2365_
timestamp 1701859473
transform 1 0 5450 0 -1 8070
box -12 -8 32 272
use FILL  FILL_0__2366_
timestamp 1701859473
transform -1 0 5670 0 -1 8070
box -12 -8 32 272
use FILL  FILL_0__2367_
timestamp 1701859473
transform 1 0 2630 0 -1 7550
box -12 -8 32 272
use FILL  FILL_0__2368_
timestamp 1701859473
transform -1 0 5470 0 -1 7030
box -12 -8 32 272
use FILL  FILL_0__2369_
timestamp 1701859473
transform 1 0 5170 0 1 7550
box -12 -8 32 272
use FILL  FILL_0__2370_
timestamp 1701859473
transform -1 0 5210 0 -1 8590
box -12 -8 32 272
use FILL  FILL_0__2371_
timestamp 1701859473
transform 1 0 5890 0 -1 9110
box -12 -8 32 272
use FILL  FILL_0__2372_
timestamp 1701859473
transform 1 0 6050 0 1 9110
box -12 -8 32 272
use FILL  FILL_0__2373_
timestamp 1701859473
transform -1 0 6130 0 -1 9630
box -12 -8 32 272
use FILL  FILL_0__2374_
timestamp 1701859473
transform 1 0 10 0 -1 9110
box -12 -8 32 272
use FILL  FILL_0__2375_
timestamp 1701859473
transform -1 0 4150 0 1 5470
box -12 -8 32 272
use FILL  FILL_0__2376_
timestamp 1701859473
transform 1 0 4490 0 -1 5990
box -12 -8 32 272
use FILL  FILL_0__2377_
timestamp 1701859473
transform -1 0 3910 0 -1 6510
box -12 -8 32 272
use FILL  FILL_0__2378_
timestamp 1701859473
transform 1 0 3650 0 -1 6510
box -12 -8 32 272
use FILL  FILL_0__2379_
timestamp 1701859473
transform -1 0 4970 0 1 6510
box -12 -8 32 272
use FILL  FILL_0__2380_
timestamp 1701859473
transform -1 0 4750 0 -1 8590
box -12 -8 32 272
use FILL  FILL_0__2381_
timestamp 1701859473
transform 1 0 3810 0 -1 8590
box -12 -8 32 272
use FILL  FILL_0__2382_
timestamp 1701859473
transform -1 0 4510 0 -1 8590
box -12 -8 32 272
use FILL  FILL_0__2383_
timestamp 1701859473
transform -1 0 5590 0 1 8590
box -12 -8 32 272
use FILL  FILL_0__2384_
timestamp 1701859473
transform -1 0 5810 0 1 8590
box -12 -8 32 272
use FILL  FILL_0__2385_
timestamp 1701859473
transform 1 0 1190 0 -1 10150
box -12 -8 32 272
use FILL  FILL_0__2386_
timestamp 1701859473
transform 1 0 5450 0 -1 7550
box -12 -8 32 272
use FILL  FILL_0__2387_
timestamp 1701859473
transform 1 0 5430 0 -1 9110
box -12 -8 32 272
use FILL  FILL_0__2388_
timestamp 1701859473
transform -1 0 5230 0 -1 9110
box -12 -8 32 272
use FILL  FILL_0__2389_
timestamp 1701859473
transform -1 0 5010 0 -1 9630
box -12 -8 32 272
use FILL  FILL_0__2390_
timestamp 1701859473
transform 1 0 5070 0 1 9630
box -12 -8 32 272
use FILL  FILL_0__2391_
timestamp 1701859473
transform -1 0 5290 0 1 9630
box -12 -8 32 272
use FILL  FILL_0__2392_
timestamp 1701859473
transform 1 0 1390 0 -1 10150
box -12 -8 32 272
use FILL  FILL_0__2393_
timestamp 1701859473
transform -1 0 5250 0 -1 7550
box -12 -8 32 272
use FILL  FILL_0__2394_
timestamp 1701859473
transform 1 0 5330 0 1 8590
box -12 -8 32 272
use FILL  FILL_0__2395_
timestamp 1701859473
transform -1 0 5690 0 -1 9110
box -12 -8 32 272
use FILL  FILL_0__2396_
timestamp 1701859473
transform 1 0 5610 0 1 9110
box -12 -8 32 272
use FILL  FILL_0__2397_
timestamp 1701859473
transform 1 0 5850 0 1 9110
box -12 -8 32 272
use FILL  FILL_0__2398_
timestamp 1701859473
transform 1 0 5670 0 -1 9630
box -12 -8 32 272
use FILL  FILL_0__2399_
timestamp 1701859473
transform -1 0 3110 0 -1 5470
box -12 -8 32 272
use FILL  FILL_0__2400_
timestamp 1701859473
transform -1 0 3290 0 1 5990
box -12 -8 32 272
use FILL  FILL_0__2401_
timestamp 1701859473
transform 1 0 3210 0 -1 6510
box -12 -8 32 272
use FILL  FILL_0__2402_
timestamp 1701859473
transform -1 0 2150 0 -1 4430
box -12 -8 32 272
use FILL  FILL_0__2403_
timestamp 1701859473
transform -1 0 2550 0 1 4430
box -12 -8 32 272
use FILL  FILL_0__2404_
timestamp 1701859473
transform -1 0 2870 0 -1 5470
box -12 -8 32 272
use FILL  FILL_0__2405_
timestamp 1701859473
transform 1 0 2250 0 -1 2870
box -12 -8 32 272
use FILL  FILL_0__2406_
timestamp 1701859473
transform 1 0 2950 0 -1 3390
box -12 -8 32 272
use FILL  FILL_0__2407_
timestamp 1701859473
transform -1 0 3090 0 1 5470
box -12 -8 32 272
use FILL  FILL_0__2408_
timestamp 1701859473
transform 1 0 710 0 -1 2870
box -12 -8 32 272
use FILL  FILL_0__2409_
timestamp 1701859473
transform 1 0 730 0 -1 3910
box -12 -8 32 272
use FILL  FILL_0__2410_
timestamp 1701859473
transform 1 0 1130 0 1 4430
box -12 -8 32 272
use FILL  FILL_0__2411_
timestamp 1701859473
transform -1 0 690 0 -1 4950
box -12 -8 32 272
use FILL  FILL_0__2412_
timestamp 1701859473
transform 1 0 2370 0 -1 5990
box -12 -8 32 272
use FILL  FILL_0__2413_
timestamp 1701859473
transform 1 0 2830 0 1 5470
box -12 -8 32 272
use FILL  FILL_0__2414_
timestamp 1701859473
transform 1 0 3990 0 -1 5470
box -12 -8 32 272
use FILL  FILL_0__2415_
timestamp 1701859473
transform -1 0 3930 0 1 7030
box -12 -8 32 272
use FILL  FILL_0__2416_
timestamp 1701859473
transform 1 0 3890 0 1 4950
box -12 -8 32 272
use FILL  FILL_0__2417_
timestamp 1701859473
transform 1 0 4230 0 -1 5470
box -12 -8 32 272
use FILL  FILL_0__2418_
timestamp 1701859473
transform -1 0 1490 0 -1 4950
box -12 -8 32 272
use FILL  FILL_0__2419_
timestamp 1701859473
transform 1 0 2070 0 1 4430
box -12 -8 32 272
use FILL  FILL_0__2420_
timestamp 1701859473
transform 1 0 3730 0 1 5990
box -12 -8 32 272
use FILL  FILL_0__2421_
timestamp 1701859473
transform -1 0 3510 0 1 5990
box -12 -8 32 272
use FILL  FILL_0__2422_
timestamp 1701859473
transform -1 0 3390 0 -1 5990
box -12 -8 32 272
use FILL  FILL_0__2423_
timestamp 1701859473
transform -1 0 3610 0 -1 5990
box -12 -8 32 272
use FILL  FILL_0__2424_
timestamp 1701859473
transform 1 0 3150 0 -1 5990
box -12 -8 32 272
use FILL  FILL_0__2425_
timestamp 1701859473
transform 1 0 4290 0 1 5990
box -12 -8 32 272
use FILL  FILL_0__2426_
timestamp 1701859473
transform 1 0 3890 0 -1 7030
box -12 -8 32 272
use FILL  FILL_0__2427_
timestamp 1701859473
transform 1 0 4710 0 1 5990
box -12 -8 32 272
use FILL  FILL_0__2428_
timestamp 1701859473
transform 1 0 4470 0 1 5990
box -12 -8 32 272
use FILL  FILL_0__2429_
timestamp 1701859473
transform -1 0 4150 0 -1 6510
box -12 -8 32 272
use FILL  FILL_0__2430_
timestamp 1701859473
transform 1 0 4710 0 1 6510
box -12 -8 32 272
use FILL  FILL_0__2431_
timestamp 1701859473
transform -1 0 4810 0 -1 7030
box -12 -8 32 272
use FILL  FILL_0__2432_
timestamp 1701859473
transform 1 0 5030 0 -1 7030
box -12 -8 32 272
use FILL  FILL_0__2433_
timestamp 1701859473
transform -1 0 4290 0 -1 8070
box -12 -8 32 272
use FILL  FILL_0__2434_
timestamp 1701859473
transform 1 0 4770 0 1 7550
box -12 -8 32 272
use FILL  FILL_0__2435_
timestamp 1701859473
transform 1 0 4110 0 1 7030
box -12 -8 32 272
use FILL  FILL_0__2436_
timestamp 1701859473
transform -1 0 4550 0 -1 7550
box -12 -8 32 272
use FILL  FILL_0__2437_
timestamp 1701859473
transform -1 0 4530 0 -1 8070
box -12 -8 32 272
use FILL  FILL_0__2438_
timestamp 1701859473
transform -1 0 4770 0 -1 8070
box -12 -8 32 272
use FILL  FILL_0__2439_
timestamp 1701859473
transform -1 0 5010 0 -1 8070
box -12 -8 32 272
use FILL  FILL_0__2440_
timestamp 1701859473
transform 1 0 4550 0 1 10150
box -12 -8 32 272
use FILL  FILL_0__2441_
timestamp 1701859473
transform 1 0 3830 0 -1 7550
box -12 -8 32 272
use FILL  FILL_0__2442_
timestamp 1701859473
transform -1 0 4050 0 -1 8070
box -12 -8 32 272
use FILL  FILL_0__2443_
timestamp 1701859473
transform -1 0 3830 0 1 8070
box -12 -8 32 272
use FILL  FILL_0__2444_
timestamp 1701859473
transform 1 0 3570 0 1 8070
box -12 -8 32 272
use FILL  FILL_0__2445_
timestamp 1701859473
transform -1 0 4550 0 1 7550
box -12 -8 32 272
use FILL  FILL_0__2446_
timestamp 1701859473
transform 1 0 4470 0 1 8070
box -12 -8 32 272
use FILL  FILL_0__2447_
timestamp 1701859473
transform 1 0 4210 0 1 9110
box -12 -8 32 272
use FILL  FILL_0__2448_
timestamp 1701859473
transform 1 0 4870 0 1 9110
box -12 -8 32 272
use FILL  FILL_0__2449_
timestamp 1701859473
transform 1 0 5130 0 1 9110
box -12 -8 32 272
use FILL  FILL_0__2450_
timestamp 1701859473
transform 1 0 5370 0 1 9110
box -12 -8 32 272
use FILL  FILL_0__2451_
timestamp 1701859473
transform -1 0 5250 0 -1 9630
box -12 -8 32 272
use FILL  FILL_0__2452_
timestamp 1701859473
transform -1 0 5170 0 -1 10670
box -12 -8 32 272
use FILL  FILL_0__2453_
timestamp 1701859473
transform 1 0 3710 0 -1 10150
box -12 -8 32 272
use FILL  FILL_0__2454_
timestamp 1701859473
transform 1 0 3830 0 1 7550
box -12 -8 32 272
use FILL  FILL_0__2455_
timestamp 1701859473
transform 1 0 3790 0 -1 8070
box -12 -8 32 272
use FILL  FILL_0__2456_
timestamp 1701859473
transform -1 0 3570 0 -1 8070
box -12 -8 32 272
use FILL  FILL_0__2457_
timestamp 1701859473
transform 1 0 3330 0 1 8070
box -12 -8 32 272
use FILL  FILL_0__2458_
timestamp 1701859473
transform -1 0 4270 0 -1 8590
box -12 -8 32 272
use FILL  FILL_0__2459_
timestamp 1701859473
transform -1 0 4430 0 -1 11190
box -12 -8 32 272
use FILL  FILL_0__2460_
timestamp 1701859473
transform 1 0 4070 0 -1 10670
box -12 -8 32 272
use FILL  FILL_0__2461_
timestamp 1701859473
transform 1 0 4250 0 -1 9110
box -12 -8 32 272
use FILL  FILL_0__2462_
timestamp 1701859473
transform -1 0 4510 0 -1 9110
box -12 -8 32 272
use FILL  FILL_0__2463_
timestamp 1701859473
transform -1 0 4750 0 -1 9110
box -12 -8 32 272
use FILL  FILL_0__2464_
timestamp 1701859473
transform -1 0 4990 0 -1 9110
box -12 -8 32 272
use FILL  FILL_0__2465_
timestamp 1701859473
transform -1 0 4850 0 -1 11190
box -12 -8 32 272
use FILL  FILL_0__2466_
timestamp 1701859473
transform -1 0 3930 0 -1 10150
box -12 -8 32 272
use FILL  FILL_0__2467_
timestamp 1701859473
transform -1 0 4030 0 -1 9630
box -12 -8 32 272
use FILL  FILL_0__2468_
timestamp 1701859473
transform -1 0 4290 0 -1 9630
box -12 -8 32 272
use FILL  FILL_0__2469_
timestamp 1701859473
transform -1 0 4150 0 1 9630
box -12 -8 32 272
use FILL  FILL_0__2470_
timestamp 1701859473
transform -1 0 4390 0 1 9630
box -12 -8 32 272
use FILL  FILL_0__2471_
timestamp 1701859473
transform -1 0 4970 0 -1 10670
box -12 -8 32 272
use FILL  FILL_0__2472_
timestamp 1701859473
transform 1 0 3930 0 1 9630
box -12 -8 32 272
use FILL  FILL_0__2473_
timestamp 1701859473
transform 1 0 4490 0 -1 9630
box -12 -8 32 272
use FILL  FILL_0__2474_
timestamp 1701859473
transform -1 0 4770 0 -1 9630
box -12 -8 32 272
use FILL  FILL_0__2475_
timestamp 1701859473
transform 1 0 4610 0 1 9630
box -12 -8 32 272
use FILL  FILL_0__2476_
timestamp 1701859473
transform -1 0 4850 0 1 9630
box -12 -8 32 272
use FILL  FILL_0__2477_
timestamp 1701859473
transform 1 0 4790 0 1 10670
box -12 -8 32 272
use FILL  FILL_0__2478_
timestamp 1701859473
transform 1 0 3030 0 1 5990
box -12 -8 32 272
use FILL  FILL_0__2479_
timestamp 1701859473
transform -1 0 2590 0 1 5990
box -12 -8 32 272
use FILL  FILL_0__2480_
timestamp 1701859473
transform -1 0 2610 0 -1 5990
box -12 -8 32 272
use FILL  FILL_0__2481_
timestamp 1701859473
transform -1 0 2850 0 -1 5990
box -12 -8 32 272
use FILL  FILL_0__2482_
timestamp 1701859473
transform 1 0 1430 0 -1 5990
box -12 -8 32 272
use FILL  FILL_0__2483_
timestamp 1701859473
transform 1 0 2250 0 1 6510
box -12 -8 32 272
use FILL  FILL_0__2484_
timestamp 1701859473
transform -1 0 1870 0 1 6510
box -12 -8 32 272
use FILL  FILL_0__2485_
timestamp 1701859473
transform -1 0 2070 0 1 6510
box -12 -8 32 272
use FILL  FILL_0__2486_
timestamp 1701859473
transform 1 0 2270 0 -1 7030
box -12 -8 32 272
use FILL  FILL_0__2487_
timestamp 1701859473
transform 1 0 2030 0 -1 7030
box -12 -8 32 272
use FILL  FILL_0__2488_
timestamp 1701859473
transform -1 0 1830 0 -1 7030
box -12 -8 32 272
use FILL  FILL_0__2489_
timestamp 1701859473
transform 1 0 1330 0 -1 7030
box -12 -8 32 272
use FILL  FILL_0__2490_
timestamp 1701859473
transform -1 0 930 0 1 5470
box -12 -8 32 272
use FILL  FILL_0__2491_
timestamp 1701859473
transform 1 0 1130 0 1 5470
box -12 -8 32 272
use FILL  FILL_0__2492_
timestamp 1701859473
transform -1 0 1990 0 -1 6510
box -12 -8 32 272
use FILL  FILL_0__2493_
timestamp 1701859473
transform 1 0 1870 0 1 5990
box -12 -8 32 272
use FILL  FILL_0__2494_
timestamp 1701859473
transform -1 0 1430 0 1 5990
box -12 -8 32 272
use FILL  FILL_0__2495_
timestamp 1701859473
transform 1 0 1170 0 1 5990
box -12 -8 32 272
use FILL  FILL_0__2496_
timestamp 1701859473
transform 1 0 1570 0 -1 7030
box -12 -8 32 272
use FILL  FILL_0__2497_
timestamp 1701859473
transform -1 0 1770 0 -1 7550
box -12 -8 32 272
use FILL  FILL_0__2498_
timestamp 1701859473
transform 1 0 710 0 1 8070
box -12 -8 32 272
use FILL  FILL_0__2499_
timestamp 1701859473
transform 1 0 2390 0 1 7550
box -12 -8 32 272
use FILL  FILL_0__2500_
timestamp 1701859473
transform 1 0 1810 0 1 7550
box -12 -8 32 272
use FILL  FILL_0__2501_
timestamp 1701859473
transform 1 0 1590 0 1 7550
box -12 -8 32 272
use FILL  FILL_0__2502_
timestamp 1701859473
transform -1 0 1130 0 1 7550
box -12 -8 32 272
use FILL  FILL_0__2503_
timestamp 1701859473
transform -1 0 1370 0 1 8070
box -12 -8 32 272
use FILL  FILL_0__2504_
timestamp 1701859473
transform -1 0 1790 0 1 8070
box -12 -8 32 272
use FILL  FILL_0__2505_
timestamp 1701859473
transform 1 0 1130 0 1 8070
box -12 -8 32 272
use FILL  FILL_0__2506_
timestamp 1701859473
transform -1 0 1650 0 -1 8070
box -12 -8 32 272
use FILL  FILL_0__2507_
timestamp 1701859473
transform 1 0 1390 0 -1 8070
box -12 -8 32 272
use FILL  FILL_0__2508_
timestamp 1701859473
transform 1 0 910 0 1 8070
box -12 -8 32 272
use FILL  FILL_0__2509_
timestamp 1701859473
transform 1 0 470 0 -1 8590
box -12 -8 32 272
use FILL  FILL_0__2510_
timestamp 1701859473
transform -1 0 1410 0 1 9110
box -12 -8 32 272
use FILL  FILL_0__2511_
timestamp 1701859473
transform -1 0 1350 0 -1 9630
box -12 -8 32 272
use FILL  FILL_0__2512_
timestamp 1701859473
transform 1 0 910 0 -1 9630
box -12 -8 32 272
use FILL  FILL_0__2513_
timestamp 1701859473
transform -1 0 910 0 1 8590
box -12 -8 32 272
use FILL  FILL_0__2514_
timestamp 1701859473
transform 1 0 1990 0 -1 8590
box -12 -8 32 272
use FILL  FILL_0__2515_
timestamp 1701859473
transform 1 0 1110 0 -1 9110
box -12 -8 32 272
use FILL  FILL_0__2516_
timestamp 1701859473
transform -1 0 950 0 1 9110
box -12 -8 32 272
use FILL  FILL_0__2517_
timestamp 1701859473
transform -1 0 710 0 1 9110
box -12 -8 32 272
use FILL  FILL_0__2518_
timestamp 1701859473
transform 1 0 1570 0 -1 9630
box -12 -8 32 272
use FILL  FILL_0__2519_
timestamp 1701859473
transform 1 0 1670 0 1 9630
box -12 -8 32 272
use FILL  FILL_0__2520_
timestamp 1701859473
transform -1 0 2510 0 -1 9110
box -12 -8 32 272
use FILL  FILL_0__2521_
timestamp 1701859473
transform 1 0 2250 0 -1 9110
box -12 -8 32 272
use FILL  FILL_0__2522_
timestamp 1701859473
transform -1 0 1870 0 1 9630
box -12 -8 32 272
use FILL  FILL_0__2523_
timestamp 1701859473
transform -1 0 2090 0 1 9630
box -12 -8 32 272
use FILL  FILL_0__2524_
timestamp 1701859473
transform -1 0 1830 0 -1 9110
box -12 -8 32 272
use FILL  FILL_0__2525_
timestamp 1701859473
transform 1 0 710 0 -1 8590
box -12 -8 32 272
use FILL  FILL_0__2526_
timestamp 1701859473
transform -1 0 1610 0 -1 8590
box -12 -8 32 272
use FILL  FILL_0__2527_
timestamp 1701859473
transform -1 0 1150 0 -1 8590
box -12 -8 32 272
use FILL  FILL_0__2528_
timestamp 1701859473
transform -1 0 930 0 -1 8590
box -12 -8 32 272
use FILL  FILL_0__2529_
timestamp 1701859473
transform -1 0 1170 0 1 9110
box -12 -8 32 272
use FILL  FILL_0__2530_
timestamp 1701859473
transform -1 0 7430 0 -1 6510
box -12 -8 32 272
use FILL  FILL_0__2531_
timestamp 1701859473
transform 1 0 7850 0 1 7550
box -12 -8 32 272
use FILL  FILL_0__2532_
timestamp 1701859473
transform -1 0 9750 0 1 2870
box -12 -8 32 272
use FILL  FILL_0__2533_
timestamp 1701859473
transform -1 0 8830 0 1 4430
box -12 -8 32 272
use FILL  FILL_0__2534_
timestamp 1701859473
transform -1 0 9230 0 -1 5470
box -12 -8 32 272
use FILL  FILL_0__2535_
timestamp 1701859473
transform 1 0 10 0 -1 4950
box -12 -8 32 272
use FILL  FILL_0__2536_
timestamp 1701859473
transform 1 0 570 0 1 4950
box -12 -8 32 272
use FILL  FILL_0__2537_
timestamp 1701859473
transform 1 0 710 0 1 3390
box -12 -8 32 272
use FILL  FILL_0__2538_
timestamp 1701859473
transform -1 0 270 0 -1 3910
box -12 -8 32 272
use FILL  FILL_0__2539_
timestamp 1701859473
transform -1 0 30 0 1 4950
box -12 -8 32 272
use FILL  FILL_0__2540_
timestamp 1701859473
transform 1 0 2970 0 1 2350
box -12 -8 32 272
use FILL  FILL_0__2541_
timestamp 1701859473
transform -1 0 3230 0 1 2870
box -12 -8 32 272
use FILL  FILL_0__2542_
timestamp 1701859473
transform -1 0 2230 0 -1 6510
box -12 -8 32 272
use FILL  FILL_0__2543_
timestamp 1701859473
transform 1 0 790 0 1 4950
box -12 -8 32 272
use FILL  FILL_0__2544_
timestamp 1701859473
transform 1 0 1350 0 1 4430
box -12 -8 32 272
use FILL  FILL_0__2545_
timestamp 1701859473
transform 1 0 1210 0 -1 5470
box -12 -8 32 272
use FILL  FILL_0__2546_
timestamp 1701859473
transform -1 0 1950 0 -1 5470
box -12 -8 32 272
use FILL  FILL_0__2547_
timestamp 1701859473
transform 1 0 1890 0 -1 4430
box -12 -8 32 272
use FILL  FILL_0__2548_
timestamp 1701859473
transform 1 0 1010 0 1 4950
box -12 -8 32 272
use FILL  FILL_0__2549_
timestamp 1701859473
transform 1 0 1230 0 1 4950
box -12 -8 32 272
use FILL  FILL_0__2550_
timestamp 1701859473
transform -1 0 1710 0 -1 5470
box -12 -8 32 272
use FILL  FILL_0__2551_
timestamp 1701859473
transform 1 0 2490 0 -1 9630
box -12 -8 32 272
use FILL  FILL_0__2552_
timestamp 1701859473
transform 1 0 3330 0 -1 5470
box -12 -8 32 272
use FILL  FILL_0__2553_
timestamp 1701859473
transform -1 0 2710 0 -1 6510
box -12 -8 32 272
use FILL  FILL_0__2554_
timestamp 1701859473
transform -1 0 3170 0 1 6510
box -12 -8 32 272
use FILL  FILL_0__2555_
timestamp 1701859473
transform -1 0 3410 0 1 6510
box -12 -8 32 272
use FILL  FILL_0__2556_
timestamp 1701859473
transform -1 0 2730 0 1 6510
box -12 -8 32 272
use FILL  FILL_0__2557_
timestamp 1701859473
transform 1 0 2430 0 -1 6510
box -12 -8 32 272
use FILL  FILL_0__2558_
timestamp 1701859473
transform 1 0 3170 0 -1 7550
box -12 -8 32 272
use FILL  FILL_0__2559_
timestamp 1701859473
transform 1 0 3370 0 -1 7550
box -12 -8 32 272
use FILL  FILL_0__2560_
timestamp 1701859473
transform -1 0 3430 0 1 7030
box -12 -8 32 272
use FILL  FILL_0__2561_
timestamp 1701859473
transform -1 0 1450 0 1 4950
box -12 -8 32 272
use FILL  FILL_0__2562_
timestamp 1701859473
transform 1 0 3170 0 1 7030
box -12 -8 32 272
use FILL  FILL_0__2563_
timestamp 1701859473
transform 1 0 3730 0 1 5470
box -12 -8 32 272
use FILL  FILL_0__2564_
timestamp 1701859473
transform -1 0 3610 0 1 6510
box -12 -8 32 272
use FILL  FILL_0__2565_
timestamp 1701859473
transform 1 0 3670 0 1 7030
box -12 -8 32 272
use FILL  FILL_0__2566_
timestamp 1701859473
transform 1 0 3130 0 1 7550
box -12 -8 32 272
use FILL  FILL_0__2567_
timestamp 1701859473
transform 1 0 3090 0 -1 8070
box -12 -8 32 272
use FILL  FILL_0__2568_
timestamp 1701859473
transform -1 0 2910 0 -1 8590
box -12 -8 32 272
use FILL  FILL_0__2569_
timestamp 1701859473
transform 1 0 2670 0 -1 8590
box -12 -8 32 272
use FILL  FILL_0__2570_
timestamp 1701859473
transform 1 0 2850 0 -1 8070
box -12 -8 32 272
use FILL  FILL_0__2571_
timestamp 1701859473
transform -1 0 3810 0 -1 9630
box -12 -8 32 272
use FILL  FILL_0__2572_
timestamp 1701859473
transform -1 0 3830 0 -1 5990
box -12 -8 32 272
use FILL  FILL_0__2573_
timestamp 1701859473
transform -1 0 3690 0 -1 7030
box -12 -8 32 272
use FILL  FILL_0__2574_
timestamp 1701859473
transform 1 0 3410 0 -1 6510
box -12 -8 32 272
use FILL  FILL_0__2575_
timestamp 1701859473
transform 1 0 3310 0 -1 8070
box -12 -8 32 272
use FILL  FILL_0__2576_
timestamp 1701859473
transform -1 0 3350 0 -1 8590
box -12 -8 32 272
use FILL  FILL_0__2577_
timestamp 1701859473
transform 1 0 3230 0 1 9110
box -12 -8 32 272
use FILL  FILL_0__2578_
timestamp 1701859473
transform 1 0 3730 0 1 9110
box -12 -8 32 272
use FILL  FILL_0__2579_
timestamp 1701859473
transform -1 0 2710 0 -1 9630
box -12 -8 32 272
use FILL  FILL_0__2580_
timestamp 1701859473
transform -1 0 4070 0 -1 9110
box -12 -8 32 272
use FILL  FILL_0__2581_
timestamp 1701859473
transform -1 0 3990 0 1 9110
box -12 -8 32 272
use FILL  FILL_0__2582_
timestamp 1701859473
transform 1 0 3490 0 1 9110
box -12 -8 32 272
use FILL  FILL_0__2583_
timestamp 1701859473
transform 1 0 2990 0 1 9110
box -12 -8 32 272
use FILL  FILL_0__2584_
timestamp 1701859473
transform 1 0 2750 0 1 9110
box -12 -8 32 272
use FILL  FILL_0__2585_
timestamp 1701859473
transform 1 0 3850 0 -1 9110
box -12 -8 32 272
use FILL  FILL_0__2586_
timestamp 1701859473
transform 1 0 3010 0 1 9630
box -12 -8 32 272
use FILL  FILL_0__2587_
timestamp 1701859473
transform 1 0 3590 0 -1 9110
box -12 -8 32 272
use FILL  FILL_0__2588_
timestamp 1701859473
transform 1 0 3190 0 1 8590
box -12 -8 32 272
use FILL  FILL_0__2589_
timestamp 1701859473
transform 1 0 3030 0 -1 10150
box -12 -8 32 272
use FILL  FILL_0__2590_
timestamp 1701859473
transform 1 0 2770 0 -1 10150
box -12 -8 32 272
use FILL  FILL_0__2591_
timestamp 1701859473
transform -1 0 3530 0 -1 11190
box -12 -8 32 272
use FILL  FILL_0__2592_
timestamp 1701859473
transform -1 0 3590 0 -1 9630
box -12 -8 32 272
use FILL  FILL_0__2593_
timestamp 1701859473
transform -1 0 3110 0 -1 9630
box -12 -8 32 272
use FILL  FILL_0__2594_
timestamp 1701859473
transform -1 0 3270 0 -1 10150
box -12 -8 32 272
use FILL  FILL_0__2595_
timestamp 1701859473
transform 1 0 2990 0 -1 11190
box -12 -8 32 272
use FILL  FILL_0__2596_
timestamp 1701859473
transform 1 0 3270 0 -1 11190
box -12 -8 32 272
use FILL  FILL_0__2597_
timestamp 1701859473
transform 1 0 2730 0 -1 10670
box -12 -8 32 272
use FILL  FILL_0__2598_
timestamp 1701859473
transform -1 0 3470 0 1 9630
box -12 -8 32 272
use FILL  FILL_0__2599_
timestamp 1701859473
transform -1 0 3250 0 1 9630
box -12 -8 32 272
use FILL  FILL_0__2600_
timestamp 1701859473
transform -1 0 2970 0 1 10150
box -12 -8 32 272
use FILL  FILL_0__2601_
timestamp 1701859473
transform 1 0 2930 0 -1 10670
box -12 -8 32 272
use FILL  FILL_0__2602_
timestamp 1701859473
transform -1 0 3190 0 -1 10670
box -12 -8 32 272
use FILL  FILL_0__2603_
timestamp 1701859473
transform 1 0 3390 0 -1 10670
box -12 -8 32 272
use FILL  FILL_0__2604_
timestamp 1701859473
transform 1 0 3190 0 1 10150
box -12 -8 32 272
use FILL  FILL_0__2605_
timestamp 1701859473
transform 1 0 2310 0 1 10670
box -12 -8 32 272
use FILL  FILL_0__2606_
timestamp 1701859473
transform 1 0 2510 0 1 10670
box -12 -8 32 272
use FILL  FILL_0__2607_
timestamp 1701859473
transform -1 0 2750 0 1 10670
box -12 -8 32 272
use FILL  FILL_0__2608_
timestamp 1701859473
transform -1 0 3710 0 1 9630
box -12 -8 32 272
use FILL  FILL_0__2609_
timestamp 1701859473
transform -1 0 2330 0 1 9630
box -12 -8 32 272
use FILL  FILL_0__2610_
timestamp 1701859473
transform -1 0 2550 0 -1 10150
box -12 -8 32 272
use FILL  FILL_0__2611_
timestamp 1701859473
transform -1 0 2270 0 -1 10670
box -12 -8 32 272
use FILL  FILL_0__2612_
timestamp 1701859473
transform 1 0 2490 0 -1 10670
box -12 -8 32 272
use FILL  FILL_0__2613_
timestamp 1701859473
transform 1 0 1810 0 1 10670
box -12 -8 32 272
use FILL  FILL_0__2614_
timestamp 1701859473
transform 1 0 1810 0 -1 10670
box -12 -8 32 272
use FILL  FILL_0__2615_
timestamp 1701859473
transform -1 0 2330 0 -1 11190
box -12 -8 32 272
use FILL  FILL_0__2616_
timestamp 1701859473
transform -1 0 3350 0 -1 9630
box -12 -8 32 272
use FILL  FILL_0__2617_
timestamp 1701859473
transform 1 0 2250 0 -1 9630
box -12 -8 32 272
use FILL  FILL_0__2618_
timestamp 1701859473
transform -1 0 2530 0 1 10150
box -12 -8 32 272
use FILL  FILL_0__2619_
timestamp 1701859473
transform 1 0 2030 0 1 10670
box -12 -8 32 272
use FILL  FILL_0__2620_
timestamp 1701859473
transform 1 0 2070 0 -1 11190
box -12 -8 32 272
use FILL  FILL_0__2621_
timestamp 1701859473
transform -1 0 1350 0 1 5470
box -12 -8 32 272
use FILL  FILL_0__2622_
timestamp 1701859473
transform -1 0 1190 0 -1 5990
box -12 -8 32 272
use FILL  FILL_0__2623_
timestamp 1701859473
transform 1 0 2410 0 -1 5470
box -12 -8 32 272
use FILL  FILL_0__2624_
timestamp 1701859473
transform -1 0 2370 0 1 5470
box -12 -8 32 272
use FILL  FILL_0__2625_
timestamp 1701859473
transform 1 0 2170 0 -1 5470
box -12 -8 32 272
use FILL  FILL_0__2626_
timestamp 1701859473
transform -1 0 910 0 -1 5470
box -12 -8 32 272
use FILL  FILL_0__2627_
timestamp 1701859473
transform -1 0 1430 0 1 3910
box -12 -8 32 272
use FILL  FILL_0__2628_
timestamp 1701859473
transform 1 0 1110 0 1 3910
box -12 -8 32 272
use FILL  FILL_0__2629_
timestamp 1701859473
transform -1 0 710 0 -1 5470
box -12 -8 32 272
use FILL  FILL_0__2630_
timestamp 1701859473
transform 1 0 690 0 -1 5990
box -12 -8 32 272
use FILL  FILL_0__2631_
timestamp 1701859473
transform -1 0 690 0 1 5990
box -12 -8 32 272
use FILL  FILL_0__2632_
timestamp 1701859473
transform 1 0 2070 0 1 10150
box -12 -8 32 272
use FILL  FILL_0__2633_
timestamp 1701859473
transform -1 0 2310 0 1 10150
box -12 -8 32 272
use FILL  FILL_0__2634_
timestamp 1701859473
transform 1 0 2270 0 -1 10150
box -12 -8 32 272
use FILL  FILL_0__2635_
timestamp 1701859473
transform 1 0 2050 0 -1 10150
box -12 -8 32 272
use FILL  FILL_0__2636_
timestamp 1701859473
transform -1 0 690 0 -1 10150
box -12 -8 32 272
use FILL  FILL_0__2637_
timestamp 1701859473
transform -1 0 490 0 1 6510
box -12 -8 32 272
use FILL  FILL_0__2638_
timestamp 1701859473
transform -1 0 270 0 1 6510
box -12 -8 32 272
use FILL  FILL_0__2639_
timestamp 1701859473
transform -1 0 250 0 -1 6510
box -12 -8 32 272
use FILL  FILL_0__2640_
timestamp 1701859473
transform -1 0 250 0 1 5990
box -12 -8 32 272
use FILL  FILL_0__2641_
timestamp 1701859473
transform 1 0 10 0 -1 7550
box -12 -8 32 272
use FILL  FILL_0__2642_
timestamp 1701859473
transform -1 0 350 0 1 4950
box -12 -8 32 272
use FILL  FILL_0__2643_
timestamp 1701859473
transform -1 0 2490 0 1 6510
box -12 -8 32 272
use FILL  FILL_0__2644_
timestamp 1701859473
transform 1 0 2530 0 -1 7030
box -12 -8 32 272
use FILL  FILL_0__2645_
timestamp 1701859473
transform 1 0 2710 0 1 7030
box -12 -8 32 272
use FILL  FILL_0__2646_
timestamp 1701859473
transform 1 0 2010 0 1 7030
box -12 -8 32 272
use FILL  FILL_0__2647_
timestamp 1701859473
transform 1 0 690 0 1 7550
box -12 -8 32 272
use FILL  FILL_0__2648_
timestamp 1701859473
transform 1 0 230 0 1 7550
box -12 -8 32 272
use FILL  FILL_0__2649_
timestamp 1701859473
transform 1 0 210 0 -1 7550
box -12 -8 32 272
use FILL  FILL_0__2650_
timestamp 1701859473
transform -1 0 690 0 -1 7550
box -12 -8 32 272
use FILL  FILL_0__2651_
timestamp 1701859473
transform 1 0 430 0 -1 7550
box -12 -8 32 272
use FILL  FILL_0__2652_
timestamp 1701859473
transform 1 0 430 0 1 7030
box -12 -8 32 272
use FILL  FILL_0__2653_
timestamp 1701859473
transform 1 0 10 0 1 7550
box -12 -8 32 272
use FILL  FILL_0__2654_
timestamp 1701859473
transform -1 0 490 0 1 7550
box -12 -8 32 272
use FILL  FILL_0__2655_
timestamp 1701859473
transform 1 0 1810 0 1 7030
box -12 -8 32 272
use FILL  FILL_0__2656_
timestamp 1701859473
transform 1 0 1450 0 -1 5470
box -12 -8 32 272
use FILL  FILL_0__2657_
timestamp 1701859473
transform -1 0 1650 0 1 5990
box -12 -8 32 272
use FILL  FILL_0__2658_
timestamp 1701859473
transform -1 0 2130 0 1 5470
box -12 -8 32 272
use FILL  FILL_0__2659_
timestamp 1701859473
transform 1 0 1890 0 -1 5990
box -12 -8 32 272
use FILL  FILL_0__2660_
timestamp 1701859473
transform -1 0 1890 0 1 5470
box -12 -8 32 272
use FILL  FILL_0__2661_
timestamp 1701859473
transform -1 0 1570 0 1 5470
box -12 -8 32 272
use FILL  FILL_0__2662_
timestamp 1701859473
transform 1 0 670 0 1 5470
box -12 -8 32 272
use FILL  FILL_0__2663_
timestamp 1701859473
transform -1 0 950 0 -1 5990
box -12 -8 32 272
use FILL  FILL_0__2664_
timestamp 1701859473
transform 1 0 670 0 -1 7030
box -12 -8 32 272
use FILL  FILL_0__2665_
timestamp 1701859473
transform 1 0 1130 0 -1 7030
box -12 -8 32 272
use FILL  FILL_0__2666_
timestamp 1701859473
transform 1 0 1330 0 1 7030
box -12 -8 32 272
use FILL  FILL_0__2667_
timestamp 1701859473
transform 1 0 870 0 -1 7030
box -12 -8 32 272
use FILL  FILL_0__2668_
timestamp 1701859473
transform -1 0 2670 0 1 7550
box -12 -8 32 272
use FILL  FILL_0__2669_
timestamp 1701859473
transform 1 0 2610 0 -1 8070
box -12 -8 32 272
use FILL  FILL_0__2670_
timestamp 1701859473
transform 1 0 1870 0 -1 8070
box -12 -8 32 272
use FILL  FILL_0__2671_
timestamp 1701859473
transform -1 0 1370 0 1 7550
box -12 -8 32 272
use FILL  FILL_0__2672_
timestamp 1701859473
transform 1 0 1090 0 -1 7550
box -12 -8 32 272
use FILL  FILL_0__2673_
timestamp 1701859473
transform -1 0 1290 0 -1 7550
box -12 -8 32 272
use FILL  FILL_0__2674_
timestamp 1701859473
transform 1 0 1570 0 1 7030
box -12 -8 32 272
use FILL  FILL_0__2675_
timestamp 1701859473
transform 1 0 1510 0 -1 7550
box -12 -8 32 272
use FILL  FILL_0__2676_
timestamp 1701859473
transform -1 0 1950 0 -1 7550
box -12 -8 32 272
use FILL  FILL_0__2677_
timestamp 1701859473
transform 1 0 2350 0 -1 8070
box -12 -8 32 272
use FILL  FILL_0__2678_
timestamp 1701859473
transform -1 0 2130 0 -1 8070
box -12 -8 32 272
use FILL  FILL_0__2679_
timestamp 1701859473
transform -1 0 1570 0 1 8070
box -12 -8 32 272
use FILL  FILL_0__2680_
timestamp 1701859473
transform -1 0 250 0 -1 8590
box -12 -8 32 272
use FILL  FILL_0__2681_
timestamp 1701859473
transform 1 0 870 0 -1 7550
box -12 -8 32 272
use FILL  FILL_0__2682_
timestamp 1701859473
transform -1 0 250 0 -1 8070
box -12 -8 32 272
use FILL  FILL_0__2683_
timestamp 1701859473
transform -1 0 30 0 -1 9630
box -12 -8 32 272
use FILL  FILL_0__2684_
timestamp 1701859473
transform -1 0 30 0 1 10150
box -12 -8 32 272
use FILL  FILL_0__2685_
timestamp 1701859473
transform 1 0 910 0 1 5990
box -12 -8 32 272
use FILL  FILL_0__2686_
timestamp 1701859473
transform 1 0 890 0 1 7550
box -12 -8 32 272
use FILL  FILL_0__2687_
timestamp 1701859473
transform -1 0 890 0 -1 10150
box -12 -8 32 272
use FILL  FILL_0__2688_
timestamp 1701859473
transform 1 0 10 0 -1 10150
box -12 -8 32 272
use FILL  FILL_0__2689_
timestamp 1701859473
transform 1 0 230 0 -1 9630
box -12 -8 32 272
use FILL  FILL_0__2690_
timestamp 1701859473
transform 1 0 230 0 1 9110
box -12 -8 32 272
use FILL  FILL_0__2691_
timestamp 1701859473
transform 1 0 2690 0 1 8590
box -12 -8 32 272
use FILL  FILL_0__2692_
timestamp 1701859473
transform 1 0 2450 0 1 8590
box -12 -8 32 272
use FILL  FILL_0__2693_
timestamp 1701859473
transform -1 0 1110 0 -1 9630
box -12 -8 32 272
use FILL  FILL_0__2694_
timestamp 1701859473
transform 1 0 690 0 -1 9630
box -12 -8 32 272
use FILL  FILL_0__2695_
timestamp 1701859473
transform 1 0 10 0 1 9630
box -12 -8 32 272
use FILL  FILL_0__2696_
timestamp 1701859473
transform -1 0 490 0 -1 10150
box -12 -8 32 272
use FILL  FILL_0__2697_
timestamp 1701859473
transform 1 0 230 0 -1 10150
box -12 -8 32 272
use FILL  FILL_0__2698_
timestamp 1701859473
transform 1 0 250 0 1 9630
box -12 -8 32 272
use FILL  FILL_0__2699_
timestamp 1701859473
transform 1 0 470 0 -1 9630
box -12 -8 32 272
use FILL  FILL_0__2700_
timestamp 1701859473
transform 1 0 490 0 1 9630
box -12 -8 32 272
use FILL  FILL_0__2701_
timestamp 1701859473
transform -1 0 710 0 -1 10670
box -12 -8 32 272
use FILL  FILL_0__2702_
timestamp 1701859473
transform 1 0 3430 0 1 8590
box -12 -8 32 272
use FILL  FILL_0__2703_
timestamp 1701859473
transform -1 0 2970 0 1 8590
box -12 -8 32 272
use FILL  FILL_0__2704_
timestamp 1701859473
transform -1 0 1450 0 1 9630
box -12 -8 32 272
use FILL  FILL_0__2705_
timestamp 1701859473
transform 1 0 1190 0 1 9630
box -12 -8 32 272
use FILL  FILL_0__2706_
timestamp 1701859473
transform 1 0 210 0 1 10150
box -12 -8 32 272
use FILL  FILL_0__2707_
timestamp 1701859473
transform -1 0 450 0 1 10150
box -12 -8 32 272
use FILL  FILL_0__2708_
timestamp 1701859473
transform 1 0 650 0 1 10150
box -12 -8 32 272
use FILL  FILL_0__2709_
timestamp 1701859473
transform -1 0 470 0 -1 10670
box -12 -8 32 272
use FILL  FILL_0__2710_
timestamp 1701859473
transform 1 0 1650 0 1 10150
box -12 -8 32 272
use FILL  FILL_0__2711_
timestamp 1701859473
transform 1 0 2190 0 1 8590
box -12 -8 32 272
use FILL  FILL_0__2712_
timestamp 1701859473
transform -1 0 1970 0 1 8590
box -12 -8 32 272
use FILL  FILL_0__2713_
timestamp 1701859473
transform -1 0 1830 0 -1 9630
box -12 -8 32 272
use FILL  FILL_0__2714_
timestamp 1701859473
transform 1 0 1590 0 -1 10150
box -12 -8 32 272
use FILL  FILL_0__2715_
timestamp 1701859473
transform 1 0 910 0 1 10150
box -12 -8 32 272
use FILL  FILL_0__2716_
timestamp 1701859473
transform 1 0 1150 0 1 10150
box -12 -8 32 272
use FILL  FILL_0__2717_
timestamp 1701859473
transform 1 0 1410 0 1 10150
box -12 -8 32 272
use FILL  FILL_0__2718_
timestamp 1701859473
transform -1 0 9990 0 1 4950
box -12 -8 32 272
use FILL  FILL_0__2719_
timestamp 1701859473
transform -1 0 9750 0 1 4950
box -12 -8 32 272
use FILL  FILL_0__2720_
timestamp 1701859473
transform -1 0 4530 0 1 4950
box -12 -8 32 272
use FILL  FILL_0__2721_
timestamp 1701859473
transform -1 0 7290 0 -1 2350
box -12 -8 32 272
use FILL  FILL_0__2722_
timestamp 1701859473
transform 1 0 9930 0 -1 790
box -12 -8 32 272
use FILL  FILL_0__2723_
timestamp 1701859473
transform -1 0 7050 0 1 1830
box -12 -8 32 272
use FILL  FILL_0__2724_
timestamp 1701859473
transform -1 0 7050 0 -1 2350
box -12 -8 32 272
use FILL  FILL_0__2725_
timestamp 1701859473
transform 1 0 6910 0 1 3390
box -12 -8 32 272
use FILL  FILL_0__2726_
timestamp 1701859473
transform -1 0 7150 0 1 3390
box -12 -8 32 272
use FILL  FILL_0__2727_
timestamp 1701859473
transform -1 0 5370 0 1 3390
box -12 -8 32 272
use FILL  FILL_0__2728_
timestamp 1701859473
transform -1 0 5590 0 1 3390
box -12 -8 32 272
use FILL  FILL_0__2729_
timestamp 1701859473
transform -1 0 6690 0 -1 3910
box -12 -8 32 272
use FILL  FILL_0__2730_
timestamp 1701859473
transform 1 0 8190 0 -1 3910
box -12 -8 32 272
use FILL  FILL_0__2731_
timestamp 1701859473
transform 1 0 9210 0 1 1830
box -12 -8 32 272
use FILL  FILL_0__2732_
timestamp 1701859473
transform 1 0 7650 0 1 1830
box -12 -8 32 272
use FILL  FILL_0__2733_
timestamp 1701859473
transform 1 0 8530 0 1 2350
box -12 -8 32 272
use FILL  FILL_0__2734_
timestamp 1701859473
transform 1 0 7110 0 -1 5470
box -12 -8 32 272
use FILL  FILL_0__2735_
timestamp 1701859473
transform 1 0 7190 0 -1 2870
box -12 -8 32 272
use FILL  FILL_0__2736_
timestamp 1701859473
transform -1 0 7470 0 1 1310
box -12 -8 32 272
use FILL  FILL_0__2737_
timestamp 1701859473
transform 1 0 8530 0 1 1830
box -12 -8 32 272
use FILL  FILL_0__2738_
timestamp 1701859473
transform -1 0 7910 0 -1 2870
box -12 -8 32 272
use FILL  FILL_0__2739_
timestamp 1701859473
transform -1 0 7730 0 1 2870
box -12 -8 32 272
use FILL  FILL_0__2740_
timestamp 1701859473
transform -1 0 6510 0 -1 1830
box -12 -8 32 272
use FILL  FILL_0__2741_
timestamp 1701859473
transform 1 0 6710 0 -1 1830
box -12 -8 32 272
use FILL  FILL_0__2742_
timestamp 1701859473
transform -1 0 8150 0 -1 2870
box -12 -8 32 272
use FILL  FILL_0__2743_
timestamp 1701859473
transform -1 0 8170 0 1 2870
box -12 -8 32 272
use FILL  FILL_0__2744_
timestamp 1701859473
transform -1 0 7290 0 -1 270
box -12 -8 32 272
use FILL  FILL_0__2745_
timestamp 1701859473
transform -1 0 7250 0 1 1830
box -12 -8 32 272
use FILL  FILL_0__2746_
timestamp 1701859473
transform 1 0 7910 0 1 2870
box -12 -8 32 272
use FILL  FILL_0__2747_
timestamp 1701859473
transform -1 0 7710 0 -1 2350
box -12 -8 32 272
use FILL  FILL_0__2748_
timestamp 1701859473
transform 1 0 7890 0 -1 2350
box -12 -8 32 272
use FILL  FILL_0__2749_
timestamp 1701859473
transform 1 0 5850 0 1 1830
box -12 -8 32 272
use FILL  FILL_0__2750_
timestamp 1701859473
transform -1 0 6610 0 -1 1310
box -12 -8 32 272
use FILL  FILL_0__2751_
timestamp 1701859473
transform -1 0 6330 0 1 1830
box -12 -8 32 272
use FILL  FILL_0__2752_
timestamp 1701859473
transform -1 0 7690 0 1 2350
box -12 -8 32 272
use FILL  FILL_0__2753_
timestamp 1701859473
transform -1 0 7430 0 1 2350
box -12 -8 32 272
use FILL  FILL_0__2754_
timestamp 1701859473
transform 1 0 8770 0 -1 4950
box -12 -8 32 272
use FILL  FILL_0__2755_
timestamp 1701859473
transform 1 0 9670 0 1 790
box -12 -8 32 272
use FILL  FILL_0__2756_
timestamp 1701859473
transform -1 0 9910 0 1 790
box -12 -8 32 272
use FILL  FILL_0__2757_
timestamp 1701859473
transform 1 0 10610 0 -1 2870
box -12 -8 32 272
use FILL  FILL_0__2758_
timestamp 1701859473
transform -1 0 9110 0 -1 2870
box -12 -8 32 272
use FILL  FILL_0__2759_
timestamp 1701859473
transform 1 0 9030 0 1 4430
box -12 -8 32 272
use FILL  FILL_0__2760_
timestamp 1701859473
transform 1 0 10370 0 -1 790
box -12 -8 32 272
use FILL  FILL_0__2761_
timestamp 1701859473
transform 1 0 10130 0 -1 790
box -12 -8 32 272
use FILL  FILL_0__2762_
timestamp 1701859473
transform -1 0 10810 0 -1 1830
box -12 -8 32 272
use FILL  FILL_0__2763_
timestamp 1701859473
transform 1 0 6550 0 1 1830
box -12 -8 32 272
use FILL  FILL_0__2764_
timestamp 1701859473
transform -1 0 6810 0 1 1830
box -12 -8 32 272
use FILL  FILL_0__2765_
timestamp 1701859473
transform -1 0 10110 0 1 1830
box -12 -8 32 272
use FILL  FILL_0__2766_
timestamp 1701859473
transform -1 0 9930 0 -1 1830
box -12 -8 32 272
use FILL  FILL_0__2767_
timestamp 1701859473
transform -1 0 10350 0 -1 1830
box -12 -8 32 272
use FILL  FILL_0__2768_
timestamp 1701859473
transform -1 0 10330 0 1 1830
box -12 -8 32 272
use FILL  FILL_0__2769_
timestamp 1701859473
transform -1 0 10790 0 1 2350
box -12 -8 32 272
use FILL  FILL_0__2770_
timestamp 1701859473
transform -1 0 10570 0 -1 1830
box -12 -8 32 272
use FILL  FILL_0__2771_
timestamp 1701859473
transform 1 0 10990 0 1 2350
box -12 -8 32 272
use FILL  FILL_0__2772_
timestamp 1701859473
transform -1 0 10650 0 1 4950
box -12 -8 32 272
use FILL  FILL_0__2773_
timestamp 1701859473
transform 1 0 10390 0 -1 3910
box -12 -8 32 272
use FILL  FILL_0__2774_
timestamp 1701859473
transform -1 0 10690 0 -1 2350
box -12 -8 32 272
use FILL  FILL_0__2775_
timestamp 1701859473
transform -1 0 9050 0 -1 1310
box -12 -8 32 272
use FILL  FILL_0__2776_
timestamp 1701859473
transform 1 0 10590 0 -1 790
box -12 -8 32 272
use FILL  FILL_0__2777_
timestamp 1701859473
transform -1 0 8350 0 -1 270
box -12 -8 32 272
use FILL  FILL_0__2778_
timestamp 1701859473
transform 1 0 10890 0 1 270
box -12 -8 32 272
use FILL  FILL_0__2779_
timestamp 1701859473
transform 1 0 8970 0 -1 1830
box -12 -8 32 272
use FILL  FILL_0__2780_
timestamp 1701859473
transform -1 0 9990 0 1 1310
box -12 -8 32 272
use FILL  FILL_0__2781_
timestamp 1701859473
transform 1 0 10130 0 -1 1310
box -12 -8 32 272
use FILL  FILL_0__2782_
timestamp 1701859473
transform 1 0 8750 0 1 1830
box -12 -8 32 272
use FILL  FILL_0__2783_
timestamp 1701859473
transform 1 0 8310 0 -1 1310
box -12 -8 32 272
use FILL  FILL_0__2784_
timestamp 1701859473
transform 1 0 8550 0 -1 1310
box -12 -8 32 272
use FILL  FILL_0__2785_
timestamp 1701859473
transform 1 0 8770 0 -1 1830
box -12 -8 32 272
use FILL  FILL_0__2786_
timestamp 1701859473
transform -1 0 9250 0 -1 1310
box -12 -8 32 272
use FILL  FILL_0__2787_
timestamp 1701859473
transform -1 0 9450 0 -1 1830
box -12 -8 32 272
use FILL  FILL_0__2788_
timestamp 1701859473
transform 1 0 10130 0 -1 1830
box -12 -8 32 272
use FILL  FILL_0__2789_
timestamp 1701859473
transform 1 0 10210 0 1 1310
box -12 -8 32 272
use FILL  FILL_0__2790_
timestamp 1701859473
transform -1 0 10010 0 -1 2350
box -12 -8 32 272
use FILL  FILL_0__2791_
timestamp 1701859473
transform 1 0 9770 0 -1 2350
box -12 -8 32 272
use FILL  FILL_0__2792_
timestamp 1701859473
transform -1 0 10230 0 -1 2350
box -12 -8 32 272
use FILL  FILL_0__2793_
timestamp 1701859473
transform -1 0 10470 0 -1 2350
box -12 -8 32 272
use FILL  FILL_0__2794_
timestamp 1701859473
transform -1 0 10890 0 -1 2350
box -12 -8 32 272
use FILL  FILL_0__2795_
timestamp 1701859473
transform -1 0 10850 0 -1 2870
box -12 -8 32 272
use FILL  FILL_0__2796_
timestamp 1701859473
transform -1 0 10190 0 -1 2870
box -12 -8 32 272
use FILL  FILL_0__2797_
timestamp 1701859473
transform -1 0 9690 0 -1 1830
box -12 -8 32 272
use FILL  FILL_0__2798_
timestamp 1701859473
transform -1 0 10570 0 1 2350
box -12 -8 32 272
use FILL  FILL_0__2799_
timestamp 1701859473
transform 1 0 10350 0 -1 2870
box -12 -8 32 272
use FILL  FILL_0__2800_
timestamp 1701859473
transform -1 0 10370 0 -1 4430
box -12 -8 32 272
use FILL  FILL_0__2801_
timestamp 1701859473
transform -1 0 9330 0 -1 2870
box -12 -8 32 272
use FILL  FILL_0__2802_
timestamp 1701859473
transform -1 0 7190 0 -1 1830
box -12 -8 32 272
use FILL  FILL_0__2803_
timestamp 1701859473
transform 1 0 8390 0 -1 2870
box -12 -8 32 272
use FILL  FILL_0__2804_
timestamp 1701859473
transform -1 0 9450 0 -1 3390
box -12 -8 32 272
use FILL  FILL_0__2805_
timestamp 1701859473
transform -1 0 9750 0 -1 2870
box -12 -8 32 272
use FILL  FILL_0__2806_
timestamp 1701859473
transform 1 0 9510 0 -1 2870
box -12 -8 32 272
use FILL  FILL_0__2807_
timestamp 1701859473
transform 1 0 8850 0 -1 2350
box -12 -8 32 272
use FILL  FILL_0__2808_
timestamp 1701859473
transform 1 0 8610 0 -1 2350
box -12 -8 32 272
use FILL  FILL_0__2809_
timestamp 1701859473
transform 1 0 10330 0 1 2350
box -12 -8 32 272
use FILL  FILL_0__2810_
timestamp 1701859473
transform -1 0 10110 0 1 2350
box -12 -8 32 272
use FILL  FILL_0__2811_
timestamp 1701859473
transform 1 0 4890 0 -1 4430
box -12 -8 32 272
use FILL  FILL_0__2812_
timestamp 1701859473
transform -1 0 8850 0 1 4950
box -12 -8 32 272
use FILL  FILL_0__2813_
timestamp 1701859473
transform 1 0 8950 0 1 3390
box -12 -8 32 272
use FILL  FILL_0__2814_
timestamp 1701859473
transform -1 0 8770 0 -1 4430
box -12 -8 32 272
use FILL  FILL_0__2815_
timestamp 1701859473
transform -1 0 8550 0 1 3910
box -12 -8 32 272
use FILL  FILL_0__2816_
timestamp 1701859473
transform -1 0 8170 0 1 4950
box -12 -8 32 272
use FILL  FILL_0__2817_
timestamp 1701859473
transform 1 0 8610 0 1 4950
box -12 -8 32 272
use FILL  FILL_0__2818_
timestamp 1701859473
transform 1 0 8310 0 -1 4430
box -12 -8 32 272
use FILL  FILL_0__2819_
timestamp 1701859473
transform 1 0 8510 0 -1 4430
box -12 -8 32 272
use FILL  FILL_0__2820_
timestamp 1701859473
transform -1 0 9470 0 1 2350
box -12 -8 32 272
use FILL  FILL_0__2821_
timestamp 1701859473
transform 1 0 8990 0 1 2350
box -12 -8 32 272
use FILL  FILL_0__2822_
timestamp 1701859473
transform -1 0 8990 0 1 1830
box -12 -8 32 272
use FILL  FILL_0__2823_
timestamp 1701859473
transform -1 0 8770 0 1 2350
box -12 -8 32 272
use FILL  FILL_0__2824_
timestamp 1701859473
transform 1 0 9890 0 -1 3390
box -12 -8 32 272
use FILL  FILL_0__2825_
timestamp 1701859473
transform -1 0 10610 0 -1 3390
box -12 -8 32 272
use FILL  FILL_0__2826_
timestamp 1701859473
transform 1 0 9470 0 1 790
box -12 -8 32 272
use FILL  FILL_0__2827_
timestamp 1701859473
transform -1 0 9210 0 -1 1830
box -12 -8 32 272
use FILL  FILL_0__2828_
timestamp 1701859473
transform 1 0 6930 0 -1 1830
box -12 -8 32 272
use FILL  FILL_0__2829_
timestamp 1701859473
transform -1 0 9950 0 1 2870
box -12 -8 32 272
use FILL  FILL_0__2830_
timestamp 1701859473
transform 1 0 8250 0 -1 3390
box -12 -8 32 272
use FILL  FILL_0__2831_
timestamp 1701859473
transform 1 0 8290 0 1 3910
box -12 -8 32 272
use FILL  FILL_0__2832_
timestamp 1701859473
transform -1 0 9270 0 1 2350
box -12 -8 32 272
use FILL  FILL_0__2833_
timestamp 1701859473
transform -1 0 9210 0 -1 3390
box -12 -8 32 272
use FILL  FILL_0__2834_
timestamp 1701859473
transform -1 0 8970 0 -1 3390
box -12 -8 32 272
use FILL  FILL_0__2835_
timestamp 1701859473
transform -1 0 9270 0 1 790
box -12 -8 32 272
use FILL  FILL_0__2836_
timestamp 1701859473
transform 1 0 8850 0 1 1310
box -12 -8 32 272
use FILL  FILL_0__2837_
timestamp 1701859473
transform -1 0 9530 0 1 1310
box -12 -8 32 272
use FILL  FILL_0__2838_
timestamp 1701859473
transform -1 0 9650 0 1 3390
box -12 -8 32 272
use FILL  FILL_0__2839_
timestamp 1701859473
transform -1 0 9690 0 -1 3390
box -12 -8 32 272
use FILL  FILL_0__2840_
timestamp 1701859473
transform 1 0 9010 0 -1 270
box -12 -8 32 272
use FILL  FILL_0__2841_
timestamp 1701859473
transform -1 0 8810 0 -1 270
box -12 -8 32 272
use FILL  FILL_0__2842_
timestamp 1701859473
transform 1 0 9230 0 -1 270
box -12 -8 32 272
use FILL  FILL_0__2843_
timestamp 1701859473
transform 1 0 9470 0 -1 270
box -12 -8 32 272
use FILL  FILL_0__2844_
timestamp 1701859473
transform 1 0 9270 0 1 270
box -12 -8 32 272
use FILL  FILL_0__2845_
timestamp 1701859473
transform -1 0 9950 0 1 270
box -12 -8 32 272
use FILL  FILL_0__2846_
timestamp 1701859473
transform 1 0 9690 0 1 270
box -12 -8 32 272
use FILL  FILL_0__2847_
timestamp 1701859473
transform -1 0 11090 0 -1 10670
box -12 -8 32 272
use FILL  FILL_0__2848_
timestamp 1701859473
transform -1 0 10570 0 -1 1310
box -12 -8 32 272
use FILL  FILL_0__2849_
timestamp 1701859473
transform -1 0 10910 0 1 1310
box -12 -8 32 272
use FILL  FILL_0__2850_
timestamp 1701859473
transform -1 0 11050 0 -1 1830
box -12 -8 32 272
use FILL  FILL_0__2851_
timestamp 1701859473
transform 1 0 10650 0 -1 3910
box -12 -8 32 272
use FILL  FILL_0__2852_
timestamp 1701859473
transform -1 0 8850 0 1 270
box -12 -8 32 272
use FILL  FILL_0__2853_
timestamp 1701859473
transform -1 0 9070 0 1 270
box -12 -8 32 272
use FILL  FILL_0__2854_
timestamp 1701859473
transform 1 0 10570 0 1 790
box -12 -8 32 272
use FILL  FILL_0__2855_
timestamp 1701859473
transform -1 0 9770 0 1 1310
box -12 -8 32 272
use FILL  FILL_0__2856_
timestamp 1701859473
transform -1 0 10430 0 1 1310
box -12 -8 32 272
use FILL  FILL_0__2857_
timestamp 1701859473
transform -1 0 10670 0 1 1310
box -12 -8 32 272
use FILL  FILL_0__2858_
timestamp 1701859473
transform -1 0 11030 0 1 1830
box -12 -8 32 272
use FILL  FILL_0__2859_
timestamp 1701859473
transform 1 0 10890 0 -1 3910
box -12 -8 32 272
use FILL  FILL_0__2860_
timestamp 1701859473
transform 1 0 10810 0 -1 3390
box -12 -8 32 272
use FILL  FILL_0__2861_
timestamp 1701859473
transform 1 0 9690 0 -1 270
box -12 -8 32 272
use FILL  FILL_0__2862_
timestamp 1701859473
transform 1 0 8550 0 -1 270
box -12 -8 32 272
use FILL  FILL_0__2863_
timestamp 1701859473
transform -1 0 10190 0 1 270
box -12 -8 32 272
use FILL  FILL_0__2864_
timestamp 1701859473
transform 1 0 10430 0 1 270
box -12 -8 32 272
use FILL  FILL_0__2865_
timestamp 1701859473
transform -1 0 10670 0 1 270
box -12 -8 32 272
use FILL  FILL_0__2866_
timestamp 1701859473
transform -1 0 11050 0 -1 790
box -12 -8 32 272
use FILL  FILL_0__2867_
timestamp 1701859473
transform 1 0 11010 0 -1 3390
box -12 -8 32 272
use FILL  FILL_0__2868_
timestamp 1701859473
transform 1 0 10990 0 1 790
box -12 -8 32 272
use FILL  FILL_0__2869_
timestamp 1701859473
transform 1 0 10110 0 1 790
box -12 -8 32 272
use FILL  FILL_0__2870_
timestamp 1701859473
transform -1 0 10330 0 1 790
box -12 -8 32 272
use FILL  FILL_0__2871_
timestamp 1701859473
transform -1 0 10770 0 1 790
box -12 -8 32 272
use FILL  FILL_0__2872_
timestamp 1701859473
transform -1 0 11110 0 1 1310
box -12 -8 32 272
use FILL  FILL_0__2873_
timestamp 1701859473
transform -1 0 9890 0 1 3390
box -12 -8 32 272
use FILL  FILL_0__2874_
timestamp 1701859473
transform -1 0 10130 0 1 3390
box -12 -8 32 272
use FILL  FILL_0__2875_
timestamp 1701859473
transform -1 0 10710 0 -1 4950
box -12 -8 32 272
use FILL  FILL_0__2876_
timestamp 1701859473
transform -1 0 9670 0 1 1830
box -12 -8 32 272
use FILL  FILL_0__2877_
timestamp 1701859473
transform 1 0 9850 0 1 1830
box -12 -8 32 272
use FILL  FILL_0__2878_
timestamp 1701859473
transform 1 0 9670 0 -1 1310
box -12 -8 32 272
use FILL  FILL_0__2879_
timestamp 1701859473
transform -1 0 9910 0 -1 1310
box -12 -8 32 272
use FILL  FILL_0__2880_
timestamp 1701859473
transform 1 0 9410 0 1 1830
box -12 -8 32 272
use FILL  FILL_0__2881_
timestamp 1701859473
transform 1 0 10790 0 -1 790
box -12 -8 32 272
use FILL  FILL_0__2882_
timestamp 1701859473
transform -1 0 9470 0 -1 1310
box -12 -8 32 272
use FILL  FILL_0__2883_
timestamp 1701859473
transform -1 0 10370 0 -1 1310
box -12 -8 32 272
use FILL  FILL_0__2884_
timestamp 1701859473
transform 1 0 11010 0 -1 1310
box -12 -8 32 272
use FILL  FILL_0__2885_
timestamp 1701859473
transform -1 0 10790 0 -1 1310
box -12 -8 32 272
use FILL  FILL_0__2886_
timestamp 1701859473
transform 1 0 10550 0 1 1830
box -12 -8 32 272
use FILL  FILL_0__2887_
timestamp 1701859473
transform 1 0 10110 0 -1 4430
box -12 -8 32 272
use FILL  FILL_0__2888_
timestamp 1701859473
transform -1 0 3930 0 1 5470
box -12 -8 32 272
use FILL  FILL_0__2889_
timestamp 1701859473
transform 1 0 6050 0 1 2350
box -12 -8 32 272
use FILL  FILL_0__2890_
timestamp 1701859473
transform -1 0 8330 0 1 5990
box -12 -8 32 272
use FILL  FILL_0__2891_
timestamp 1701859473
transform -1 0 8130 0 1 5990
box -12 -8 32 272
use FILL  FILL_0__2892_
timestamp 1701859473
transform 1 0 7350 0 -1 5470
box -12 -8 32 272
use FILL  FILL_0__2893_
timestamp 1701859473
transform 1 0 7170 0 1 5470
box -12 -8 32 272
use FILL  FILL_0__2894_
timestamp 1701859473
transform 1 0 6450 0 -1 6510
box -12 -8 32 272
use FILL  FILL_0__2895_
timestamp 1701859473
transform 1 0 6590 0 1 6510
box -12 -8 32 272
use FILL  FILL_0__2896_
timestamp 1701859473
transform -1 0 7850 0 -1 5470
box -12 -8 32 272
use FILL  FILL_0__2897_
timestamp 1701859473
transform 1 0 7650 0 1 5470
box -12 -8 32 272
use FILL  FILL_0__2898_
timestamp 1701859473
transform 1 0 7170 0 -1 6510
box -12 -8 32 272
use FILL  FILL_0__2899_
timestamp 1701859473
transform 1 0 6690 0 -1 6510
box -12 -8 32 272
use FILL  FILL_0__2900_
timestamp 1701859473
transform -1 0 6230 0 -1 6510
box -12 -8 32 272
use FILL  FILL_0__2901_
timestamp 1701859473
transform 1 0 5970 0 -1 6510
box -12 -8 32 272
use FILL  FILL_0__2902_
timestamp 1701859473
transform -1 0 7890 0 1 5990
box -12 -8 32 272
use FILL  FILL_0__2903_
timestamp 1701859473
transform 1 0 7170 0 1 5990
box -12 -8 32 272
use FILL  FILL_0__2904_
timestamp 1701859473
transform 1 0 8290 0 -1 5470
box -12 -8 32 272
use FILL  FILL_0__2905_
timestamp 1701859473
transform 1 0 8310 0 1 5470
box -12 -8 32 272
use FILL  FILL_0__2906_
timestamp 1701859473
transform 1 0 8050 0 -1 5990
box -12 -8 32 272
use FILL  FILL_0__2907_
timestamp 1701859473
transform -1 0 7830 0 -1 5990
box -12 -8 32 272
use FILL  FILL_0__2908_
timestamp 1701859473
transform -1 0 8150 0 -1 4950
box -12 -8 32 272
use FILL  FILL_0__2909_
timestamp 1701859473
transform 1 0 3290 0 -1 4430
box -12 -8 32 272
use FILL  FILL_0__2910_
timestamp 1701859473
transform -1 0 6450 0 -1 4430
box -12 -8 32 272
use FILL  FILL_0__2911_
timestamp 1701859473
transform -1 0 6790 0 1 4430
box -12 -8 32 272
use FILL  FILL_0__2912_
timestamp 1701859473
transform 1 0 8570 0 -1 4950
box -12 -8 32 272
use FILL  FILL_0__2913_
timestamp 1701859473
transform -1 0 6750 0 -1 4950
box -12 -8 32 272
use FILL  FILL_0__2914_
timestamp 1701859473
transform 1 0 7010 0 -1 8070
box -12 -8 32 272
use FILL  FILL_0__2915_
timestamp 1701859473
transform 1 0 7130 0 -1 5990
box -12 -8 32 272
use FILL  FILL_0__2916_
timestamp 1701859473
transform 1 0 6890 0 -1 5990
box -12 -8 32 272
use FILL  FILL_0__2917_
timestamp 1701859473
transform -1 0 6270 0 -1 5990
box -12 -8 32 272
use FILL  FILL_0__2918_
timestamp 1701859473
transform 1 0 6190 0 1 5470
box -12 -8 32 272
use FILL  FILL_0__2919_
timestamp 1701859473
transform 1 0 6110 0 1 4950
box -12 -8 32 272
use FILL  FILL_0__2920_
timestamp 1701859473
transform 1 0 5870 0 1 4950
box -12 -8 32 272
use FILL  FILL_0__2921_
timestamp 1701859473
transform -1 0 7330 0 -1 3910
box -12 -8 32 272
use FILL  FILL_0__2922_
timestamp 1701859473
transform -1 0 7370 0 1 3910
box -12 -8 32 272
use FILL  FILL_0__2923_
timestamp 1701859473
transform -1 0 6690 0 -1 4430
box -12 -8 32 272
use FILL  FILL_0__2924_
timestamp 1701859473
transform 1 0 6310 0 1 4950
box -12 -8 32 272
use FILL  FILL_0__2925_
timestamp 1701859473
transform 1 0 7210 0 1 7550
box -12 -8 32 272
use FILL  FILL_0__2926_
timestamp 1701859473
transform -1 0 7450 0 1 4430
box -12 -8 32 272
use FILL  FILL_0__2927_
timestamp 1701859473
transform 1 0 7230 0 -1 4950
box -12 -8 32 272
use FILL  FILL_0__2928_
timestamp 1701859473
transform 1 0 6970 0 -1 4950
box -12 -8 32 272
use FILL  FILL_0__2929_
timestamp 1701859473
transform -1 0 6550 0 1 4950
box -12 -8 32 272
use FILL  FILL_0__2930_
timestamp 1701859473
transform 1 0 6090 0 1 1830
box -12 -8 32 272
use FILL  FILL_0__2931_
timestamp 1701859473
transform 1 0 6970 0 -1 2870
box -12 -8 32 272
use FILL  FILL_0__2932_
timestamp 1701859473
transform 1 0 5130 0 -1 4430
box -12 -8 32 272
use FILL  FILL_0__2933_
timestamp 1701859473
transform 1 0 5330 0 -1 4430
box -12 -8 32 272
use FILL  FILL_0__2934_
timestamp 1701859473
transform 1 0 5570 0 -1 4430
box -12 -8 32 272
use FILL  FILL_0__2935_
timestamp 1701859473
transform 1 0 6390 0 1 6510
box -12 -8 32 272
use FILL  FILL_0__2936_
timestamp 1701859473
transform 1 0 6270 0 -1 4950
box -12 -8 32 272
use FILL  FILL_0__2937_
timestamp 1701859473
transform 1 0 6490 0 -1 4950
box -12 -8 32 272
use FILL  FILL_0__2938_
timestamp 1701859473
transform 1 0 4970 0 1 4950
box -12 -8 32 272
use FILL  FILL_0__2939_
timestamp 1701859473
transform 1 0 4750 0 1 4950
box -12 -8 32 272
use FILL  FILL_0__2940_
timestamp 1701859473
transform -1 0 5810 0 -1 5470
box -12 -8 32 272
use FILL  FILL_0__2941_
timestamp 1701859473
transform 1 0 5570 0 -1 5470
box -12 -8 32 272
use FILL  FILL_0__2942_
timestamp 1701859473
transform -1 0 9270 0 1 4430
box -12 -8 32 272
use FILL  FILL_0__2943_
timestamp 1701859473
transform 1 0 6230 0 -1 4430
box -12 -8 32 272
use FILL  FILL_0__2944_
timestamp 1701859473
transform -1 0 6250 0 1 3910
box -12 -8 32 272
use FILL  FILL_0__2945_
timestamp 1701859473
transform -1 0 6330 0 1 4430
box -12 -8 32 272
use FILL  FILL_0__2946_
timestamp 1701859473
transform 1 0 6090 0 1 4430
box -12 -8 32 272
use FILL  FILL_0__2947_
timestamp 1701859473
transform -1 0 6490 0 -1 5990
box -12 -8 32 272
use FILL  FILL_0__2948_
timestamp 1701859473
transform 1 0 6030 0 -1 5990
box -12 -8 32 272
use FILL  FILL_0__2949_
timestamp 1701859473
transform -1 0 5850 0 -1 5990
box -12 -8 32 272
use FILL  FILL_0__2950_
timestamp 1701859473
transform 1 0 5710 0 1 5470
box -12 -8 32 272
use FILL  FILL_0__2951_
timestamp 1701859473
transform -1 0 5970 0 1 5470
box -12 -8 32 272
use FILL  FILL_0__2952_
timestamp 1701859473
transform -1 0 6050 0 -1 4950
box -12 -8 32 272
use FILL  FILL_0__2953_
timestamp 1701859473
transform -1 0 4330 0 1 4950
box -12 -8 32 272
use FILL  FILL_0__2954_
timestamp 1701859473
transform -1 0 6590 0 1 4430
box -12 -8 32 272
use FILL  FILL_0__2955_
timestamp 1701859473
transform -1 0 5870 0 1 4430
box -12 -8 32 272
use FILL  FILL_0__2956_
timestamp 1701859473
transform 1 0 5150 0 1 4430
box -12 -8 32 272
use FILL  FILL_0__2957_
timestamp 1701859473
transform 1 0 5090 0 -1 4950
box -12 -8 32 272
use FILL  FILL_0__2958_
timestamp 1701859473
transform -1 0 5410 0 1 4430
box -12 -8 32 272
use FILL  FILL_0__2959_
timestamp 1701859473
transform 1 0 6910 0 -1 5470
box -12 -8 32 272
use FILL  FILL_0__2960_
timestamp 1701859473
transform -1 0 6450 0 1 5470
box -12 -8 32 272
use FILL  FILL_0__2961_
timestamp 1701859473
transform 1 0 6210 0 -1 5470
box -12 -8 32 272
use FILL  FILL_0__2962_
timestamp 1701859473
transform -1 0 6470 0 -1 5470
box -12 -8 32 272
use FILL  FILL_0__2963_
timestamp 1701859473
transform -1 0 6710 0 -1 5470
box -12 -8 32 272
use FILL  FILL_0__2964_
timestamp 1701859473
transform -1 0 5350 0 -1 4950
box -12 -8 32 272
use FILL  FILL_0__2965_
timestamp 1701859473
transform 1 0 4850 0 -1 4950
box -12 -8 32 272
use FILL  FILL_0__2966_
timestamp 1701859473
transform -1 0 6310 0 1 2350
box -12 -8 32 272
use FILL  FILL_0__2967_
timestamp 1701859473
transform 1 0 7570 0 1 3910
box -12 -8 32 272
use FILL  FILL_0__2968_
timestamp 1701859473
transform -1 0 6890 0 -1 3910
box -12 -8 32 272
use FILL  FILL_0__2969_
timestamp 1701859473
transform -1 0 7110 0 -1 3910
box -12 -8 32 272
use FILL  FILL_0__2970_
timestamp 1701859473
transform -1 0 7150 0 1 3910
box -12 -8 32 272
use FILL  FILL_0__2971_
timestamp 1701859473
transform -1 0 6670 0 1 3910
box -12 -8 32 272
use FILL  FILL_0__2972_
timestamp 1701859473
transform 1 0 6890 0 1 3910
box -12 -8 32 272
use FILL  FILL_0__2973_
timestamp 1701859473
transform -1 0 7010 0 1 4430
box -12 -8 32 272
use FILL  FILL_0__2974_
timestamp 1701859473
transform 1 0 6910 0 -1 4430
box -12 -8 32 272
use FILL  FILL_0__2975_
timestamp 1701859473
transform -1 0 7670 0 -1 4430
box -12 -8 32 272
use FILL  FILL_0__2976_
timestamp 1701859473
transform -1 0 7430 0 -1 4430
box -12 -8 32 272
use FILL  FILL_0__2977_
timestamp 1701859473
transform 1 0 7150 0 -1 4430
box -12 -8 32 272
use FILL  FILL_0__2978_
timestamp 1701859473
transform 1 0 7210 0 1 4430
box -12 -8 32 272
use FILL  FILL_0__2979_
timestamp 1701859473
transform -1 0 3550 0 -1 4950
box -12 -8 32 272
use FILL  FILL_0__2980_
timestamp 1701859473
transform -1 0 2930 0 1 7550
box -12 -8 32 272
use FILL  FILL_0__2981_
timestamp 1701859473
transform 1 0 3450 0 1 4950
box -12 -8 32 272
use FILL  FILL_0__2982_
timestamp 1701859473
transform 1 0 9510 0 1 6510
box -12 -8 32 272
use FILL  FILL_0__2983_
timestamp 1701859473
transform 1 0 1830 0 1 4430
box -12 -8 32 272
use FILL  FILL_0__2984_
timestamp 1701859473
transform -1 0 3450 0 -1 3910
box -12 -8 32 272
use FILL  FILL_0__2985_
timestamp 1701859473
transform 1 0 3610 0 1 4430
box -12 -8 32 272
use FILL  FILL_0__2986_
timestamp 1701859473
transform -1 0 5810 0 -1 4430
box -12 -8 32 272
use FILL  FILL_0__2987_
timestamp 1701859473
transform -1 0 5630 0 1 4430
box -12 -8 32 272
use FILL  FILL_0__2988_
timestamp 1701859473
transform 1 0 9290 0 1 6510
box -12 -8 32 272
use FILL  FILL_0__2989_
timestamp 1701859473
transform 1 0 5910 0 1 6510
box -12 -8 32 272
use FILL  FILL_0__2990_
timestamp 1701859473
transform -1 0 6170 0 1 6510
box -12 -8 32 272
use FILL  FILL_0__2991_
timestamp 1701859473
transform 1 0 7070 0 1 6510
box -12 -8 32 272
use FILL  FILL_0__2992_
timestamp 1701859473
transform 1 0 9590 0 1 7030
box -12 -8 32 272
use FILL  FILL_0__2993_
timestamp 1701859473
transform 1 0 9790 0 1 7030
box -12 -8 32 272
use FILL  FILL_0__2994_
timestamp 1701859473
transform -1 0 10710 0 -1 7550
box -12 -8 32 272
use FILL  FILL_0__2995_
timestamp 1701859473
transform -1 0 7510 0 -1 7550
box -12 -8 32 272
use FILL  FILL_0__2996_
timestamp 1701859473
transform 1 0 7410 0 1 7550
box -12 -8 32 272
use FILL  FILL_0__2997_
timestamp 1701859473
transform -1 0 7290 0 -1 7550
box -12 -8 32 272
use FILL  FILL_0__2998_
timestamp 1701859473
transform -1 0 6350 0 -1 7550
box -12 -8 32 272
use FILL  FILL_0__2999_
timestamp 1701859473
transform 1 0 6070 0 1 7550
box -12 -8 32 272
use FILL  FILL_0__3000_
timestamp 1701859473
transform -1 0 5910 0 -1 7550
box -12 -8 32 272
use FILL  FILL_0__3001_
timestamp 1701859473
transform -1 0 5690 0 -1 7550
box -12 -8 32 272
use FILL  FILL_0__3002_
timestamp 1701859473
transform -1 0 6110 0 -1 7550
box -12 -8 32 272
use FILL  FILL_0__3003_
timestamp 1701859473
transform -1 0 6290 0 1 7550
box -12 -8 32 272
use FILL  FILL_0__3004_
timestamp 1701859473
transform 1 0 8090 0 1 7550
box -12 -8 32 272
use FILL  FILL_0__3005_
timestamp 1701859473
transform 1 0 10910 0 -1 7550
box -12 -8 32 272
use FILL  FILL_0__3006_
timestamp 1701859473
transform -1 0 10390 0 1 7550
box -12 -8 32 272
use FILL  FILL_0__3007_
timestamp 1701859473
transform 1 0 6910 0 1 7030
box -12 -8 32 272
use FILL  FILL_0__3008_
timestamp 1701859473
transform -1 0 6470 0 1 7030
box -12 -8 32 272
use FILL  FILL_0__3009_
timestamp 1701859473
transform -1 0 5870 0 -1 7030
box -12 -8 32 272
use FILL  FILL_0__3010_
timestamp 1701859473
transform 1 0 6090 0 -1 7030
box -12 -8 32 272
use FILL  FILL_0__3011_
timestamp 1701859473
transform 1 0 6670 0 1 7030
box -12 -8 32 272
use FILL  FILL_0__3012_
timestamp 1701859473
transform -1 0 7790 0 -1 7030
box -12 -8 32 272
use FILL  FILL_0__3013_
timestamp 1701859473
transform 1 0 8230 0 -1 7030
box -12 -8 32 272
use FILL  FILL_0__3014_
timestamp 1701859473
transform 1 0 10590 0 1 7550
box -12 -8 32 272
use FILL  FILL_0__3015_
timestamp 1701859473
transform -1 0 6310 0 -1 7030
box -12 -8 32 272
use FILL  FILL_0__3016_
timestamp 1701859473
transform -1 0 7190 0 1 7030
box -12 -8 32 272
use FILL  FILL_0__3017_
timestamp 1701859473
transform 1 0 6530 0 -1 7030
box -12 -8 32 272
use FILL  FILL_0__3018_
timestamp 1701859473
transform -1 0 6830 0 -1 7030
box -12 -8 32 272
use FILL  FILL_0__3019_
timestamp 1701859473
transform -1 0 7070 0 -1 7030
box -12 -8 32 272
use FILL  FILL_0__3020_
timestamp 1701859473
transform 1 0 8230 0 1 7030
box -12 -8 32 272
use FILL  FILL_0__3021_
timestamp 1701859473
transform -1 0 9290 0 -1 8070
box -12 -8 32 272
use FILL  FILL_0__3022_
timestamp 1701859473
transform 1 0 9470 0 -1 8070
box -12 -8 32 272
use FILL  FILL_0__3023_
timestamp 1701859473
transform -1 0 5690 0 1 6510
box -12 -8 32 272
use FILL  FILL_0__3024_
timestamp 1701859473
transform 1 0 5430 0 1 6510
box -12 -8 32 272
use FILL  FILL_0__3025_
timestamp 1701859473
transform -1 0 5450 0 -1 6510
box -12 -8 32 272
use FILL  FILL_0__3026_
timestamp 1701859473
transform 1 0 10870 0 -1 5990
box -12 -8 32 272
use FILL  FILL_0__3027_
timestamp 1701859473
transform -1 0 11110 0 -1 5990
box -12 -8 32 272
use FILL  FILL_0__3028_
timestamp 1701859473
transform -1 0 9730 0 -1 8070
box -12 -8 32 272
use FILL  FILL_0__3029_
timestamp 1701859473
transform -1 0 7050 0 -1 7550
box -12 -8 32 272
use FILL  FILL_0__3030_
timestamp 1701859473
transform -1 0 8030 0 -1 7030
box -12 -8 32 272
use FILL  FILL_0__3031_
timestamp 1701859473
transform 1 0 8010 0 1 7030
box -12 -8 32 272
use FILL  FILL_0__3032_
timestamp 1701859473
transform 1 0 7630 0 1 7550
box -12 -8 32 272
use FILL  FILL_0__3033_
timestamp 1701859473
transform -1 0 6710 0 1 8070
box -12 -8 32 272
use FILL  FILL_0__3034_
timestamp 1701859473
transform -1 0 7690 0 -1 8070
box -12 -8 32 272
use FILL  FILL_0__3035_
timestamp 1701859473
transform 1 0 7430 0 -1 8070
box -12 -8 32 272
use FILL  FILL_0__3036_
timestamp 1701859473
transform -1 0 6910 0 1 8070
box -12 -8 32 272
use FILL  FILL_0__3037_
timestamp 1701859473
transform -1 0 6470 0 1 8070
box -12 -8 32 272
use FILL  FILL_0__3038_
timestamp 1701859473
transform -1 0 7090 0 1 8070
box -12 -8 32 272
use FILL  FILL_0__3039_
timestamp 1701859473
transform 1 0 7310 0 1 8070
box -12 -8 32 272
use FILL  FILL_0__3040_
timestamp 1701859473
transform 1 0 9650 0 1 7550
box -12 -8 32 272
use FILL  FILL_0__3041_
timestamp 1701859473
transform -1 0 9510 0 -1 6510
box -12 -8 32 272
use FILL  FILL_0__3042_
timestamp 1701859473
transform 1 0 7210 0 -1 8070
box -12 -8 32 272
use FILL  FILL_0__3043_
timestamp 1701859473
transform -1 0 6530 0 1 7550
box -12 -8 32 272
use FILL  FILL_0__3044_
timestamp 1701859473
transform -1 0 6570 0 -1 7550
box -12 -8 32 272
use FILL  FILL_0__3045_
timestamp 1701859473
transform 1 0 6790 0 -1 7550
box -12 -8 32 272
use FILL  FILL_0__3046_
timestamp 1701859473
transform -1 0 7750 0 1 6510
box -12 -8 32 272
use FILL  FILL_0__3047_
timestamp 1701859473
transform 1 0 9090 0 1 6510
box -12 -8 32 272
use FILL  FILL_0__3048_
timestamp 1701859473
transform 1 0 9710 0 -1 6510
box -12 -8 32 272
use FILL  FILL_0__3049_
timestamp 1701859473
transform -1 0 6790 0 1 7550
box -12 -8 32 272
use FILL  FILL_0__3050_
timestamp 1701859473
transform -1 0 7010 0 1 7550
box -12 -8 32 272
use FILL  FILL_0__3051_
timestamp 1701859473
transform -1 0 7750 0 1 7030
box -12 -8 32 272
use FILL  FILL_0__3052_
timestamp 1701859473
transform 1 0 7450 0 1 7030
box -12 -8 32 272
use FILL  FILL_0__3053_
timestamp 1701859473
transform 1 0 7290 0 -1 7030
box -12 -8 32 272
use FILL  FILL_0__3054_
timestamp 1701859473
transform -1 0 7550 0 -1 7030
box -12 -8 32 272
use FILL  FILL_0__3055_
timestamp 1701859473
transform 1 0 7970 0 1 6510
box -12 -8 32 272
use FILL  FILL_0__3056_
timestamp 1701859473
transform -1 0 9490 0 1 5470
box -12 -8 32 272
use FILL  FILL_0__3057_
timestamp 1701859473
transform -1 0 9250 0 1 5470
box -12 -8 32 272
use FILL  FILL_0__3058_
timestamp 1701859473
transform 1 0 8670 0 -1 7550
box -12 -8 32 272
use FILL  FILL_0__3059_
timestamp 1701859473
transform -1 0 8550 0 -1 5990
box -12 -8 32 272
use FILL  FILL_0__3060_
timestamp 1701859473
transform 1 0 9730 0 1 6510
box -12 -8 32 272
use FILL  FILL_0__3061_
timestamp 1701859473
transform 1 0 9970 0 1 6510
box -12 -8 32 272
use FILL  FILL_0__3062_
timestamp 1701859473
transform -1 0 9590 0 -1 7550
box -12 -8 32 272
use FILL  FILL_0__3063_
timestamp 1701859473
transform 1 0 9330 0 -1 7550
box -12 -8 32 272
use FILL  FILL_0__3064_
timestamp 1701859473
transform -1 0 10290 0 -1 7030
box -12 -8 32 272
use FILL  FILL_0__3065_
timestamp 1701859473
transform -1 0 10530 0 -1 7030
box -12 -8 32 272
use FILL  FILL_0__3066_
timestamp 1701859473
transform -1 0 8450 0 -1 7550
box -12 -8 32 272
use FILL  FILL_0__3067_
timestamp 1701859473
transform 1 0 8190 0 -1 7550
box -12 -8 32 272
use FILL  FILL_0__3068_
timestamp 1701859473
transform 1 0 10150 0 -1 5990
box -12 -8 32 272
use FILL  FILL_0__3069_
timestamp 1701859473
transform 1 0 10390 0 -1 5990
box -12 -8 32 272
use FILL  FILL_0__3070_
timestamp 1701859473
transform 1 0 8850 0 -1 7550
box -12 -8 32 272
use FILL  FILL_0__3071_
timestamp 1701859473
transform -1 0 9110 0 -1 7550
box -12 -8 32 272
use FILL  FILL_0__3072_
timestamp 1701859473
transform -1 0 9730 0 1 5990
box -12 -8 32 272
use FILL  FILL_0__3073_
timestamp 1701859473
transform -1 0 9950 0 1 5990
box -12 -8 32 272
use FILL  FILL_0__3074_
timestamp 1701859473
transform 1 0 8770 0 1 5990
box -12 -8 32 272
use FILL  FILL_0__3075_
timestamp 1701859473
transform 1 0 8770 0 -1 5990
box -12 -8 32 272
use FILL  FILL_0__3076_
timestamp 1701859473
transform 1 0 10670 0 1 6510
box -12 -8 32 272
use FILL  FILL_0__3077_
timestamp 1701859473
transform 1 0 10870 0 1 6510
box -12 -8 32 272
use FILL  FILL_0__3078_
timestamp 1701859473
transform -1 0 8670 0 -1 7030
box -12 -8 32 272
use FILL  FILL_0__3079_
timestamp 1701859473
transform -1 0 8450 0 -1 7030
box -12 -8 32 272
use FILL  FILL_0__3080_
timestamp 1701859473
transform 1 0 10930 0 -1 8590
box -12 -8 32 272
use FILL  FILL_0__3081_
timestamp 1701859473
transform -1 0 10930 0 -1 270
box -12 -8 32 272
use FILL  FILL_0__3082_
timestamp 1701859473
transform 1 0 10030 0 -1 8590
box -12 -8 32 272
use FILL  FILL_0__3083_
timestamp 1701859473
transform -1 0 9810 0 -1 8590
box -12 -8 32 272
use FILL  FILL_0__3084_
timestamp 1701859473
transform -1 0 8990 0 1 7550
box -12 -8 32 272
use FILL  FILL_0__3085_
timestamp 1701859473
transform 1 0 8890 0 1 7030
box -12 -8 32 272
use FILL  FILL_0__3086_
timestamp 1701859473
transform -1 0 10650 0 1 5990
box -12 -8 32 272
use FILL  FILL_0__3087_
timestamp 1701859473
transform 1 0 10850 0 1 5990
box -12 -8 32 272
use FILL  FILL_0__3088_
timestamp 1701859473
transform 1 0 8210 0 1 8070
box -12 -8 32 272
use FILL  FILL_0__3089_
timestamp 1701859473
transform -1 0 7990 0 1 8070
box -12 -8 32 272
use FILL  FILL_0__3090_
timestamp 1701859473
transform -1 0 11090 0 1 4950
box -12 -8 32 272
use FILL  FILL_0__3091_
timestamp 1701859473
transform 1 0 10830 0 1 4950
box -12 -8 32 272
use FILL  FILL_0__3092_
timestamp 1701859473
transform 1 0 8750 0 -1 5470
box -12 -8 32 272
use FILL  FILL_0__3093_
timestamp 1701859473
transform -1 0 8990 0 -1 5470
box -12 -8 32 272
use FILL  FILL_0__3094_
timestamp 1701859473
transform -1 0 10190 0 -1 5470
box -12 -8 32 272
use FILL  FILL_0__3095_
timestamp 1701859473
transform 1 0 10130 0 1 5470
box -12 -8 32 272
use FILL  FILL_0__3096_
timestamp 1701859473
transform 1 0 8870 0 1 6510
box -12 -8 32 272
use FILL  FILL_0__3097_
timestamp 1701859473
transform -1 0 8650 0 1 6510
box -12 -8 32 272
use FILL  FILL_0__3098_
timestamp 1701859473
transform -1 0 10350 0 1 8070
box -12 -8 32 272
use FILL  FILL_0__3099_
timestamp 1701859473
transform -1 0 11110 0 -1 8070
box -12 -8 32 272
use FILL  FILL_0__3100_
timestamp 1701859473
transform 1 0 10110 0 1 8070
box -12 -8 32 272
use FILL  FILL_0__3101_
timestamp 1701859473
transform 1 0 10250 0 -1 8590
box -12 -8 32 272
use FILL  FILL_0__3102_
timestamp 1701859473
transform 1 0 8330 0 -1 8070
box -12 -8 32 272
use FILL  FILL_0__3103_
timestamp 1701859473
transform -1 0 8310 0 1 7550
box -12 -8 32 272
use FILL  FILL_0__3104_
timestamp 1701859473
transform -1 0 11110 0 1 6510
box -12 -8 32 272
use FILL  FILL_0__3105_
timestamp 1701859473
transform -1 0 10910 0 -1 4950
box -12 -8 32 272
use FILL  FILL_0__3106_
timestamp 1701859473
transform 1 0 9330 0 -1 8590
box -12 -8 32 272
use FILL  FILL_0__3107_
timestamp 1701859473
transform -1 0 9570 0 -1 8590
box -12 -8 32 272
use FILL  FILL_0__3108_
timestamp 1701859473
transform 1 0 9930 0 1 5470
box -12 -8 32 272
use FILL  FILL_0__3109_
timestamp 1701859473
transform -1 0 9710 0 1 5470
box -12 -8 32 272
use FILL  FILL_0__3110_
timestamp 1701859473
transform 1 0 8350 0 -1 6510
box -12 -8 32 272
use FILL  FILL_0__3111_
timestamp 1701859473
transform -1 0 8130 0 -1 6510
box -12 -8 32 272
use FILL  FILL_0__3112_
timestamp 1701859473
transform 1 0 470 0 -1 2870
box -12 -8 32 272
use FILL  FILL_0__3113_
timestamp 1701859473
transform 1 0 10 0 -1 2870
box -12 -8 32 272
use FILL  FILL_0__3114_
timestamp 1701859473
transform -1 0 270 0 -1 2870
box -12 -8 32 272
use FILL  FILL_0__3115_
timestamp 1701859473
transform -1 0 1150 0 1 2350
box -12 -8 32 272
use FILL  FILL_0__3116_
timestamp 1701859473
transform 1 0 910 0 -1 2350
box -12 -8 32 272
use FILL  FILL_0__3117_
timestamp 1701859473
transform 1 0 1990 0 -1 1310
box -12 -8 32 272
use FILL  FILL_0__3118_
timestamp 1701859473
transform -1 0 1370 0 -1 2350
box -12 -8 32 272
use FILL  FILL_0__3119_
timestamp 1701859473
transform -1 0 1130 0 -1 2350
box -12 -8 32 272
use FILL  FILL_0__3120_
timestamp 1701859473
transform -1 0 430 0 1 2350
box -12 -8 32 272
use FILL  FILL_0__3121_
timestamp 1701859473
transform 1 0 210 0 1 2870
box -12 -8 32 272
use FILL  FILL_0__3122_
timestamp 1701859473
transform 1 0 2470 0 -1 3390
box -12 -8 32 272
use FILL  FILL_0__3123_
timestamp 1701859473
transform 1 0 490 0 1 3390
box -12 -8 32 272
use FILL  FILL_0__3124_
timestamp 1701859473
transform -1 0 270 0 1 3390
box -12 -8 32 272
use FILL  FILL_0__3125_
timestamp 1701859473
transform -1 0 690 0 -1 2350
box -12 -8 32 272
use FILL  FILL_0__3126_
timestamp 1701859473
transform -1 0 1390 0 1 2350
box -12 -8 32 272
use FILL  FILL_0__3127_
timestamp 1701859473
transform -1 0 910 0 1 2350
box -12 -8 32 272
use FILL  FILL_0__3128_
timestamp 1701859473
transform -1 0 1850 0 1 2350
box -12 -8 32 272
use FILL  FILL_0__3129_
timestamp 1701859473
transform -1 0 1610 0 -1 2350
box -12 -8 32 272
use FILL  FILL_0__3130_
timestamp 1701859473
transform -1 0 1630 0 1 2350
box -12 -8 32 272
use FILL  FILL_0__3131_
timestamp 1701859473
transform -1 0 670 0 1 2350
box -12 -8 32 272
use FILL  FILL_0__3132_
timestamp 1701859473
transform 1 0 430 0 1 2870
box -12 -8 32 272
use FILL  FILL_0__3133_
timestamp 1701859473
transform 1 0 490 0 -1 3910
box -12 -8 32 272
use FILL  FILL_0__3134_
timestamp 1701859473
transform -1 0 1170 0 1 3390
box -12 -8 32 272
use FILL  FILL_0__3135_
timestamp 1701859473
transform 1 0 930 0 1 3390
box -12 -8 32 272
use FILL  FILL_0__3136_
timestamp 1701859473
transform -1 0 510 0 -1 3390
box -12 -8 32 272
use FILL  FILL_0__3137_
timestamp 1701859473
transform 1 0 230 0 -1 3390
box -12 -8 32 272
use FILL  FILL_0__3138_
timestamp 1701859473
transform -1 0 1630 0 1 4430
box -12 -8 32 272
use FILL  FILL_0__3139_
timestamp 1701859473
transform -1 0 1830 0 -1 3390
box -12 -8 32 272
use FILL  FILL_0__3140_
timestamp 1701859473
transform -1 0 250 0 1 3910
box -12 -8 32 272
use FILL  FILL_0__3141_
timestamp 1701859473
transform 1 0 690 0 1 4430
box -12 -8 32 272
use FILL  FILL_0__3142_
timestamp 1701859473
transform 1 0 930 0 1 4430
box -12 -8 32 272
use FILL  FILL_0__3143_
timestamp 1701859473
transform 1 0 950 0 -1 4430
box -12 -8 32 272
use FILL  FILL_0__3144_
timestamp 1701859473
transform -1 0 1190 0 -1 4430
box -12 -8 32 272
use FILL  FILL_0__3145_
timestamp 1701859473
transform -1 0 470 0 1 3910
box -12 -8 32 272
use FILL  FILL_0__3146_
timestamp 1701859473
transform -1 0 690 0 1 3910
box -12 -8 32 272
use FILL  FILL_0__3147_
timestamp 1701859473
transform 1 0 470 0 -1 4430
box -12 -8 32 272
use FILL  FILL_0__3148_
timestamp 1701859473
transform -1 0 730 0 -1 4430
box -12 -8 32 272
use FILL  FILL_0__3149_
timestamp 1701859473
transform -1 0 30 0 -1 3910
box -12 -8 32 272
use FILL  FILL_0__3150_
timestamp 1701859473
transform -1 0 890 0 1 3910
box -12 -8 32 272
use FILL  FILL_0__3151_
timestamp 1701859473
transform 1 0 10 0 1 3910
box -12 -8 32 272
use FILL  FILL_0__3152_
timestamp 1701859473
transform 1 0 10 0 -1 4430
box -12 -8 32 272
use FILL  FILL_0__3153_
timestamp 1701859473
transform -1 0 250 0 -1 4430
box -12 -8 32 272
use FILL  FILL_0__3154_
timestamp 1701859473
transform -1 0 750 0 -1 3390
box -12 -8 32 272
use FILL  FILL_0__3155_
timestamp 1701859473
transform -1 0 30 0 1 2870
box -12 -8 32 272
use FILL  FILL_0__3156_
timestamp 1701859473
transform 1 0 10 0 -1 3390
box -12 -8 32 272
use FILL  FILL_0__3157_
timestamp 1701859473
transform -1 0 30 0 1 3390
box -12 -8 32 272
use FILL  FILL_0__3158_
timestamp 1701859473
transform 1 0 10 0 1 4430
box -12 -8 32 272
use FILL  FILL_0__3159_
timestamp 1701859473
transform 1 0 230 0 1 4430
box -12 -8 32 272
use FILL  FILL_0__3160_
timestamp 1701859473
transform -1 0 470 0 1 4430
box -12 -8 32 272
use FILL  FILL_0__3161_
timestamp 1701859473
transform 1 0 4110 0 -1 7030
box -12 -8 32 272
use FILL  FILL_0__3162_
timestamp 1701859473
transform -1 0 4350 0 -1 7030
box -12 -8 32 272
use FILL  FILL_0__3163_
timestamp 1701859473
transform 1 0 4570 0 -1 7030
box -12 -8 32 272
use FILL  FILL_0__3164_
timestamp 1701859473
transform 1 0 4810 0 1 7030
box -12 -8 32 272
use FILL  FILL_0__3165_
timestamp 1701859473
transform 1 0 4070 0 1 7550
box -12 -8 32 272
use FILL  FILL_0__3166_
timestamp 1701859473
transform -1 0 4310 0 1 7550
box -12 -8 32 272
use FILL  FILL_0__3167_
timestamp 1701859473
transform 1 0 4790 0 -1 10150
box -12 -8 32 272
use FILL  FILL_0__3168_
timestamp 1701859473
transform 1 0 4990 0 -1 10150
box -12 -8 32 272
use FILL  FILL_0__3169_
timestamp 1701859473
transform -1 0 3630 0 -1 10670
box -12 -8 32 272
use FILL  FILL_0__3170_
timestamp 1701859473
transform -1 0 3850 0 -1 10670
box -12 -8 32 272
use FILL  FILL_0__3171_
timestamp 1701859473
transform 1 0 4270 0 -1 10670
box -12 -8 32 272
use FILL  FILL_0__3172_
timestamp 1701859473
transform -1 0 4510 0 -1 10670
box -12 -8 32 272
use FILL  FILL_0__3173_
timestamp 1701859473
transform 1 0 4110 0 1 10150
box -12 -8 32 272
use FILL  FILL_0__3174_
timestamp 1701859473
transform -1 0 4350 0 1 10150
box -12 -8 32 272
use FILL  FILL_0__3175_
timestamp 1701859473
transform 1 0 5450 0 1 10150
box -12 -8 32 272
use FILL  FILL_0__3176_
timestamp 1701859473
transform 1 0 5210 0 1 10150
box -12 -8 32 272
use FILL  FILL_0__3177_
timestamp 1701859473
transform -1 0 1690 0 -1 5990
box -12 -8 32 272
use FILL  FILL_0__3178_
timestamp 1701859473
transform 1 0 2130 0 -1 5990
box -12 -8 32 272
use FILL  FILL_0__3179_
timestamp 1701859473
transform -1 0 1410 0 1 6510
box -12 -8 32 272
use FILL  FILL_0__3180_
timestamp 1701859473
transform -1 0 1630 0 1 6510
box -12 -8 32 272
use FILL  FILL_0__3181_
timestamp 1701859473
transform -1 0 490 0 -1 6510
box -12 -8 32 272
use FILL  FILL_0__3182_
timestamp 1701859473
transform -1 0 890 0 -1 6510
box -12 -8 32 272
use FILL  FILL_0__3183_
timestamp 1701859473
transform 1 0 250 0 1 8070
box -12 -8 32 272
use FILL  FILL_0__3184_
timestamp 1701859473
transform -1 0 490 0 1 8070
box -12 -8 32 272
use FILL  FILL_0__3185_
timestamp 1701859473
transform -1 0 30 0 -1 8590
box -12 -8 32 272
use FILL  FILL_0__3186_
timestamp 1701859473
transform -1 0 30 0 1 8070
box -12 -8 32 272
use FILL  FILL_0__3187_
timestamp 1701859473
transform 1 0 650 0 -1 9110
box -12 -8 32 272
use FILL  FILL_0__3188_
timestamp 1701859473
transform 1 0 870 0 -1 9110
box -12 -8 32 272
use FILL  FILL_0__3189_
timestamp 1701859473
transform 1 0 2050 0 -1 9630
box -12 -8 32 272
use FILL  FILL_0__3190_
timestamp 1701859473
transform 1 0 2290 0 1 9110
box -12 -8 32 272
use FILL  FILL_0__3191_
timestamp 1701859473
transform 1 0 1350 0 -1 9110
box -12 -8 32 272
use FILL  FILL_0__3192_
timestamp 1701859473
transform -1 0 1590 0 -1 9110
box -12 -8 32 272
use FILL  FILL_0__3324_
timestamp 1701859473
transform 1 0 5530 0 1 8070
box -12 -8 32 272
use FILL  FILL_0__3325_
timestamp 1701859473
transform -1 0 6250 0 1 8070
box -12 -8 32 272
use FILL  FILL_0__3326_
timestamp 1701859473
transform -1 0 6150 0 -1 8070
box -12 -8 32 272
use FILL  FILL_0__3327_
timestamp 1701859473
transform -1 0 6110 0 -1 8590
box -12 -8 32 272
use FILL  FILL_0__3328_
timestamp 1701859473
transform -1 0 6010 0 1 8070
box -12 -8 32 272
use FILL  FILL_0__3329_
timestamp 1701859473
transform 1 0 5770 0 1 8070
box -12 -8 32 272
use FILL  FILL_0__3330_
timestamp 1701859473
transform -1 0 6950 0 1 8590
box -12 -8 32 272
use FILL  FILL_0__3331_
timestamp 1701859473
transform 1 0 7230 0 -1 8590
box -12 -8 32 272
use FILL  FILL_0__3332_
timestamp 1701859473
transform 1 0 6950 0 -1 8590
box -12 -8 32 272
use FILL  FILL_0__3333_
timestamp 1701859473
transform 1 0 10150 0 1 8590
box -12 -8 32 272
use FILL  FILL_0__3334_
timestamp 1701859473
transform 1 0 9270 0 1 8590
box -12 -8 32 272
use FILL  FILL_0__3335_
timestamp 1701859473
transform 1 0 7810 0 -1 10150
box -12 -8 32 272
use FILL  FILL_0__3336_
timestamp 1701859473
transform -1 0 6650 0 1 9630
box -12 -8 32 272
use FILL  FILL_0__3337_
timestamp 1701859473
transform -1 0 6170 0 1 9630
box -12 -8 32 272
use FILL  FILL_0__3338_
timestamp 1701859473
transform 1 0 7130 0 -1 10150
box -12 -8 32 272
use FILL  FILL_0__3339_
timestamp 1701859473
transform -1 0 8010 0 1 10150
box -12 -8 32 272
use FILL  FILL_0__3340_
timestamp 1701859473
transform 1 0 7770 0 1 10150
box -12 -8 32 272
use FILL  FILL_0__3341_
timestamp 1701859473
transform 1 0 7530 0 1 10150
box -12 -8 32 272
use FILL  FILL_0__3342_
timestamp 1701859473
transform 1 0 6750 0 -1 11190
box -12 -8 32 272
use FILL  FILL_0__3343_
timestamp 1701859473
transform -1 0 7350 0 -1 10150
box -12 -8 32 272
use FILL  FILL_0__3344_
timestamp 1701859473
transform 1 0 7570 0 -1 10150
box -12 -8 32 272
use FILL  FILL_0__3345_
timestamp 1701859473
transform -1 0 8950 0 1 9630
box -12 -8 32 272
use FILL  FILL_0__3346_
timestamp 1701859473
transform 1 0 8470 0 1 10150
box -12 -8 32 272
use FILL  FILL_0__3347_
timestamp 1701859473
transform -1 0 8250 0 1 10150
box -12 -8 32 272
use FILL  FILL_0__3348_
timestamp 1701859473
transform 1 0 9070 0 -1 10670
box -12 -8 32 272
use FILL  FILL_0__3349_
timestamp 1701859473
transform 1 0 7810 0 1 9630
box -12 -8 32 272
use FILL  FILL_0__3350_
timestamp 1701859473
transform 1 0 7510 0 -1 8590
box -12 -8 32 272
use FILL  FILL_0__3351_
timestamp 1701859473
transform -1 0 7690 0 1 8590
box -12 -8 32 272
use FILL  FILL_0__3352_
timestamp 1701859473
transform -1 0 8150 0 -1 9110
box -12 -8 32 272
use FILL  FILL_0__3353_
timestamp 1701859473
transform 1 0 8030 0 -1 10150
box -12 -8 32 272
use FILL  FILL_0__3354_
timestamp 1701859473
transform 1 0 7710 0 -1 10670
box -12 -8 32 272
use FILL  FILL_0__3355_
timestamp 1701859473
transform -1 0 7490 0 -1 10670
box -12 -8 32 272
use FILL  FILL_0__3356_
timestamp 1701859473
transform 1 0 7270 0 -1 10670
box -12 -8 32 272
use FILL  FILL_0__3357_
timestamp 1701859473
transform 1 0 7090 0 1 10670
box -12 -8 32 272
use FILL  FILL_0__3358_
timestamp 1701859473
transform 1 0 7350 0 1 10670
box -12 -8 32 272
use FILL  FILL_0__3359_
timestamp 1701859473
transform 1 0 7590 0 1 10670
box -12 -8 32 272
use FILL  FILL_0__3360_
timestamp 1701859473
transform -1 0 7850 0 1 10670
box -12 -8 32 272
use FILL  FILL_0__3361_
timestamp 1701859473
transform 1 0 8870 0 -1 10670
box -12 -8 32 272
use FILL  FILL_0__3362_
timestamp 1701859473
transform 1 0 7930 0 -1 10670
box -12 -8 32 272
use FILL  FILL_0__3363_
timestamp 1701859473
transform 1 0 8050 0 1 10670
box -12 -8 32 272
use FILL  FILL_0__3364_
timestamp 1701859473
transform 1 0 7890 0 -1 11190
box -12 -8 32 272
use FILL  FILL_0__3365_
timestamp 1701859473
transform -1 0 7430 0 -1 11190
box -12 -8 32 272
use FILL  FILL_0__3366_
timestamp 1701859473
transform 1 0 6950 0 -1 11190
box -12 -8 32 272
use FILL  FILL_0__3367_
timestamp 1701859473
transform 1 0 6830 0 1 10670
box -12 -8 32 272
use FILL  FILL_0__3368_
timestamp 1701859473
transform 1 0 7170 0 -1 11190
box -12 -8 32 272
use FILL  FILL_0__3369_
timestamp 1701859473
transform 1 0 7650 0 -1 11190
box -12 -8 32 272
use FILL  FILL_0__3370_
timestamp 1701859473
transform 1 0 8170 0 -1 10670
box -12 -8 32 272
use FILL  FILL_0__3371_
timestamp 1701859473
transform 1 0 8270 0 1 10670
box -12 -8 32 272
use FILL  FILL_0__3372_
timestamp 1701859473
transform 1 0 9450 0 1 10670
box -12 -8 32 272
use FILL  FILL_0__3373_
timestamp 1701859473
transform -1 0 6550 0 -1 11190
box -12 -8 32 272
use FILL  FILL_0__3374_
timestamp 1701859473
transform 1 0 5650 0 1 10670
box -12 -8 32 272
use FILL  FILL_0__3375_
timestamp 1701859473
transform -1 0 5910 0 1 10670
box -12 -8 32 272
use FILL  FILL_0__3376_
timestamp 1701859473
transform -1 0 6130 0 1 10670
box -12 -8 32 272
use FILL  FILL_0__3377_
timestamp 1701859473
transform 1 0 6370 0 1 10670
box -12 -8 32 272
use FILL  FILL_0__3378_
timestamp 1701859473
transform 1 0 6310 0 -1 11190
box -12 -8 32 272
use FILL  FILL_0__3379_
timestamp 1701859473
transform 1 0 8630 0 -1 10670
box -12 -8 32 272
use FILL  FILL_0__3380_
timestamp 1701859473
transform 1 0 8750 0 1 10670
box -12 -8 32 272
use FILL  FILL_0__3381_
timestamp 1701859473
transform -1 0 6630 0 1 10670
box -12 -8 32 272
use FILL  FILL_0__3382_
timestamp 1701859473
transform 1 0 6090 0 -1 10670
box -12 -8 32 272
use FILL  FILL_0__3383_
timestamp 1701859473
transform -1 0 6350 0 -1 10670
box -12 -8 32 272
use FILL  FILL_0__3384_
timestamp 1701859473
transform -1 0 6790 0 -1 10670
box -12 -8 32 272
use FILL  FILL_0__3385_
timestamp 1701859473
transform 1 0 6550 0 -1 10670
box -12 -8 32 272
use FILL  FILL_0__3386_
timestamp 1701859473
transform 1 0 7030 0 -1 10670
box -12 -8 32 272
use FILL  FILL_0__3387_
timestamp 1701859473
transform 1 0 8390 0 -1 10670
box -12 -8 32 272
use FILL  FILL_0__3388_
timestamp 1701859473
transform 1 0 8510 0 1 10670
box -12 -8 32 272
use FILL  FILL_0__3389_
timestamp 1701859473
transform 1 0 10170 0 -1 10670
box -12 -8 32 272
use FILL  FILL_0__3390_
timestamp 1701859473
transform 1 0 9730 0 -1 10670
box -12 -8 32 272
use FILL  FILL_0__3391_
timestamp 1701859473
transform 1 0 9930 0 -1 10670
box -12 -8 32 272
use FILL  FILL_0__3392_
timestamp 1701859473
transform 1 0 10390 0 -1 10670
box -12 -8 32 272
use FILL  FILL_0__3393_
timestamp 1701859473
transform -1 0 11130 0 -1 10150
box -12 -8 32 272
use FILL  FILL_0__3394_
timestamp 1701859473
transform 1 0 7310 0 1 10150
box -12 -8 32 272
use FILL  FILL_0__3395_
timestamp 1701859473
transform 1 0 6370 0 1 10150
box -12 -8 32 272
use FILL  FILL_0__3396_
timestamp 1701859473
transform -1 0 6630 0 1 10150
box -12 -8 32 272
use FILL  FILL_0__3397_
timestamp 1701859473
transform -1 0 6950 0 -1 10150
box -12 -8 32 272
use FILL  FILL_0__3398_
timestamp 1701859473
transform 1 0 6230 0 -1 10150
box -12 -8 32 272
use FILL  FILL_0__3399_
timestamp 1701859473
transform -1 0 6710 0 -1 10150
box -12 -8 32 272
use FILL  FILL_0__3400_
timestamp 1701859473
transform -1 0 6890 0 1 10150
box -12 -8 32 272
use FILL  FILL_0__3401_
timestamp 1701859473
transform 1 0 7070 0 1 10150
box -12 -8 32 272
use FILL  FILL_0__3402_
timestamp 1701859473
transform -1 0 9010 0 1 10150
box -12 -8 32 272
use FILL  FILL_0__3403_
timestamp 1701859473
transform 1 0 9450 0 1 10150
box -12 -8 32 272
use FILL  FILL_0__3404_
timestamp 1701859473
transform -1 0 5710 0 1 9630
box -12 -8 32 272
use FILL  FILL_0__3405_
timestamp 1701859473
transform -1 0 5990 0 -1 10150
box -12 -8 32 272
use FILL  FILL_0__3406_
timestamp 1701859473
transform 1 0 6350 0 -1 9630
box -12 -8 32 272
use FILL  FILL_0__3407_
timestamp 1701859473
transform -1 0 6570 0 -1 9630
box -12 -8 32 272
use FILL  FILL_0__3408_
timestamp 1701859473
transform 1 0 6830 0 1 9630
box -12 -8 32 272
use FILL  FILL_0__3409_
timestamp 1701859473
transform -1 0 6450 0 -1 10150
box -12 -8 32 272
use FILL  FILL_0__3410_
timestamp 1701859473
transform 1 0 9190 0 -1 10150
box -12 -8 32 272
use FILL  FILL_0__3411_
timestamp 1701859473
transform 1 0 9210 0 1 10150
box -12 -8 32 272
use FILL  FILL_0__3412_
timestamp 1701859473
transform 1 0 9930 0 1 10150
box -12 -8 32 272
use FILL  FILL_0__3413_
timestamp 1701859473
transform -1 0 5950 0 1 9630
box -12 -8 32 272
use FILL  FILL_0__3414_
timestamp 1701859473
transform 1 0 8090 0 1 9110
box -12 -8 32 272
use FILL  FILL_0__3415_
timestamp 1701859473
transform 1 0 6370 0 1 9630
box -12 -8 32 272
use FILL  FILL_0__3416_
timestamp 1701859473
transform 1 0 7210 0 1 8590
box -12 -8 32 272
use FILL  FILL_0__3417_
timestamp 1701859473
transform 1 0 7290 0 -1 9110
box -12 -8 32 272
use FILL  FILL_0__3418_
timestamp 1701859473
transform -1 0 7430 0 -1 9630
box -12 -8 32 272
use FILL  FILL_0__3419_
timestamp 1701859473
transform 1 0 7190 0 -1 9630
box -12 -8 32 272
use FILL  FILL_0__3420_
timestamp 1701859473
transform -1 0 6770 0 -1 9630
box -12 -8 32 272
use FILL  FILL_0__3421_
timestamp 1701859473
transform -1 0 6990 0 -1 9630
box -12 -8 32 272
use FILL  FILL_0__3422_
timestamp 1701859473
transform -1 0 7090 0 1 9630
box -12 -8 32 272
use FILL  FILL_0__3423_
timestamp 1701859473
transform -1 0 8150 0 -1 9630
box -12 -8 32 272
use FILL  FILL_0__3424_
timestamp 1701859473
transform -1 0 7670 0 -1 9630
box -12 -8 32 272
use FILL  FILL_0__3425_
timestamp 1701859473
transform -1 0 7330 0 1 9630
box -12 -8 32 272
use FILL  FILL_0__3426_
timestamp 1701859473
transform -1 0 8970 0 -1 10150
box -12 -8 32 272
use FILL  FILL_0__3427_
timestamp 1701859473
transform 1 0 8730 0 -1 10150
box -12 -8 32 272
use FILL  FILL_0__3428_
timestamp 1701859473
transform 1 0 7410 0 1 8590
box -12 -8 32 272
use FILL  FILL_0__3429_
timestamp 1701859473
transform 1 0 7490 0 -1 9110
box -12 -8 32 272
use FILL  FILL_0__3430_
timestamp 1701859473
transform -1 0 7710 0 -1 9110
box -12 -8 32 272
use FILL  FILL_0__3431_
timestamp 1701859473
transform 1 0 7630 0 1 9110
box -12 -8 32 272
use FILL  FILL_0__3432_
timestamp 1701859473
transform 1 0 7870 0 1 9110
box -12 -8 32 272
use FILL  FILL_0__3433_
timestamp 1701859473
transform -1 0 7910 0 -1 9630
box -12 -8 32 272
use FILL  FILL_0__3434_
timestamp 1701859473
transform 1 0 7550 0 1 9630
box -12 -8 32 272
use FILL  FILL_0__3435_
timestamp 1701859473
transform 1 0 10170 0 1 10150
box -12 -8 32 272
use FILL  FILL_0__3436_
timestamp 1701859473
transform -1 0 10170 0 -1 10150
box -12 -8 32 272
use FILL  FILL_0__3437_
timestamp 1701859473
transform 1 0 10610 0 1 10150
box -12 -8 32 272
use FILL  FILL_0__3438_
timestamp 1701859473
transform 1 0 10390 0 1 10150
box -12 -8 32 272
use FILL  FILL_0__3439_
timestamp 1701859473
transform 1 0 10830 0 1 10150
box -12 -8 32 272
use FILL  FILL_0__3440_
timestamp 1701859473
transform -1 0 10650 0 -1 10150
box -12 -8 32 272
use FILL  FILL_0__3441_
timestamp 1701859473
transform -1 0 10510 0 1 9630
box -12 -8 32 272
use FILL  FILL_0__3442_
timestamp 1701859473
transform -1 0 10390 0 -1 10150
box -12 -8 32 272
use FILL  FILL_0__3443_
timestamp 1701859473
transform -1 0 10950 0 1 9630
box -12 -8 32 272
use FILL  FILL_0__3444_
timestamp 1701859473
transform -1 0 8350 0 -1 9630
box -12 -8 32 272
use FILL  FILL_0__3445_
timestamp 1701859473
transform -1 0 8050 0 1 9630
box -12 -8 32 272
use FILL  FILL_0__3446_
timestamp 1701859473
transform 1 0 8490 0 1 9630
box -12 -8 32 272
use FILL  FILL_0__3447_
timestamp 1701859473
transform 1 0 8270 0 1 9630
box -12 -8 32 272
use FILL  FILL_0__3448_
timestamp 1701859473
transform -1 0 8710 0 1 9630
box -12 -8 32 272
use FILL  FILL_0__3449_
timestamp 1701859473
transform -1 0 9750 0 1 10150
box -12 -8 32 272
use FILL  FILL_0__3450_
timestamp 1701859473
transform -1 0 9710 0 -1 10150
box -12 -8 32 272
use FILL  FILL_0__3451_
timestamp 1701859473
transform 1 0 9430 0 -1 10150
box -12 -8 32 272
use FILL  FILL_0__3452_
timestamp 1701859473
transform -1 0 9170 0 1 9630
box -12 -8 32 272
use FILL  FILL_0__3453_
timestamp 1701859473
transform -1 0 9930 0 -1 10150
box -12 -8 32 272
use FILL  FILL_0__3454_
timestamp 1701859473
transform 1 0 9370 0 1 9630
box -12 -8 32 272
use FILL  FILL_0__3455_
timestamp 1701859473
transform 1 0 9590 0 1 9630
box -12 -8 32 272
use FILL  FILL_0__3456_
timestamp 1701859473
transform -1 0 10290 0 1 9630
box -12 -8 32 272
use FILL  FILL_0__3457_
timestamp 1701859473
transform -1 0 9830 0 1 9630
box -12 -8 32 272
use FILL  FILL_0__3458_
timestamp 1701859473
transform -1 0 10070 0 1 9630
box -12 -8 32 272
use FILL  FILL_0__3459_
timestamp 1701859473
transform -1 0 10210 0 -1 9630
box -12 -8 32 272
use FILL  FILL_0__3460_
timestamp 1701859473
transform 1 0 10870 0 -1 10150
box -12 -8 32 272
use FILL  FILL_0__3461_
timestamp 1701859473
transform -1 0 11110 0 -1 9630
box -12 -8 32 272
use FILL  FILL_0__3462_
timestamp 1701859473
transform -1 0 10650 0 -1 9630
box -12 -8 32 272
use FILL  FILL_0__3463_
timestamp 1701859473
transform 1 0 10330 0 -1 11190
box -12 -8 32 272
use FILL  FILL_0__3464_
timestamp 1701859473
transform 1 0 9670 0 -1 11190
box -12 -8 32 272
use FILL  FILL_0__3465_
timestamp 1701859473
transform 1 0 9910 0 -1 11190
box -12 -8 32 272
use FILL  FILL_0__3466_
timestamp 1701859473
transform 1 0 10090 0 -1 11190
box -12 -8 32 272
use FILL  FILL_0__3467_
timestamp 1701859473
transform -1 0 11070 0 1 10670
box -12 -8 32 272
use FILL  FILL_0__3468_
timestamp 1701859473
transform 1 0 10570 0 1 10670
box -12 -8 32 272
use FILL  FILL_0__3469_
timestamp 1701859473
transform 1 0 9290 0 -1 10670
box -12 -8 32 272
use FILL  FILL_0__3470_
timestamp 1701859473
transform 1 0 9530 0 -1 10670
box -12 -8 32 272
use FILL  FILL_0__3471_
timestamp 1701859473
transform 1 0 9670 0 1 10670
box -12 -8 32 272
use FILL  FILL_0__3472_
timestamp 1701859473
transform -1 0 9930 0 1 10670
box -12 -8 32 272
use FILL  FILL_0__3473_
timestamp 1701859473
transform 1 0 8550 0 -1 11190
box -12 -8 32 272
use FILL  FILL_0__3474_
timestamp 1701859473
transform 1 0 8110 0 -1 11190
box -12 -8 32 272
use FILL  FILL_0__3475_
timestamp 1701859473
transform 1 0 8350 0 -1 11190
box -12 -8 32 272
use FILL  FILL_0__3476_
timestamp 1701859473
transform -1 0 8790 0 -1 11190
box -12 -8 32 272
use FILL  FILL_0__3477_
timestamp 1701859473
transform 1 0 9010 0 -1 11190
box -12 -8 32 272
use FILL  FILL_0__3478_
timestamp 1701859473
transform 1 0 8990 0 1 10670
box -12 -8 32 272
use FILL  FILL_0__3479_
timestamp 1701859473
transform 1 0 8270 0 -1 10150
box -12 -8 32 272
use FILL  FILL_0__3480_
timestamp 1701859473
transform -1 0 8530 0 -1 10150
box -12 -8 32 272
use FILL  FILL_0__3481_
timestamp 1701859473
transform -1 0 8310 0 1 9110
box -12 -8 32 272
use FILL  FILL_0__3482_
timestamp 1701859473
transform -1 0 8530 0 1 9110
box -12 -8 32 272
use FILL  FILL_0__3483_
timestamp 1701859473
transform 1 0 8710 0 1 10150
box -12 -8 32 272
use FILL  FILL_0__3484_
timestamp 1701859473
transform -1 0 10010 0 -1 9630
box -12 -8 32 272
use FILL  FILL_0__3485_
timestamp 1701859473
transform 1 0 11030 0 1 10150
box -12 -8 32 272
use FILL  FILL_0__3486_
timestamp 1701859473
transform 1 0 10370 0 1 9110
box -12 -8 32 272
use FILL  FILL_0__3487_
timestamp 1701859473
transform 1 0 10410 0 -1 9630
box -12 -8 32 272
use FILL  FILL_0__3488_
timestamp 1701859473
transform -1 0 10710 0 1 9630
box -12 -8 32 272
use FILL  FILL_0__3489_
timestamp 1701859473
transform 1 0 10550 0 -1 11190
box -12 -8 32 272
use FILL  FILL_0__3490_
timestamp 1701859473
transform 1 0 11010 0 -1 11190
box -12 -8 32 272
use FILL  FILL_0__3491_
timestamp 1701859473
transform -1 0 10810 0 -1 11190
box -12 -8 32 272
use FILL  FILL_0__3492_
timestamp 1701859473
transform -1 0 10370 0 1 10670
box -12 -8 32 272
use FILL  FILL_0__3493_
timestamp 1701859473
transform -1 0 10150 0 1 10670
box -12 -8 32 272
use FILL  FILL_0__3494_
timestamp 1701859473
transform 1 0 9250 0 1 10670
box -12 -8 32 272
use FILL  FILL_0__3495_
timestamp 1701859473
transform -1 0 9450 0 -1 11190
box -12 -8 32 272
use FILL  FILL_0__3496_
timestamp 1701859473
transform 1 0 9210 0 -1 11190
box -12 -8 32 272
use FILL  FILL_0__3497_
timestamp 1701859473
transform -1 0 9310 0 -1 9630
box -12 -8 32 272
use FILL  FILL_0__3498_
timestamp 1701859473
transform -1 0 8810 0 1 9110
box -12 -8 32 272
use FILL  FILL_0__3499_
timestamp 1701859473
transform 1 0 8330 0 -1 9110
box -12 -8 32 272
use FILL  FILL_0__3500_
timestamp 1701859473
transform 1 0 9710 0 1 9110
box -12 -8 32 272
use FILL  FILL_0__3501_
timestamp 1701859473
transform -1 0 9950 0 1 9110
box -12 -8 32 272
use FILL  FILL_0__3502_
timestamp 1701859473
transform -1 0 8210 0 -1 8590
box -12 -8 32 272
use FILL  FILL_0__3503_
timestamp 1701859473
transform -1 0 8590 0 -1 9630
box -12 -8 32 272
use FILL  FILL_0__3504_
timestamp 1701859473
transform 1 0 8810 0 -1 9630
box -12 -8 32 272
use FILL  FILL_0__3505_
timestamp 1701859473
transform -1 0 9070 0 -1 9630
box -12 -8 32 272
use FILL  FILL_0__3506_
timestamp 1701859473
transform -1 0 8590 0 1 8590
box -12 -8 32 272
use FILL  FILL_0__3507_
timestamp 1701859473
transform 1 0 10670 0 -1 9110
box -12 -8 32 272
use FILL  FILL_0__3508_
timestamp 1701859473
transform 1 0 10430 0 -1 9110
box -12 -8 32 272
use FILL  FILL_0__3509_
timestamp 1701859473
transform 1 0 8370 0 1 8590
box -12 -8 32 272
use FILL  FILL_0__3510_
timestamp 1701859473
transform -1 0 8830 0 1 8590
box -12 -8 32 272
use FILL  FILL_0__3511_
timestamp 1701859473
transform 1 0 9890 0 -1 270
box -12 -8 32 272
use FILL  FILL_0__3512_
timestamp 1701859473
transform 1 0 10890 0 -1 9110
box -12 -8 32 272
use FILL  FILL_0__3513_
timestamp 1701859473
transform 1 0 10870 0 -1 9630
box -12 -8 32 272
use FILL  FILL_0__3514_
timestamp 1701859473
transform 1 0 10830 0 1 10670
box -12 -8 32 272
use FILL  FILL_0__3515_
timestamp 1701859473
transform -1 0 10630 0 -1 10670
box -12 -8 32 272
use FILL  FILL_0__3516_
timestamp 1701859473
transform 1 0 10850 0 -1 10670
box -12 -8 32 272
use FILL  FILL_0__3517_
timestamp 1701859473
transform 1 0 9530 0 -1 9630
box -12 -8 32 272
use FILL  FILL_0__3518_
timestamp 1701859473
transform 1 0 9750 0 -1 9630
box -12 -8 32 272
use FILL  FILL_0__3519_
timestamp 1701859473
transform 1 0 9030 0 1 9110
box -12 -8 32 272
use FILL  FILL_0__3520_
timestamp 1701859473
transform -1 0 9270 0 1 9110
box -12 -8 32 272
use FILL  FILL_0__3521_
timestamp 1701859473
transform 1 0 6510 0 1 8590
box -12 -8 32 272
use FILL  FILL_0__3522_
timestamp 1701859473
transform 1 0 7910 0 -1 9110
box -12 -8 32 272
use FILL  FILL_0__3523_
timestamp 1701859473
transform 1 0 6710 0 1 8590
box -12 -8 32 272
use FILL  FILL_0__3524_
timestamp 1701859473
transform 1 0 7430 0 1 9110
box -12 -8 32 272
use FILL  FILL_0__3525_
timestamp 1701859473
transform 1 0 6970 0 1 9110
box -12 -8 32 272
use FILL  FILL_0__3526_
timestamp 1701859473
transform -1 0 7210 0 1 9110
box -12 -8 32 272
use FILL  FILL_0__3539_
timestamp 1701859473
transform 1 0 11070 0 -1 7030
box -12 -8 32 272
use FILL  FILL_0__3540_
timestamp 1701859473
transform 1 0 4570 0 1 10670
box -12 -8 32 272
use FILL  FILL_0__3541_
timestamp 1701859473
transform -1 0 30 0 1 5990
box -12 -8 32 272
use FILL  FILL_0__3542_
timestamp 1701859473
transform -1 0 30 0 -1 8070
box -12 -8 32 272
use FILL  FILL_0__3543_
timestamp 1701859473
transform -1 0 30 0 1 8590
box -12 -8 32 272
use FILL  FILL_0__3544_
timestamp 1701859473
transform -1 0 30 0 1 9110
box -12 -8 32 272
use FILL  FILL_0__3545_
timestamp 1701859473
transform -1 0 1870 0 -1 11190
box -12 -8 32 272
use FILL  FILL_0__3546_
timestamp 1701859473
transform -1 0 490 0 1 9110
box -12 -8 32 272
use FILL  FILL_0__3547_
timestamp 1701859473
transform 1 0 4610 0 -1 11190
box -12 -8 32 272
use FILL  FILL_0__3548_
timestamp 1701859473
transform 1 0 5210 0 1 10670
box -12 -8 32 272
use FILL  FILL_0__3549_
timestamp 1701859473
transform -1 0 4210 0 -1 11190
box -12 -8 32 272
use FILL  FILL_0__3550_
timestamp 1701859473
transform -1 0 5050 0 -1 11190
box -12 -8 32 272
use FILL  FILL_0__3551_
timestamp 1701859473
transform 1 0 5450 0 -1 11190
box -12 -8 32 272
use FILL  FILL_0__3552_
timestamp 1701859473
transform 1 0 5230 0 -1 11190
box -12 -8 32 272
use FILL  FILL_0__3553_
timestamp 1701859473
transform -1 0 30 0 -1 5990
box -12 -8 32 272
use FILL  FILL_0__3554_
timestamp 1701859473
transform -1 0 230 0 1 7030
box -12 -8 32 272
use FILL  FILL_0__3555_
timestamp 1701859473
transform -1 0 5010 0 1 10670
box -12 -8 32 272
use FILL  FILL_0__3556_
timestamp 1701859473
transform 1 0 6150 0 1 10150
box -12 -8 32 272
use FILL  FILL_0__3557_
timestamp 1701859473
transform -1 0 5690 0 -1 11190
box -12 -8 32 272
use FILL  FILL_0__3558_
timestamp 1701859473
transform 1 0 6090 0 -1 11190
box -12 -8 32 272
use FILL  FILL_0__3559_
timestamp 1701859473
transform -1 0 4750 0 -1 10670
box -12 -8 32 272
use FILL  FILL_0__3560_
timestamp 1701859473
transform 1 0 5430 0 1 10670
box -12 -8 32 272
use FILL  FILL_0__3561_
timestamp 1701859473
transform 1 0 5870 0 -1 11190
box -12 -8 32 272
use FILL  FILL_0__3562_
timestamp 1701859473
transform 1 0 5670 0 1 10150
box -12 -8 32 272
use FILL  FILL_0__3563_
timestamp 1701859473
transform 1 0 5130 0 1 3390
box -12 -8 32 272
use FILL  FILL_0_BUFX2_insert0
timestamp 1701859473
transform 1 0 5750 0 -1 10150
box -12 -8 32 272
use FILL  FILL_0_BUFX2_insert1
timestamp 1701859473
transform 1 0 6510 0 1 2350
box -12 -8 32 272
use FILL  FILL_0_BUFX2_insert2
timestamp 1701859473
transform 1 0 5350 0 -1 1830
box -12 -8 32 272
use FILL  FILL_0_BUFX2_insert3
timestamp 1701859473
transform -1 0 490 0 -1 5470
box -12 -8 32 272
use FILL  FILL_0_BUFX2_insert4
timestamp 1701859473
transform 1 0 3230 0 1 4950
box -12 -8 32 272
use FILL  FILL_0_BUFX2_insert5
timestamp 1701859473
transform 1 0 1290 0 -1 1830
box -12 -8 32 272
use FILL  FILL_0_BUFX2_insert6
timestamp 1701859473
transform -1 0 30 0 -1 11190
box -12 -8 32 272
use FILL  FILL_0_BUFX2_insert7
timestamp 1701859473
transform 1 0 1590 0 1 10670
box -12 -8 32 272
use FILL  FILL_0_BUFX2_insert8
timestamp 1701859473
transform 1 0 1550 0 1 1830
box -12 -8 32 272
use FILL  FILL_0_BUFX2_insert9
timestamp 1701859473
transform 1 0 1850 0 -1 3910
box -12 -8 32 272
use FILL  FILL_0_BUFX2_insert10
timestamp 1701859473
transform 1 0 1670 0 -1 4430
box -12 -8 32 272
use FILL  FILL_0_BUFX2_insert11
timestamp 1701859473
transform -1 0 1650 0 -1 3910
box -12 -8 32 272
use FILL  FILL_0_BUFX2_insert12
timestamp 1701859473
transform -1 0 1430 0 -1 3910
box -12 -8 32 272
use FILL  FILL_0_BUFX2_insert13
timestamp 1701859473
transform -1 0 1330 0 -1 1310
box -12 -8 32 272
use FILL  FILL_0_BUFX2_insert14
timestamp 1701859473
transform -1 0 3570 0 1 3390
box -12 -8 32 272
use FILL  FILL_0_BUFX2_insert15
timestamp 1701859473
transform 1 0 4450 0 -1 5470
box -12 -8 32 272
use FILL  FILL_0_BUFX2_insert16
timestamp 1701859473
transform 1 0 1250 0 -1 4950
box -12 -8 32 272
use FILL  FILL_0_BUFX2_insert17
timestamp 1701859473
transform 1 0 3530 0 1 1310
box -12 -8 32 272
use FILL  FILL_0_BUFX2_insert18
timestamp 1701859473
transform -1 0 9670 0 1 2350
box -12 -8 32 272
use FILL  FILL_0_BUFX2_insert19
timestamp 1701859473
transform -1 0 8410 0 -1 790
box -12 -8 32 272
use FILL  FILL_0_BUFX2_insert20
timestamp 1701859473
transform 1 0 9870 0 1 2350
box -12 -8 32 272
use FILL  FILL_0_BUFX2_insert21
timestamp 1701859473
transform -1 0 7710 0 -1 1310
box -12 -8 32 272
use FILL  FILL_0_BUFX2_insert22
timestamp 1701859473
transform -1 0 3110 0 -1 2870
box -12 -8 32 272
use FILL  FILL_0_BUFX2_insert23
timestamp 1701859473
transform -1 0 2650 0 -1 4950
box -12 -8 32 272
use FILL  FILL_0_BUFX2_insert24
timestamp 1701859473
transform -1 0 3550 0 -1 4430
box -12 -8 32 272
use FILL  FILL_0_BUFX2_insert25
timestamp 1701859473
transform 1 0 4290 0 1 4430
box -12 -8 32 272
use FILL  FILL_0_BUFX2_insert26
timestamp 1701859473
transform 1 0 4110 0 1 2870
box -12 -8 32 272
use FILL  FILL_0_BUFX2_insert27
timestamp 1701859473
transform 1 0 9510 0 1 4950
box -12 -8 32 272
use FILL  FILL_0_BUFX2_insert28
timestamp 1701859473
transform -1 0 7390 0 -1 5990
box -12 -8 32 272
use FILL  FILL_0_BUFX2_insert29
timestamp 1701859473
transform -1 0 1190 0 1 6510
box -12 -8 32 272
use FILL  FILL_0_BUFX2_insert30
timestamp 1701859473
transform -1 0 8690 0 -1 3910
box -12 -8 32 272
use FILL  FILL_0_BUFX2_insert31
timestamp 1701859473
transform -1 0 9470 0 1 3910
box -12 -8 32 272
use FILL  FILL_0_BUFX2_insert32
timestamp 1701859473
transform 1 0 5770 0 -1 3910
box -12 -8 32 272
use FILL  FILL_0_BUFX2_insert33
timestamp 1701859473
transform -1 0 9450 0 -1 4950
box -12 -8 32 272
use FILL  FILL_0_BUFX2_insert34
timestamp 1701859473
transform 1 0 5110 0 1 8590
box -12 -8 32 272
use FILL  FILL_0_BUFX2_insert35
timestamp 1701859473
transform -1 0 5870 0 1 7550
box -12 -8 32 272
use FILL  FILL_0_BUFX2_insert36
timestamp 1701859473
transform -1 0 1110 0 1 8590
box -12 -8 32 272
use FILL  FILL_0_BUFX2_insert37
timestamp 1701859473
transform -1 0 9490 0 1 8590
box -12 -8 32 272
use FILL  FILL_0_BUFX2_insert49
timestamp 1701859473
transform -1 0 2950 0 1 6510
box -12 -8 32 272
use FILL  FILL_0_BUFX2_insert50
timestamp 1701859473
transform 1 0 2250 0 -1 8590
box -12 -8 32 272
use FILL  FILL_0_BUFX2_insert51
timestamp 1701859473
transform 1 0 3110 0 -1 8590
box -12 -8 32 272
use FILL  FILL_0_BUFX2_insert52
timestamp 1701859473
transform 1 0 3290 0 1 5470
box -12 -8 32 272
use FILL  FILL_0_BUFX2_insert53
timestamp 1701859473
transform -1 0 11130 0 1 9110
box -12 -8 32 272
use FILL  FILL_0_BUFX2_insert54
timestamp 1701859473
transform -1 0 9070 0 1 8590
box -12 -8 32 272
use FILL  FILL_0_BUFX2_insert55
timestamp 1701859473
transform -1 0 9510 0 1 9110
box -12 -8 32 272
use FILL  FILL_0_BUFX2_insert56
timestamp 1701859473
transform -1 0 10170 0 1 9110
box -12 -8 32 272
use FILL  FILL_0_BUFX2_insert57
timestamp 1701859473
transform -1 0 11130 0 -1 2350
box -12 -8 32 272
use FILL  FILL_0_BUFX2_insert58
timestamp 1701859473
transform -1 0 8870 0 1 2870
box -12 -8 32 272
use FILL  FILL_0_BUFX2_insert59
timestamp 1701859473
transform -1 0 7450 0 1 1830
box -12 -8 32 272
use FILL  FILL_0_BUFX2_insert60
timestamp 1701859473
transform 1 0 10790 0 1 1830
box -12 -8 32 272
use FILL  FILL_0_BUFX2_insert61
timestamp 1701859473
transform -1 0 11070 0 1 2870
box -12 -8 32 272
use FILL  FILL_0_BUFX2_insert62
timestamp 1701859473
transform 1 0 2110 0 1 3910
box -12 -8 32 272
use FILL  FILL_0_BUFX2_insert63
timestamp 1701859473
transform 1 0 2030 0 1 3390
box -12 -8 32 272
use FILL  FILL_0_BUFX2_insert64
timestamp 1701859473
transform -1 0 1690 0 1 3910
box -12 -8 32 272
use FILL  FILL_0_BUFX2_insert65
timestamp 1701859473
transform -1 0 1630 0 1 3390
box -12 -8 32 272
use FILL  FILL_0_BUFX2_insert66
timestamp 1701859473
transform -1 0 4210 0 1 1310
box -12 -8 32 272
use FILL  FILL_0_BUFX2_insert67
timestamp 1701859473
transform -1 0 3510 0 -1 10150
box -12 -8 32 272
use FILL  FILL_0_BUFX2_insert68
timestamp 1701859473
transform -1 0 7070 0 1 2870
box -12 -8 32 272
use FILL  FILL_0_BUFX2_insert69
timestamp 1701859473
transform -1 0 5550 0 -1 3390
box -12 -8 32 272
use FILL  FILL_0_BUFX2_insert70
timestamp 1701859473
transform -1 0 3570 0 -1 1830
box -12 -8 32 272
use FILL  FILL_0_BUFX2_insert71
timestamp 1701859473
transform -1 0 7210 0 1 2350
box -12 -8 32 272
use FILL  FILL_0_BUFX2_insert72
timestamp 1701859473
transform -1 0 6390 0 1 1310
box -12 -8 32 272
use FILL  FILL_0_BUFX2_insert73
timestamp 1701859473
transform 1 0 3510 0 1 5470
box -12 -8 32 272
use FILL  FILL_0_BUFX2_insert74
timestamp 1701859473
transform 1 0 7470 0 -1 2350
box -12 -8 32 272
use FILL  FILL_0_BUFX2_insert75
timestamp 1701859473
transform 1 0 7490 0 1 2870
box -12 -8 32 272
use FILL  FILL_0_BUFX2_insert76
timestamp 1701859473
transform 1 0 7270 0 1 2870
box -12 -8 32 272
use FILL  FILL_0_BUFX2_insert77
timestamp 1701859473
transform -1 0 3330 0 -1 2870
box -12 -8 32 272
use FILL  FILL_0_BUFX2_insert78
timestamp 1701859473
transform 1 0 1830 0 -1 2870
box -12 -8 32 272
use FILL  FILL_0_BUFX2_insert79
timestamp 1701859473
transform -1 0 2070 0 -1 2870
box -12 -8 32 272
use FILL  FILL_0_BUFX2_insert80
timestamp 1701859473
transform 1 0 2310 0 1 4430
box -12 -8 32 272
use FILL  FILL_0_BUFX2_insert81
timestamp 1701859473
transform -1 0 1910 0 1 3910
box -12 -8 32 272
use FILL  FILL_0_BUFX2_insert82
timestamp 1701859473
transform -1 0 230 0 1 8590
box -12 -8 32 272
use FILL  FILL_0_BUFX2_insert83
timestamp 1701859473
transform 1 0 4110 0 -1 10150
box -12 -8 32 272
use FILL  FILL_0_BUFX2_insert84
timestamp 1701859473
transform 1 0 4070 0 -1 7550
box -12 -8 32 272
use FILL  FILL_0_BUFX2_insert85
timestamp 1701859473
transform -1 0 30 0 -1 6510
box -12 -8 32 272
use FILL  FILL_0_BUFX2_insert86
timestamp 1701859473
transform 1 0 1830 0 -1 10150
box -12 -8 32 272
use FILL  FILL_0_CLKBUF1_insert38
timestamp 1701859473
transform 1 0 2830 0 -1 7550
box -12 -8 32 272
use FILL  FILL_0_CLKBUF1_insert39
timestamp 1701859473
transform -1 0 4630 0 -1 6510
box -12 -8 32 272
use FILL  FILL_0_CLKBUF1_insert40
timestamp 1701859473
transform -1 0 930 0 -1 4950
box -12 -8 32 272
use FILL  FILL_0_CLKBUF1_insert41
timestamp 1701859473
transform -1 0 10590 0 -1 270
box -12 -8 32 272
use FILL  FILL_0_CLKBUF1_insert42
timestamp 1701859473
transform 1 0 9650 0 -1 4950
box -12 -8 32 272
use FILL  FILL_0_CLKBUF1_insert43
timestamp 1701859473
transform -1 0 10970 0 1 7030
box -12 -8 32 272
use FILL  FILL_0_CLKBUF1_insert44
timestamp 1701859473
transform -1 0 10710 0 1 4430
box -12 -8 32 272
use FILL  FILL_0_CLKBUF1_insert45
timestamp 1701859473
transform 1 0 5630 0 -1 6510
box -12 -8 32 272
use FILL  FILL_0_CLKBUF1_insert46
timestamp 1701859473
transform 1 0 3950 0 1 5990
box -12 -8 32 272
use FILL  FILL_0_CLKBUF1_insert47
timestamp 1701859473
transform -1 0 2070 0 1 7550
box -12 -8 32 272
use FILL  FILL_0_CLKBUF1_insert48
timestamp 1701859473
transform -1 0 10750 0 -1 7030
box -12 -8 32 272
use FILL  FILL_1__1668_
timestamp 1701859473
transform 1 0 6710 0 -1 3390
box -12 -8 32 272
use FILL  FILL_1__1669_
timestamp 1701859473
transform -1 0 6750 0 -1 790
box -12 -8 32 272
use FILL  FILL_1__1670_
timestamp 1701859473
transform 1 0 6530 0 -1 2870
box -12 -8 32 272
use FILL  FILL_1__1671_
timestamp 1701859473
transform -1 0 6330 0 -1 8590
box -12 -8 32 272
use FILL  FILL_1__1672_
timestamp 1701859473
transform 1 0 5890 0 -1 10670
box -12 -8 32 272
use FILL  FILL_1__1673_
timestamp 1701859473
transform 1 0 6290 0 1 8590
box -12 -8 32 272
use FILL  FILL_1__1674_
timestamp 1701859473
transform -1 0 6370 0 -1 9110
box -12 -8 32 272
use FILL  FILL_1__1675_
timestamp 1701859473
transform 1 0 30 0 -1 5470
box -12 -8 32 272
use FILL  FILL_1__1676_
timestamp 1701859473
transform -1 0 270 0 -1 5470
box -12 -8 32 272
use FILL  FILL_1__1677_
timestamp 1701859473
transform -1 0 510 0 1 5470
box -12 -8 32 272
use FILL  FILL_1__1678_
timestamp 1701859473
transform 1 0 30 0 -1 10670
box -12 -8 32 272
use FILL  FILL_1__1679_
timestamp 1701859473
transform -1 0 250 0 -1 11190
box -12 -8 32 272
use FILL  FILL_1__1680_
timestamp 1701859473
transform 1 0 230 0 -1 10670
box -12 -8 32 272
use FILL  FILL_1__1681_
timestamp 1701859473
transform -1 0 50 0 -1 7030
box -12 -8 32 272
use FILL  FILL_1__1682_
timestamp 1701859473
transform -1 0 50 0 1 7030
box -12 -8 32 272
use FILL  FILL_1__1683_
timestamp 1701859473
transform 1 0 30 0 1 6510
box -12 -8 32 272
use FILL  FILL_1__1684_
timestamp 1701859473
transform 1 0 910 0 -1 11190
box -12 -8 32 272
use FILL  FILL_1__1685_
timestamp 1701859473
transform -1 0 1170 0 -1 11190
box -12 -8 32 272
use FILL  FILL_1__1686_
timestamp 1701859473
transform -1 0 970 0 1 10670
box -12 -8 32 272
use FILL  FILL_1__1687_
timestamp 1701859473
transform 1 0 1390 0 -1 11190
box -12 -8 32 272
use FILL  FILL_1__1688_
timestamp 1701859473
transform -1 0 1650 0 -1 11190
box -12 -8 32 272
use FILL  FILL_1__1689_
timestamp 1701859473
transform -1 0 1910 0 1 10150
box -12 -8 32 272
use FILL  FILL_1__1690_
timestamp 1701859473
transform 1 0 2070 0 1 9110
box -12 -8 32 272
use FILL  FILL_1__1691_
timestamp 1701859473
transform -1 0 2090 0 -1 9110
box -12 -8 32 272
use FILL  FILL_1__1692_
timestamp 1701859473
transform 1 0 30 0 1 790
box -12 -8 32 272
use FILL  FILL_1__1693_
timestamp 1701859473
transform 1 0 30 0 -1 1310
box -12 -8 32 272
use FILL  FILL_1__1694_
timestamp 1701859473
transform 1 0 450 0 -1 270
box -12 -8 32 272
use FILL  FILL_1__1695_
timestamp 1701859473
transform -1 0 670 0 -1 270
box -12 -8 32 272
use FILL  FILL_1__1696_
timestamp 1701859473
transform 1 0 1090 0 1 2870
box -12 -8 32 272
use FILL  FILL_1__1697_
timestamp 1701859473
transform -1 0 2750 0 -1 2870
box -12 -8 32 272
use FILL  FILL_1__1698_
timestamp 1701859473
transform -1 0 1850 0 1 3390
box -12 -8 32 272
use FILL  FILL_1__1699_
timestamp 1701859473
transform 1 0 3770 0 1 3390
box -12 -8 32 272
use FILL  FILL_1__1700_
timestamp 1701859473
transform -1 0 2570 0 -1 3910
box -12 -8 32 272
use FILL  FILL_1__1701_
timestamp 1701859473
transform -1 0 1110 0 1 270
box -12 -8 32 272
use FILL  FILL_1__1702_
timestamp 1701859473
transform 1 0 870 0 1 270
box -12 -8 32 272
use FILL  FILL_1__1703_
timestamp 1701859473
transform -1 0 1350 0 1 1830
box -12 -8 32 272
use FILL  FILL_1__1704_
timestamp 1701859473
transform -1 0 9110 0 1 2870
box -12 -8 32 272
use FILL  FILL_1__1705_
timestamp 1701859473
transform 1 0 9730 0 -1 790
box -12 -8 32 272
use FILL  FILL_1__1706_
timestamp 1701859473
transform -1 0 7950 0 -1 4950
box -12 -8 32 272
use FILL  FILL_1__1707_
timestamp 1701859473
transform 1 0 8390 0 -1 4950
box -12 -8 32 272
use FILL  FILL_1__1708_
timestamp 1701859473
transform 1 0 5010 0 -1 5990
box -12 -8 32 272
use FILL  FILL_1__1709_
timestamp 1701859473
transform -1 0 11110 0 1 5990
box -12 -8 32 272
use FILL  FILL_1__1710_
timestamp 1701859473
transform 1 0 5390 0 -1 5470
box -12 -8 32 272
use FILL  FILL_1__1711_
timestamp 1701859473
transform -1 0 5230 0 -1 5990
box -12 -8 32 272
use FILL  FILL_1__1712_
timestamp 1701859473
transform -1 0 5050 0 1 5470
box -12 -8 32 272
use FILL  FILL_1__1713_
timestamp 1701859473
transform 1 0 7910 0 1 4430
box -12 -8 32 272
use FILL  FILL_1__1714_
timestamp 1701859473
transform 1 0 7710 0 1 4950
box -12 -8 32 272
use FILL  FILL_1__1715_
timestamp 1701859473
transform -1 0 7950 0 1 4950
box -12 -8 32 272
use FILL  FILL_1__1716_
timestamp 1701859473
transform -1 0 8170 0 1 4430
box -12 -8 32 272
use FILL  FILL_1__1717_
timestamp 1701859473
transform -1 0 7950 0 1 1310
box -12 -8 32 272
use FILL  FILL_1__1718_
timestamp 1701859473
transform -1 0 5890 0 1 5990
box -12 -8 32 272
use FILL  FILL_1__1719_
timestamp 1701859473
transform -1 0 6750 0 -1 5990
box -12 -8 32 272
use FILL  FILL_1__1720_
timestamp 1701859473
transform -1 0 6730 0 1 5470
box -12 -8 32 272
use FILL  FILL_1__1721_
timestamp 1701859473
transform -1 0 6970 0 1 5470
box -12 -8 32 272
use FILL  FILL_1__1722_
timestamp 1701859473
transform -1 0 7670 0 1 4430
box -12 -8 32 272
use FILL  FILL_1__1723_
timestamp 1701859473
transform 1 0 7890 0 1 1830
box -12 -8 32 272
use FILL  FILL_1__1724_
timestamp 1701859473
transform -1 0 7930 0 -1 1310
box -12 -8 32 272
use FILL  FILL_1__1725_
timestamp 1701859473
transform 1 0 6530 0 1 5990
box -12 -8 32 272
use FILL  FILL_1__1726_
timestamp 1701859473
transform 1 0 6730 0 1 5990
box -12 -8 32 272
use FILL  FILL_1__1727_
timestamp 1701859473
transform -1 0 6970 0 1 5990
box -12 -8 32 272
use FILL  FILL_1__1728_
timestamp 1701859473
transform 1 0 7670 0 1 5990
box -12 -8 32 272
use FILL  FILL_1__1729_
timestamp 1701859473
transform -1 0 7610 0 -1 5990
box -12 -8 32 272
use FILL  FILL_1__1730_
timestamp 1701859473
transform -1 0 8090 0 1 3390
box -12 -8 32 272
use FILL  FILL_1__1731_
timestamp 1701859473
transform -1 0 7950 0 -1 270
box -12 -8 32 272
use FILL  FILL_1__1732_
timestamp 1701859473
transform -1 0 7910 0 1 5470
box -12 -8 32 272
use FILL  FILL_1__1733_
timestamp 1701859473
transform -1 0 8130 0 1 5470
box -12 -8 32 272
use FILL  FILL_1__1734_
timestamp 1701859473
transform 1 0 8090 0 -1 5470
box -12 -8 32 272
use FILL  FILL_1__1735_
timestamp 1701859473
transform 1 0 8550 0 -1 5470
box -12 -8 32 272
use FILL  FILL_1__1736_
timestamp 1701859473
transform 1 0 8390 0 1 4950
box -12 -8 32 272
use FILL  FILL_1__1737_
timestamp 1701859473
transform -1 0 8470 0 -1 3910
box -12 -8 32 272
use FILL  FILL_1__1738_
timestamp 1701859473
transform 1 0 8870 0 1 790
box -12 -8 32 272
use FILL  FILL_1__1739_
timestamp 1701859473
transform -1 0 9090 0 -1 790
box -12 -8 32 272
use FILL  FILL_1__1740_
timestamp 1701859473
transform 1 0 6450 0 1 270
box -12 -8 32 272
use FILL  FILL_1__1741_
timestamp 1701859473
transform 1 0 6350 0 1 790
box -12 -8 32 272
use FILL  FILL_1__1742_
timestamp 1701859473
transform -1 0 6290 0 -1 790
box -12 -8 32 272
use FILL  FILL_1__1743_
timestamp 1701859473
transform -1 0 2290 0 -1 3390
box -12 -8 32 272
use FILL  FILL_1__1744_
timestamp 1701859473
transform 1 0 270 0 -1 4950
box -12 -8 32 272
use FILL  FILL_1__1745_
timestamp 1701859473
transform 1 0 2090 0 -1 3910
box -12 -8 32 272
use FILL  FILL_1__1746_
timestamp 1701859473
transform -1 0 5110 0 -1 3390
box -12 -8 32 272
use FILL  FILL_1__1747_
timestamp 1701859473
transform -1 0 270 0 -1 270
box -12 -8 32 272
use FILL  FILL_1__1748_
timestamp 1701859473
transform -1 0 470 0 1 270
box -12 -8 32 272
use FILL  FILL_1__1749_
timestamp 1701859473
transform -1 0 910 0 1 1310
box -12 -8 32 272
use FILL  FILL_1__1750_
timestamp 1701859473
transform -1 0 1130 0 1 1310
box -12 -8 32 272
use FILL  FILL_1__1751_
timestamp 1701859473
transform -1 0 4490 0 -1 2870
box -12 -8 32 272
use FILL  FILL_1__1752_
timestamp 1701859473
transform 1 0 4690 0 -1 2870
box -12 -8 32 272
use FILL  FILL_1__1753_
timestamp 1701859473
transform -1 0 4310 0 1 790
box -12 -8 32 272
use FILL  FILL_1__1754_
timestamp 1701859473
transform 1 0 250 0 -1 790
box -12 -8 32 272
use FILL  FILL_1__1755_
timestamp 1701859473
transform -1 0 470 0 -1 790
box -12 -8 32 272
use FILL  FILL_1__1756_
timestamp 1701859473
transform -1 0 50 0 -1 270
box -12 -8 32 272
use FILL  FILL_1__1757_
timestamp 1701859473
transform 1 0 650 0 -1 790
box -12 -8 32 272
use FILL  FILL_1__1758_
timestamp 1701859473
transform 1 0 30 0 1 2350
box -12 -8 32 272
use FILL  FILL_1__1759_
timestamp 1701859473
transform -1 0 2530 0 -1 2870
box -12 -8 32 272
use FILL  FILL_1__1760_
timestamp 1701859473
transform 1 0 2910 0 -1 2870
box -12 -8 32 272
use FILL  FILL_1__1761_
timestamp 1701859473
transform -1 0 3230 0 -1 3390
box -12 -8 32 272
use FILL  FILL_1__1762_
timestamp 1701859473
transform -1 0 50 0 1 270
box -12 -8 32 272
use FILL  FILL_1__1763_
timestamp 1701859473
transform 1 0 30 0 -1 790
box -12 -8 32 272
use FILL  FILL_1__1764_
timestamp 1701859473
transform 1 0 470 0 1 1310
box -12 -8 32 272
use FILL  FILL_1__1765_
timestamp 1701859473
transform 1 0 1330 0 1 1310
box -12 -8 32 272
use FILL  FILL_1__1766_
timestamp 1701859473
transform -1 0 3130 0 -1 1830
box -12 -8 32 272
use FILL  FILL_1__1767_
timestamp 1701859473
transform 1 0 1430 0 -1 4430
box -12 -8 32 272
use FILL  FILL_1__1768_
timestamp 1701859473
transform 1 0 250 0 -1 1310
box -12 -8 32 272
use FILL  FILL_1__1769_
timestamp 1701859473
transform -1 0 470 0 1 1830
box -12 -8 32 272
use FILL  FILL_1__1770_
timestamp 1701859473
transform 1 0 2070 0 -1 3390
box -12 -8 32 272
use FILL  FILL_1__1771_
timestamp 1701859473
transform -1 0 2330 0 -1 3910
box -12 -8 32 272
use FILL  FILL_1__1772_
timestamp 1701859473
transform -1 0 2990 0 -1 3910
box -12 -8 32 272
use FILL  FILL_1__1773_
timestamp 1701859473
transform 1 0 3890 0 1 2870
box -12 -8 32 272
use FILL  FILL_1__1774_
timestamp 1701859473
transform -1 0 5270 0 -1 2350
box -12 -8 32 272
use FILL  FILL_1__1775_
timestamp 1701859473
transform 1 0 230 0 1 790
box -12 -8 32 272
use FILL  FILL_1__1776_
timestamp 1701859473
transform -1 0 270 0 1 1310
box -12 -8 32 272
use FILL  FILL_1__1777_
timestamp 1701859473
transform 1 0 690 0 -1 1830
box -12 -8 32 272
use FILL  FILL_1__1778_
timestamp 1701859473
transform -1 0 4410 0 1 5470
box -12 -8 32 272
use FILL  FILL_1__1779_
timestamp 1701859473
transform -1 0 6050 0 -1 5470
box -12 -8 32 272
use FILL  FILL_1__1780_
timestamp 1701859473
transform 1 0 4770 0 1 2870
box -12 -8 32 272
use FILL  FILL_1__1781_
timestamp 1701859473
transform 1 0 4350 0 1 2870
box -12 -8 32 272
use FILL  FILL_1__1782_
timestamp 1701859473
transform -1 0 50 0 1 1310
box -12 -8 32 272
use FILL  FILL_1__1783_
timestamp 1701859473
transform -1 0 1330 0 1 2870
box -12 -8 32 272
use FILL  FILL_1__1784_
timestamp 1701859473
transform -1 0 5030 0 1 2870
box -12 -8 32 272
use FILL  FILL_1__1785_
timestamp 1701859473
transform 1 0 4950 0 -1 2870
box -12 -8 32 272
use FILL  FILL_1__1786_
timestamp 1701859473
transform -1 0 5030 0 -1 2350
box -12 -8 32 272
use FILL  FILL_1__1787_
timestamp 1701859473
transform 1 0 5010 0 1 2350
box -12 -8 32 272
use FILL  FILL_1__1788_
timestamp 1701859473
transform -1 0 4810 0 -1 2350
box -12 -8 32 272
use FILL  FILL_1__1789_
timestamp 1701859473
transform 1 0 30 0 1 1830
box -12 -8 32 272
use FILL  FILL_1__1790_
timestamp 1701859473
transform -1 0 270 0 -1 2350
box -12 -8 32 272
use FILL  FILL_1__1791_
timestamp 1701859473
transform -1 0 2070 0 -1 2350
box -12 -8 32 272
use FILL  FILL_1__1792_
timestamp 1701859473
transform -1 0 3450 0 -1 2350
box -12 -8 32 272
use FILL  FILL_1__1793_
timestamp 1701859473
transform -1 0 4550 0 1 1830
box -12 -8 32 272
use FILL  FILL_1__1794_
timestamp 1701859473
transform 1 0 870 0 1 1830
box -12 -8 32 272
use FILL  FILL_1__1795_
timestamp 1701859473
transform -1 0 2130 0 1 2350
box -12 -8 32 272
use FILL  FILL_1__1796_
timestamp 1701859473
transform -1 0 1750 0 -1 1830
box -12 -8 32 272
use FILL  FILL_1__1797_
timestamp 1701859473
transform 1 0 1970 0 -1 1830
box -12 -8 32 272
use FILL  FILL_1__1798_
timestamp 1701859473
transform 1 0 890 0 -1 1310
box -12 -8 32 272
use FILL  FILL_1__1799_
timestamp 1701859473
transform 1 0 3710 0 1 3910
box -12 -8 32 272
use FILL  FILL_1__1800_
timestamp 1701859473
transform 1 0 3390 0 1 1830
box -12 -8 32 272
use FILL  FILL_1__1801_
timestamp 1701859473
transform -1 0 1130 0 1 1830
box -12 -8 32 272
use FILL  FILL_1__1802_
timestamp 1701859473
transform -1 0 3670 0 1 2350
box -12 -8 32 272
use FILL  FILL_1__1803_
timestamp 1701859473
transform -1 0 3890 0 1 2350
box -12 -8 32 272
use FILL  FILL_1__1804_
timestamp 1701859473
transform -1 0 4130 0 1 2350
box -12 -8 32 272
use FILL  FILL_1__1805_
timestamp 1701859473
transform 1 0 5430 0 1 2350
box -12 -8 32 272
use FILL  FILL_1__1806_
timestamp 1701859473
transform -1 0 4830 0 1 2350
box -12 -8 32 272
use FILL  FILL_1__1807_
timestamp 1701859473
transform -1 0 5230 0 1 2350
box -12 -8 32 272
use FILL  FILL_1__1808_
timestamp 1701859473
transform 1 0 4750 0 1 1830
box -12 -8 32 272
use FILL  FILL_1__1809_
timestamp 1701859473
transform -1 0 7110 0 -1 270
box -12 -8 32 272
use FILL  FILL_1__1810_
timestamp 1701859473
transform -1 0 7090 0 1 1310
box -12 -8 32 272
use FILL  FILL_1__1811_
timestamp 1701859473
transform 1 0 7430 0 -1 1830
box -12 -8 32 272
use FILL  FILL_1__1812_
timestamp 1701859473
transform -1 0 7510 0 -1 1310
box -12 -8 32 272
use FILL  FILL_1__1813_
timestamp 1701859473
transform 1 0 9090 0 1 790
box -12 -8 32 272
use FILL  FILL_1__1814_
timestamp 1701859473
transform -1 0 8130 0 -1 1830
box -12 -8 32 272
use FILL  FILL_1__1815_
timestamp 1701859473
transform 1 0 8330 0 1 2350
box -12 -8 32 272
use FILL  FILL_1__1816_
timestamp 1701859473
transform -1 0 9610 0 -1 2350
box -12 -8 32 272
use FILL  FILL_1__1817_
timestamp 1701859473
transform -1 0 9330 0 1 1310
box -12 -8 32 272
use FILL  FILL_1__1818_
timestamp 1701859473
transform -1 0 9530 0 1 270
box -12 -8 32 272
use FILL  FILL_1__1819_
timestamp 1701859473
transform -1 0 8350 0 -1 1830
box -12 -8 32 272
use FILL  FILL_1__1820_
timestamp 1701859473
transform -1 0 8430 0 1 1310
box -12 -8 32 272
use FILL  FILL_1__1821_
timestamp 1701859473
transform -1 0 4870 0 1 1310
box -12 -8 32 272
use FILL  FILL_1__1822_
timestamp 1701859473
transform -1 0 4670 0 -1 790
box -12 -8 32 272
use FILL  FILL_1__1823_
timestamp 1701859473
transform -1 0 4210 0 -1 790
box -12 -8 32 272
use FILL  FILL_1__1824_
timestamp 1701859473
transform 1 0 4590 0 1 2350
box -12 -8 32 272
use FILL  FILL_1__1825_
timestamp 1701859473
transform 1 0 5650 0 1 1830
box -12 -8 32 272
use FILL  FILL_1__1826_
timestamp 1701859473
transform 1 0 8150 0 -1 270
box -12 -8 32 272
use FILL  FILL_1__1827_
timestamp 1701859473
transform 1 0 9290 0 -1 790
box -12 -8 32 272
use FILL  FILL_1__1828_
timestamp 1701859473
transform 1 0 8450 0 1 270
box -12 -8 32 272
use FILL  FILL_1__1829_
timestamp 1701859473
transform 1 0 5750 0 1 270
box -12 -8 32 272
use FILL  FILL_1__1830_
timestamp 1701859473
transform 1 0 3190 0 1 4430
box -12 -8 32 272
use FILL  FILL_1__1831_
timestamp 1701859473
transform -1 0 7970 0 -1 790
box -12 -8 32 272
use FILL  FILL_1__1832_
timestamp 1701859473
transform 1 0 6470 0 -1 790
box -12 -8 32 272
use FILL  FILL_1__1833_
timestamp 1701859473
transform -1 0 670 0 1 270
box -12 -8 32 272
use FILL  FILL_1__1834_
timestamp 1701859473
transform 1 0 1110 0 -1 1310
box -12 -8 32 272
use FILL  FILL_1__1835_
timestamp 1701859473
transform -1 0 2490 0 -1 1310
box -12 -8 32 272
use FILL  FILL_1__1836_
timestamp 1701859473
transform 1 0 1050 0 1 790
box -12 -8 32 272
use FILL  FILL_1__1837_
timestamp 1701859473
transform -1 0 2450 0 1 790
box -12 -8 32 272
use FILL  FILL_1__1838_
timestamp 1701859473
transform 1 0 2190 0 1 790
box -12 -8 32 272
use FILL  FILL_1__1839_
timestamp 1701859473
transform -1 0 250 0 1 270
box -12 -8 32 272
use FILL  FILL_1__1840_
timestamp 1701859473
transform -1 0 890 0 1 2870
box -12 -8 32 272
use FILL  FILL_1__1841_
timestamp 1701859473
transform 1 0 3670 0 1 2870
box -12 -8 32 272
use FILL  FILL_1__1842_
timestamp 1701859473
transform -1 0 2930 0 -1 1830
box -12 -8 32 272
use FILL  FILL_1__1843_
timestamp 1701859473
transform -1 0 3890 0 -1 2350
box -12 -8 32 272
use FILL  FILL_1__1844_
timestamp 1701859473
transform 1 0 3790 0 -1 2870
box -12 -8 32 272
use FILL  FILL_1__1845_
timestamp 1701859473
transform -1 0 1730 0 -1 4950
box -12 -8 32 272
use FILL  FILL_1__1846_
timestamp 1701859473
transform 1 0 4090 0 1 4430
box -12 -8 32 272
use FILL  FILL_1__1847_
timestamp 1701859473
transform 1 0 3410 0 1 4430
box -12 -8 32 272
use FILL  FILL_1__1848_
timestamp 1701859473
transform 1 0 3850 0 1 4430
box -12 -8 32 272
use FILL  FILL_1__1849_
timestamp 1701859473
transform -1 0 4050 0 -1 2870
box -12 -8 32 272
use FILL  FILL_1__1850_
timestamp 1701859473
transform -1 0 870 0 1 790
box -12 -8 32 272
use FILL  FILL_1__1851_
timestamp 1701859473
transform 1 0 1530 0 -1 1830
box -12 -8 32 272
use FILL  FILL_1__1852_
timestamp 1701859473
transform -1 0 2350 0 1 2350
box -12 -8 32 272
use FILL  FILL_1__1853_
timestamp 1701859473
transform 1 0 30 0 -1 2350
box -12 -8 32 272
use FILL  FILL_1__1854_
timestamp 1701859473
transform 1 0 2270 0 -1 2350
box -12 -8 32 272
use FILL  FILL_1__1855_
timestamp 1701859473
transform -1 0 2530 0 -1 2350
box -12 -8 32 272
use FILL  FILL_1__1856_
timestamp 1701859473
transform 1 0 1430 0 -1 790
box -12 -8 32 272
use FILL  FILL_1__1857_
timestamp 1701859473
transform -1 0 2630 0 -1 790
box -12 -8 32 272
use FILL  FILL_1__1858_
timestamp 1701859473
transform 1 0 2370 0 -1 790
box -12 -8 32 272
use FILL  FILL_1__1859_
timestamp 1701859473
transform 1 0 2150 0 -1 790
box -12 -8 32 272
use FILL  FILL_1__1860_
timestamp 1701859473
transform -1 0 1690 0 -1 790
box -12 -8 32 272
use FILL  FILL_1__1861_
timestamp 1701859473
transform -1 0 1930 0 -1 790
box -12 -8 32 272
use FILL  FILL_1__1862_
timestamp 1701859473
transform -1 0 2010 0 1 270
box -12 -8 32 272
use FILL  FILL_1__1863_
timestamp 1701859473
transform 1 0 2230 0 1 270
box -12 -8 32 272
use FILL  FILL_1__1864_
timestamp 1701859473
transform 1 0 3470 0 1 270
box -12 -8 32 272
use FILL  FILL_1__1865_
timestamp 1701859473
transform 1 0 7270 0 -1 1310
box -12 -8 32 272
use FILL  FILL_1__1866_
timestamp 1701859473
transform 1 0 3630 0 -1 1310
box -12 -8 32 272
use FILL  FILL_1__1867_
timestamp 1701859473
transform 1 0 1090 0 -1 1830
box -12 -8 32 272
use FILL  FILL_1__1868_
timestamp 1701859473
transform 1 0 1530 0 1 1310
box -12 -8 32 272
use FILL  FILL_1__1869_
timestamp 1701859473
transform 1 0 1950 0 1 1310
box -12 -8 32 272
use FILL  FILL_1__1870_
timestamp 1701859473
transform -1 0 1570 0 -1 1310
box -12 -8 32 272
use FILL  FILL_1__1871_
timestamp 1701859473
transform -1 0 2690 0 -1 1310
box -12 -8 32 272
use FILL  FILL_1__1872_
timestamp 1701859473
transform -1 0 470 0 1 790
box -12 -8 32 272
use FILL  FILL_1__1873_
timestamp 1701859473
transform 1 0 650 0 1 790
box -12 -8 32 272
use FILL  FILL_1__1874_
timestamp 1701859473
transform -1 0 1290 0 1 790
box -12 -8 32 272
use FILL  FILL_1__1875_
timestamp 1701859473
transform 1 0 870 0 -1 790
box -12 -8 32 272
use FILL  FILL_1__1876_
timestamp 1701859473
transform 1 0 1190 0 -1 790
box -12 -8 32 272
use FILL  FILL_1__1877_
timestamp 1701859473
transform 1 0 2130 0 1 4950
box -12 -8 32 272
use FILL  FILL_1__1878_
timestamp 1701859473
transform 1 0 470 0 -1 1310
box -12 -8 32 272
use FILL  FILL_1__1879_
timestamp 1701859473
transform 1 0 690 0 1 1310
box -12 -8 32 272
use FILL  FILL_1__1880_
timestamp 1701859473
transform -1 0 1950 0 -1 4950
box -12 -8 32 272
use FILL  FILL_1__1881_
timestamp 1701859473
transform -1 0 2190 0 -1 4950
box -12 -8 32 272
use FILL  FILL_1__1882_
timestamp 1701859473
transform 1 0 1510 0 -1 3390
box -12 -8 32 272
use FILL  FILL_1__1883_
timestamp 1701859473
transform 1 0 990 0 -1 3390
box -12 -8 32 272
use FILL  FILL_1__1884_
timestamp 1701859473
transform -1 0 4010 0 1 3390
box -12 -8 32 272
use FILL  FILL_1__1885_
timestamp 1701859473
transform -1 0 3730 0 -1 3390
box -12 -8 32 272
use FILL  FILL_1__1886_
timestamp 1701859473
transform 1 0 3470 0 -1 3390
box -12 -8 32 272
use FILL  FILL_1__1887_
timestamp 1701859473
transform -1 0 3450 0 1 2870
box -12 -8 32 272
use FILL  FILL_1__1888_
timestamp 1701859473
transform -1 0 2490 0 1 270
box -12 -8 32 272
use FILL  FILL_1__1889_
timestamp 1701859473
transform 1 0 1630 0 -1 2870
box -12 -8 32 272
use FILL  FILL_1__1890_
timestamp 1701859473
transform -1 0 270 0 -1 1830
box -12 -8 32 272
use FILL  FILL_1__1891_
timestamp 1701859473
transform 1 0 30 0 -1 1830
box -12 -8 32 272
use FILL  FILL_1__1892_
timestamp 1701859473
transform 1 0 4870 0 -1 3390
box -12 -8 32 272
use FILL  FILL_1__1893_
timestamp 1701859473
transform 1 0 3870 0 1 1830
box -12 -8 32 272
use FILL  FILL_1__1894_
timestamp 1701859473
transform 1 0 4070 0 1 1830
box -12 -8 32 272
use FILL  FILL_1__1895_
timestamp 1701859473
transform -1 0 1810 0 1 1830
box -12 -8 32 272
use FILL  FILL_1__1896_
timestamp 1701859473
transform 1 0 1830 0 -1 2350
box -12 -8 32 272
use FILL  FILL_1__1897_
timestamp 1701859473
transform 1 0 3450 0 1 2350
box -12 -8 32 272
use FILL  FILL_1__1898_
timestamp 1701859473
transform 1 0 3230 0 1 2350
box -12 -8 32 272
use FILL  FILL_1__1899_
timestamp 1701859473
transform -1 0 3210 0 -1 2350
box -12 -8 32 272
use FILL  FILL_1__1900_
timestamp 1701859473
transform -1 0 4050 0 -1 1830
box -12 -8 32 272
use FILL  FILL_1__1901_
timestamp 1701859473
transform -1 0 690 0 1 1830
box -12 -8 32 272
use FILL  FILL_1__1902_
timestamp 1701859473
transform 1 0 4990 0 1 1830
box -12 -8 32 272
use FILL  FILL_1__1903_
timestamp 1701859473
transform 1 0 3310 0 1 1310
box -12 -8 32 272
use FILL  FILL_1__1904_
timestamp 1701859473
transform -1 0 3410 0 -1 1310
box -12 -8 32 272
use FILL  FILL_1__1905_
timestamp 1701859473
transform 1 0 2950 0 1 270
box -12 -8 32 272
use FILL  FILL_1__1906_
timestamp 1701859473
transform 1 0 230 0 1 2350
box -12 -8 32 272
use FILL  FILL_1__1907_
timestamp 1701859473
transform -1 0 2990 0 -1 2350
box -12 -8 32 272
use FILL  FILL_1__1908_
timestamp 1701859473
transform 1 0 6410 0 -1 2350
box -12 -8 32 272
use FILL  FILL_1__1909_
timestamp 1701859473
transform -1 0 6010 0 -1 2350
box -12 -8 32 272
use FILL  FILL_1__1910_
timestamp 1701859473
transform -1 0 5510 0 -1 2350
box -12 -8 32 272
use FILL  FILL_1__1911_
timestamp 1701859473
transform -1 0 670 0 1 2870
box -12 -8 32 272
use FILL  FILL_1__1912_
timestamp 1701859473
transform -1 0 3270 0 1 3910
box -12 -8 32 272
use FILL  FILL_1__1913_
timestamp 1701859473
transform -1 0 990 0 -1 2870
box -12 -8 32 272
use FILL  FILL_1__1914_
timestamp 1701859473
transform -1 0 1430 0 1 3390
box -12 -8 32 272
use FILL  FILL_1__1915_
timestamp 1701859473
transform 1 0 2510 0 1 3390
box -12 -8 32 272
use FILL  FILL_1__1916_
timestamp 1701859473
transform -1 0 3370 0 1 3390
box -12 -8 32 272
use FILL  FILL_1__1917_
timestamp 1701859473
transform -1 0 4650 0 -1 3390
box -12 -8 32 272
use FILL  FILL_1__1918_
timestamp 1701859473
transform 1 0 1690 0 1 4950
box -12 -8 32 272
use FILL  FILL_1__1919_
timestamp 1701859473
transform -1 0 1210 0 -1 2870
box -12 -8 32 272
use FILL  FILL_1__1920_
timestamp 1701859473
transform -1 0 4990 0 1 4430
box -12 -8 32 272
use FILL  FILL_1__1921_
timestamp 1701859473
transform 1 0 4750 0 1 4430
box -12 -8 32 272
use FILL  FILL_1__1922_
timestamp 1701859473
transform -1 0 4550 0 1 4430
box -12 -8 32 272
use FILL  FILL_1__1923_
timestamp 1701859473
transform 1 0 4410 0 -1 3390
box -12 -8 32 272
use FILL  FILL_1__1924_
timestamp 1701859473
transform 1 0 1910 0 1 4950
box -12 -8 32 272
use FILL  FILL_1__1925_
timestamp 1701859473
transform 1 0 6050 0 -1 4430
box -12 -8 32 272
use FILL  FILL_1__1926_
timestamp 1701859473
transform 1 0 670 0 -1 1310
box -12 -8 32 272
use FILL  FILL_1__1927_
timestamp 1701859473
transform 1 0 2910 0 -1 1310
box -12 -8 32 272
use FILL  FILL_1__1928_
timestamp 1701859473
transform -1 0 3170 0 -1 1310
box -12 -8 32 272
use FILL  FILL_1__1929_
timestamp 1701859473
transform 1 0 3350 0 1 790
box -12 -8 32 272
use FILL  FILL_1__1930_
timestamp 1701859473
transform 1 0 3170 0 1 270
box -12 -8 32 272
use FILL  FILL_1__1931_
timestamp 1701859473
transform 1 0 3770 0 1 270
box -12 -8 32 272
use FILL  FILL_1__1932_
timestamp 1701859473
transform -1 0 4010 0 1 270
box -12 -8 32 272
use FILL  FILL_1__1933_
timestamp 1701859473
transform -1 0 1810 0 1 270
box -12 -8 32 272
use FILL  FILL_1__1934_
timestamp 1701859473
transform -1 0 5430 0 1 790
box -12 -8 32 272
use FILL  FILL_1__1935_
timestamp 1701859473
transform 1 0 5550 0 -1 270
box -12 -8 32 272
use FILL  FILL_1__1936_
timestamp 1701859473
transform -1 0 8310 0 1 3390
box -12 -8 32 272
use FILL  FILL_1__1937_
timestamp 1701859473
transform -1 0 7530 0 -1 270
box -12 -8 32 272
use FILL  FILL_1__1938_
timestamp 1701859473
transform -1 0 7730 0 -1 270
box -12 -8 32 272
use FILL  FILL_1__1939_
timestamp 1701859473
transform -1 0 6650 0 -1 270
box -12 -8 32 272
use FILL  FILL_1__1940_
timestamp 1701859473
transform -1 0 5770 0 -1 270
box -12 -8 32 272
use FILL  FILL_1__1941_
timestamp 1701859473
transform 1 0 5790 0 -1 790
box -12 -8 32 272
use FILL  FILL_1__1942_
timestamp 1701859473
transform 1 0 4770 0 -1 1310
box -12 -8 32 272
use FILL  FILL_1__1943_
timestamp 1701859473
transform 1 0 8030 0 1 270
box -12 -8 32 272
use FILL  FILL_1__1944_
timestamp 1701859473
transform -1 0 8270 0 1 270
box -12 -8 32 272
use FILL  FILL_1__1945_
timestamp 1701859473
transform 1 0 7810 0 1 270
box -12 -8 32 272
use FILL  FILL_1__1946_
timestamp 1701859473
transform -1 0 6010 0 1 270
box -12 -8 32 272
use FILL  FILL_1__1947_
timestamp 1701859473
transform -1 0 6030 0 -1 790
box -12 -8 32 272
use FILL  FILL_1__1948_
timestamp 1701859473
transform 1 0 5310 0 -1 790
box -12 -8 32 272
use FILL  FILL_1__1949_
timestamp 1701859473
transform 1 0 4550 0 -1 1310
box -12 -8 32 272
use FILL  FILL_1__1950_
timestamp 1701859473
transform -1 0 8190 0 -1 790
box -12 -8 32 272
use FILL  FILL_1__1951_
timestamp 1701859473
transform 1 0 470 0 -1 2350
box -12 -8 32 272
use FILL  FILL_1__1952_
timestamp 1701859473
transform -1 0 5650 0 1 2350
box -12 -8 32 272
use FILL  FILL_1__1953_
timestamp 1701859473
transform 1 0 5750 0 -1 2350
box -12 -8 32 272
use FILL  FILL_1__1954_
timestamp 1701859473
transform 1 0 8130 0 -1 1310
box -12 -8 32 272
use FILL  FILL_1__1955_
timestamp 1701859473
transform -1 0 8670 0 1 1310
box -12 -8 32 272
use FILL  FILL_1__1956_
timestamp 1701859473
transform -1 0 6210 0 -1 1310
box -12 -8 32 272
use FILL  FILL_1__1957_
timestamp 1701859473
transform -1 0 5970 0 -1 1310
box -12 -8 32 272
use FILL  FILL_1__1958_
timestamp 1701859473
transform 1 0 5230 0 -1 1310
box -12 -8 32 272
use FILL  FILL_1__1959_
timestamp 1701859473
transform 1 0 5670 0 -1 2870
box -12 -8 32 272
use FILL  FILL_1__1960_
timestamp 1701859473
transform -1 0 6110 0 -1 2870
box -12 -8 32 272
use FILL  FILL_1__1961_
timestamp 1701859473
transform -1 0 4370 0 1 2350
box -12 -8 32 272
use FILL  FILL_1__1962_
timestamp 1701859473
transform 1 0 5830 0 1 2350
box -12 -8 32 272
use FILL  FILL_1__1963_
timestamp 1701859473
transform 1 0 5290 0 1 1310
box -12 -8 32 272
use FILL  FILL_1__1964_
timestamp 1701859473
transform 1 0 9110 0 1 1310
box -12 -8 32 272
use FILL  FILL_1__1965_
timestamp 1701859473
transform 1 0 7510 0 1 790
box -12 -8 32 272
use FILL  FILL_1__1966_
timestamp 1701859473
transform -1 0 7630 0 1 270
box -12 -8 32 272
use FILL  FILL_1__1967_
timestamp 1701859473
transform -1 0 6690 0 1 270
box -12 -8 32 272
use FILL  FILL_1__1968_
timestamp 1701859473
transform 1 0 5470 0 -1 1310
box -12 -8 32 272
use FILL  FILL_1__1969_
timestamp 1701859473
transform 1 0 5670 0 1 2870
box -12 -8 32 272
use FILL  FILL_1__1970_
timestamp 1701859473
transform 1 0 5310 0 -1 3390
box -12 -8 32 272
use FILL  FILL_1__1971_
timestamp 1701859473
transform 1 0 5750 0 1 3910
box -12 -8 32 272
use FILL  FILL_1__1972_
timestamp 1701859473
transform 1 0 5690 0 1 4950
box -12 -8 32 272
use FILL  FILL_1__1973_
timestamp 1701859473
transform -1 0 6030 0 -1 3910
box -12 -8 32 272
use FILL  FILL_1__1974_
timestamp 1701859473
transform 1 0 6210 0 -1 3910
box -12 -8 32 272
use FILL  FILL_1__1975_
timestamp 1701859473
transform -1 0 6010 0 1 3910
box -12 -8 32 272
use FILL  FILL_1__1976_
timestamp 1701859473
transform -1 0 6470 0 -1 3910
box -12 -8 32 272
use FILL  FILL_1__1977_
timestamp 1701859473
transform 1 0 6790 0 1 2870
box -12 -8 32 272
use FILL  FILL_1__1978_
timestamp 1701859473
transform -1 0 6330 0 -1 2870
box -12 -8 32 272
use FILL  FILL_1__1979_
timestamp 1701859473
transform 1 0 6370 0 1 2870
box -12 -8 32 272
use FILL  FILL_1__1980_
timestamp 1701859473
transform 1 0 6570 0 1 2870
box -12 -8 32 272
use FILL  FILL_1__1981_
timestamp 1701859473
transform 1 0 6150 0 1 2870
box -12 -8 32 272
use FILL  FILL_1__1982_
timestamp 1701859473
transform -1 0 5610 0 -1 1830
box -12 -8 32 272
use FILL  FILL_1__1983_
timestamp 1701859473
transform -1 0 4710 0 -1 270
box -12 -8 32 272
use FILL  FILL_1__1984_
timestamp 1701859473
transform -1 0 6410 0 -1 1310
box -12 -8 32 272
use FILL  FILL_1__1985_
timestamp 1701859473
transform 1 0 4970 0 -1 1310
box -12 -8 32 272
use FILL  FILL_1__1986_
timestamp 1701859473
transform 1 0 8170 0 1 790
box -12 -8 32 272
use FILL  FILL_1__1987_
timestamp 1701859473
transform 1 0 6850 0 1 1310
box -12 -8 32 272
use FILL  FILL_1__1988_
timestamp 1701859473
transform -1 0 7310 0 1 1310
box -12 -8 32 272
use FILL  FILL_1__1989_
timestamp 1701859473
transform 1 0 2670 0 -1 5470
box -12 -8 32 272
use FILL  FILL_1__1990_
timestamp 1701859473
transform 1 0 1990 0 1 1830
box -12 -8 32 272
use FILL  FILL_1__1991_
timestamp 1701859473
transform -1 0 2710 0 1 1830
box -12 -8 32 272
use FILL  FILL_1__1992_
timestamp 1701859473
transform -1 0 4110 0 -1 2350
box -12 -8 32 272
use FILL  FILL_1__1993_
timestamp 1701859473
transform -1 0 4350 0 -1 2350
box -12 -8 32 272
use FILL  FILL_1__1994_
timestamp 1701859473
transform 1 0 2450 0 1 1830
box -12 -8 32 272
use FILL  FILL_1__1995_
timestamp 1701859473
transform 1 0 2930 0 1 1830
box -12 -8 32 272
use FILL  FILL_1__1996_
timestamp 1701859473
transform -1 0 6610 0 1 790
box -12 -8 32 272
use FILL  FILL_1__1997_
timestamp 1701859473
transform -1 0 4950 0 1 790
box -12 -8 32 272
use FILL  FILL_1__1998_
timestamp 1701859473
transform 1 0 4210 0 1 270
box -12 -8 32 272
use FILL  FILL_1__1999_
timestamp 1701859473
transform -1 0 3810 0 -1 270
box -12 -8 32 272
use FILL  FILL_1__2000_
timestamp 1701859473
transform -1 0 4490 0 -1 270
box -12 -8 32 272
use FILL  FILL_1__2001_
timestamp 1701859473
transform -1 0 5870 0 -1 2870
box -12 -8 32 272
use FILL  FILL_1__2002_
timestamp 1701859473
transform -1 0 1810 0 1 2870
box -12 -8 32 272
use FILL  FILL_1__2003_
timestamp 1701859473
transform 1 0 1310 0 -1 3390
box -12 -8 32 272
use FILL  FILL_1__2004_
timestamp 1701859473
transform 1 0 2730 0 -1 3390
box -12 -8 32 272
use FILL  FILL_1__2005_
timestamp 1701859473
transform -1 0 3010 0 1 2870
box -12 -8 32 272
use FILL  FILL_1__2006_
timestamp 1701859473
transform 1 0 2750 0 1 2870
box -12 -8 32 272
use FILL  FILL_1__2007_
timestamp 1701859473
transform 1 0 6770 0 -1 2870
box -12 -8 32 272
use FILL  FILL_1__2008_
timestamp 1701859473
transform 1 0 450 0 -1 1830
box -12 -8 32 272
use FILL  FILL_1__2009_
timestamp 1701859473
transform -1 0 3970 0 -1 3390
box -12 -8 32 272
use FILL  FILL_1__2010_
timestamp 1701859473
transform -1 0 4270 0 -1 2870
box -12 -8 32 272
use FILL  FILL_1__2011_
timestamp 1701859473
transform -1 0 2010 0 1 790
box -12 -8 32 272
use FILL  FILL_1__2012_
timestamp 1701859473
transform 1 0 1510 0 1 790
box -12 -8 32 272
use FILL  FILL_1__2013_
timestamp 1701859473
transform -1 0 1770 0 1 790
box -12 -8 32 272
use FILL  FILL_1__2014_
timestamp 1701859473
transform 1 0 4430 0 1 1310
box -12 -8 32 272
use FILL  FILL_1__2015_
timestamp 1701859473
transform 1 0 3150 0 1 1830
box -12 -8 32 272
use FILL  FILL_1__2016_
timestamp 1701859473
transform -1 0 3650 0 1 1830
box -12 -8 32 272
use FILL  FILL_1__2017_
timestamp 1701859473
transform -1 0 5170 0 -1 1830
box -12 -8 32 272
use FILL  FILL_1__2018_
timestamp 1701859473
transform 1 0 4930 0 -1 1830
box -12 -8 32 272
use FILL  FILL_1__2019_
timestamp 1701859473
transform -1 0 5450 0 -1 2870
box -12 -8 32 272
use FILL  FILL_1__2020_
timestamp 1701859473
transform -1 0 5210 0 -1 2870
box -12 -8 32 272
use FILL  FILL_1__2021_
timestamp 1701859473
transform -1 0 6850 0 -1 1310
box -12 -8 32 272
use FILL  FILL_1__2022_
timestamp 1701859473
transform -1 0 7090 0 1 790
box -12 -8 32 272
use FILL  FILL_1__2023_
timestamp 1701859473
transform 1 0 8130 0 1 1830
box -12 -8 32 272
use FILL  FILL_1__2024_
timestamp 1701859473
transform -1 0 8350 0 1 1830
box -12 -8 32 272
use FILL  FILL_1__2025_
timestamp 1701859473
transform 1 0 9510 0 -1 790
box -12 -8 32 272
use FILL  FILL_1__2026_
timestamp 1701859473
transform -1 0 8650 0 1 790
box -12 -8 32 272
use FILL  FILL_1__2027_
timestamp 1701859473
transform -1 0 6850 0 1 790
box -12 -8 32 272
use FILL  FILL_1__2028_
timestamp 1701859473
transform 1 0 6950 0 -1 790
box -12 -8 32 272
use FILL  FILL_1__2029_
timestamp 1701859473
transform 1 0 7390 0 1 270
box -12 -8 32 272
use FILL  FILL_1__2030_
timestamp 1701859473
transform -1 0 7070 0 -1 1310
box -12 -8 32 272
use FILL  FILL_1__2031_
timestamp 1701859473
transform 1 0 7390 0 -1 790
box -12 -8 32 272
use FILL  FILL_1__2032_
timestamp 1701859473
transform -1 0 8690 0 1 270
box -12 -8 32 272
use FILL  FILL_1__2033_
timestamp 1701859473
transform 1 0 8170 0 1 1310
box -12 -8 32 272
use FILL  FILL_1__2034_
timestamp 1701859473
transform -1 0 8850 0 -1 1310
box -12 -8 32 272
use FILL  FILL_1__2035_
timestamp 1701859473
transform -1 0 8430 0 1 790
box -12 -8 32 272
use FILL  FILL_1__2036_
timestamp 1701859473
transform -1 0 8590 0 -1 1830
box -12 -8 32 272
use FILL  FILL_1__2037_
timestamp 1701859473
transform -1 0 8650 0 -1 790
box -12 -8 32 272
use FILL  FILL_1__2038_
timestamp 1701859473
transform 1 0 7950 0 1 790
box -12 -8 32 272
use FILL  FILL_1__2039_
timestamp 1701859473
transform 1 0 7730 0 1 790
box -12 -8 32 272
use FILL  FILL_1__2040_
timestamp 1701859473
transform -1 0 7650 0 -1 790
box -12 -8 32 272
use FILL  FILL_1__2041_
timestamp 1701859473
transform -1 0 6870 0 -1 270
box -12 -8 32 272
use FILL  FILL_1__2042_
timestamp 1701859473
transform 1 0 8850 0 -1 790
box -12 -8 32 272
use FILL  FILL_1__2043_
timestamp 1701859473
transform 1 0 7170 0 1 270
box -12 -8 32 272
use FILL  FILL_1__2044_
timestamp 1701859473
transform 1 0 6910 0 1 270
box -12 -8 32 272
use FILL  FILL_1__2045_
timestamp 1701859473
transform -1 0 6230 0 1 270
box -12 -8 32 272
use FILL  FILL_1__2046_
timestamp 1701859473
transform 1 0 6410 0 -1 270
box -12 -8 32 272
use FILL  FILL_1__2047_
timestamp 1701859473
transform -1 0 6190 0 -1 270
box -12 -8 32 272
use FILL  FILL_1__2048_
timestamp 1701859473
transform -1 0 5990 0 -1 270
box -12 -8 32 272
use FILL  FILL_1__2049_
timestamp 1701859473
transform -1 0 7170 0 -1 790
box -12 -8 32 272
use FILL  FILL_1__2050_
timestamp 1701859473
transform 1 0 1410 0 -1 2870
box -12 -8 32 272
use FILL  FILL_1__2051_
timestamp 1701859473
transform 1 0 6210 0 -1 2350
box -12 -8 32 272
use FILL  FILL_1__2052_
timestamp 1701859473
transform -1 0 6110 0 1 790
box -12 -8 32 272
use FILL  FILL_1__2053_
timestamp 1701859473
transform -1 0 4330 0 1 1830
box -12 -8 32 272
use FILL  FILL_1__2054_
timestamp 1701859473
transform 1 0 2830 0 1 1310
box -12 -8 32 272
use FILL  FILL_1__2055_
timestamp 1701859473
transform -1 0 3090 0 1 1310
box -12 -8 32 272
use FILL  FILL_1__2056_
timestamp 1701859473
transform -1 0 1810 0 -1 1310
box -12 -8 32 272
use FILL  FILL_1__2057_
timestamp 1701859473
transform 1 0 2670 0 1 790
box -12 -8 32 272
use FILL  FILL_1__2058_
timestamp 1701859473
transform 1 0 3590 0 1 790
box -12 -8 32 272
use FILL  FILL_1__2059_
timestamp 1701859473
transform 1 0 3830 0 1 790
box -12 -8 32 272
use FILL  FILL_1__2060_
timestamp 1701859473
transform -1 0 4070 0 1 790
box -12 -8 32 272
use FILL  FILL_1__2061_
timestamp 1701859473
transform -1 0 2930 0 -1 270
box -12 -8 32 272
use FILL  FILL_1__2062_
timestamp 1701859473
transform 1 0 2710 0 1 270
box -12 -8 32 272
use FILL  FILL_1__2063_
timestamp 1701859473
transform 1 0 3090 0 -1 270
box -12 -8 32 272
use FILL  FILL_1__2064_
timestamp 1701859473
transform 1 0 3330 0 -1 270
box -12 -8 32 272
use FILL  FILL_1__2065_
timestamp 1701859473
transform -1 0 3570 0 -1 270
box -12 -8 32 272
use FILL  FILL_1__2066_
timestamp 1701859473
transform -1 0 5350 0 -1 270
box -12 -8 32 272
use FILL  FILL_1__2067_
timestamp 1701859473
transform 1 0 7290 0 1 790
box -12 -8 32 272
use FILL  FILL_1__2068_
timestamp 1701859473
transform 1 0 5850 0 1 790
box -12 -8 32 272
use FILL  FILL_1__2069_
timestamp 1701859473
transform 1 0 3330 0 -1 1830
box -12 -8 32 272
use FILL  FILL_1__2070_
timestamp 1701859473
transform -1 0 3810 0 -1 1830
box -12 -8 32 272
use FILL  FILL_1__2071_
timestamp 1701859473
transform -1 0 5650 0 1 790
box -12 -8 32 272
use FILL  FILL_1__2072_
timestamp 1701859473
transform -1 0 7710 0 1 1310
box -12 -8 32 272
use FILL  FILL_1__2073_
timestamp 1701859473
transform 1 0 6590 0 1 1310
box -12 -8 32 272
use FILL  FILL_1__2074_
timestamp 1701859473
transform 1 0 1730 0 1 1310
box -12 -8 32 272
use FILL  FILL_1__2075_
timestamp 1701859473
transform -1 0 2210 0 1 1310
box -12 -8 32 272
use FILL  FILL_1__2076_
timestamp 1701859473
transform -1 0 2250 0 -1 1310
box -12 -8 32 272
use FILL  FILL_1__2077_
timestamp 1701859473
transform 1 0 4110 0 -1 1310
box -12 -8 32 272
use FILL  FILL_1__2078_
timestamp 1701859473
transform -1 0 2250 0 1 1830
box -12 -8 32 272
use FILL  FILL_1__2079_
timestamp 1701859473
transform -1 0 890 0 -1 1830
box -12 -8 32 272
use FILL  FILL_1__2080_
timestamp 1701859473
transform 1 0 2210 0 -1 1830
box -12 -8 32 272
use FILL  FILL_1__2081_
timestamp 1701859473
transform 1 0 2450 0 -1 1830
box -12 -8 32 272
use FILL  FILL_1__2082_
timestamp 1701859473
transform -1 0 2670 0 -1 1830
box -12 -8 32 272
use FILL  FILL_1__2083_
timestamp 1701859473
transform 1 0 4350 0 -1 1310
box -12 -8 32 272
use FILL  FILL_1__2084_
timestamp 1701859473
transform -1 0 5190 0 1 790
box -12 -8 32 272
use FILL  FILL_1__2085_
timestamp 1701859473
transform -1 0 5030 0 -1 270
box -12 -8 32 272
use FILL  FILL_1__2086_
timestamp 1701859473
transform -1 0 4250 0 -1 270
box -12 -8 32 272
use FILL  FILL_1__2087_
timestamp 1701859473
transform -1 0 4730 0 1 790
box -12 -8 32 272
use FILL  FILL_1__2088_
timestamp 1701859473
transform -1 0 5570 0 1 270
box -12 -8 32 272
use FILL  FILL_1__2089_
timestamp 1701859473
transform 1 0 5330 0 1 270
box -12 -8 32 272
use FILL  FILL_1__2090_
timestamp 1701859473
transform -1 0 4910 0 -1 790
box -12 -8 32 272
use FILL  FILL_1__2091_
timestamp 1701859473
transform 1 0 3130 0 1 790
box -12 -8 32 272
use FILL  FILL_1__2092_
timestamp 1701859473
transform 1 0 2690 0 -1 270
box -12 -8 32 272
use FILL  FILL_1__2093_
timestamp 1701859473
transform -1 0 2850 0 -1 790
box -12 -8 32 272
use FILL  FILL_1__2094_
timestamp 1701859473
transform 1 0 2250 0 -1 270
box -12 -8 32 272
use FILL  FILL_1__2095_
timestamp 1701859473
transform 1 0 2450 0 -1 270
box -12 -8 32 272
use FILL  FILL_1__2096_
timestamp 1701859473
transform -1 0 4910 0 1 270
box -12 -8 32 272
use FILL  FILL_1__2097_
timestamp 1701859473
transform -1 0 5130 0 1 270
box -12 -8 32 272
use FILL  FILL_1__2098_
timestamp 1701859473
transform 1 0 4670 0 1 270
box -12 -8 32 272
use FILL  FILL_1__2099_
timestamp 1701859473
transform 1 0 3990 0 -1 270
box -12 -8 32 272
use FILL  FILL_1__2100_
timestamp 1701859473
transform -1 0 5850 0 -1 1830
box -12 -8 32 272
use FILL  FILL_1__2101_
timestamp 1701859473
transform -1 0 5770 0 1 1310
box -12 -8 32 272
use FILL  FILL_1__2102_
timestamp 1701859473
transform -1 0 6170 0 1 1310
box -12 -8 32 272
use FILL  FILL_1__2103_
timestamp 1701859473
transform 1 0 5730 0 -1 1310
box -12 -8 32 272
use FILL  FILL_1__2104_
timestamp 1701859473
transform -1 0 5970 0 1 1310
box -12 -8 32 272
use FILL  FILL_1__2105_
timestamp 1701859473
transform -1 0 4270 0 -1 1830
box -12 -8 32 272
use FILL  FILL_1__2106_
timestamp 1701859473
transform 1 0 3950 0 -1 790
box -12 -8 32 272
use FILL  FILL_1__2107_
timestamp 1701859473
transform -1 0 3530 0 -1 790
box -12 -8 32 272
use FILL  FILL_1__2108_
timestamp 1701859473
transform 1 0 2890 0 1 790
box -12 -8 32 272
use FILL  FILL_1__2109_
timestamp 1701859473
transform -1 0 3310 0 -1 790
box -12 -8 32 272
use FILL  FILL_1__2110_
timestamp 1701859473
transform 1 0 3070 0 -1 790
box -12 -8 32 272
use FILL  FILL_1__2111_
timestamp 1701859473
transform -1 0 3750 0 -1 790
box -12 -8 32 272
use FILL  FILL_1__2112_
timestamp 1701859473
transform -1 0 5110 0 -1 790
box -12 -8 32 272
use FILL  FILL_1__2113_
timestamp 1701859473
transform -1 0 5090 0 1 1310
box -12 -8 32 272
use FILL  FILL_1__2114_
timestamp 1701859473
transform -1 0 5530 0 1 1310
box -12 -8 32 272
use FILL  FILL_1__2115_
timestamp 1701859473
transform -1 0 5570 0 -1 790
box -12 -8 32 272
use FILL  FILL_1__2116_
timestamp 1701859473
transform 1 0 2390 0 1 1310
box -12 -8 32 272
use FILL  FILL_1__2117_
timestamp 1701859473
transform 1 0 2590 0 1 1310
box -12 -8 32 272
use FILL  FILL_1__2118_
timestamp 1701859473
transform 1 0 3770 0 1 1310
box -12 -8 32 272
use FILL  FILL_1__2119_
timestamp 1701859473
transform -1 0 4030 0 1 1310
box -12 -8 32 272
use FILL  FILL_1__2120_
timestamp 1701859473
transform 1 0 3890 0 -1 1310
box -12 -8 32 272
use FILL  FILL_1__2121_
timestamp 1701859473
transform -1 0 4470 0 1 270
box -12 -8 32 272
use FILL  FILL_1__2122_
timestamp 1701859473
transform -1 0 2810 0 1 2350
box -12 -8 32 272
use FILL  FILL_1__2123_
timestamp 1701859473
transform 1 0 2750 0 -1 2350
box -12 -8 32 272
use FILL  FILL_1__2124_
timestamp 1701859473
transform -1 0 3650 0 -1 2350
box -12 -8 32 272
use FILL  FILL_1__2125_
timestamp 1701859473
transform 1 0 5770 0 -1 3390
box -12 -8 32 272
use FILL  FILL_1__2126_
timestamp 1701859473
transform 1 0 5450 0 1 2870
box -12 -8 32 272
use FILL  FILL_1__2127_
timestamp 1701859473
transform -1 0 5930 0 1 2870
box -12 -8 32 272
use FILL  FILL_1__2128_
timestamp 1701859473
transform 1 0 4550 0 1 2870
box -12 -8 32 272
use FILL  FILL_1__2129_
timestamp 1701859473
transform 1 0 5230 0 1 2870
box -12 -8 32 272
use FILL  FILL_1__2130_
timestamp 1701859473
transform -1 0 4590 0 -1 2350
box -12 -8 32 272
use FILL  FILL_1__2131_
timestamp 1701859473
transform 1 0 4630 0 1 1310
box -12 -8 32 272
use FILL  FILL_1__2132_
timestamp 1701859473
transform -1 0 4510 0 1 790
box -12 -8 32 272
use FILL  FILL_1__2133_
timestamp 1701859473
transform 1 0 4430 0 -1 790
box -12 -8 32 272
use FILL  FILL_1__2134_
timestamp 1701859473
transform 1 0 3550 0 -1 2870
box -12 -8 32 272
use FILL  FILL_1__2135_
timestamp 1701859473
transform 1 0 4170 0 -1 3390
box -12 -8 32 272
use FILL  FILL_1__2136_
timestamp 1701859473
transform -1 0 2710 0 1 3390
box -12 -8 32 272
use FILL  FILL_1__2137_
timestamp 1701859473
transform 1 0 2270 0 1 3390
box -12 -8 32 272
use FILL  FILL_1__2138_
timestamp 1701859473
transform 1 0 3070 0 -1 4430
box -12 -8 32 272
use FILL  FILL_1__2139_
timestamp 1701859473
transform -1 0 2850 0 -1 4430
box -12 -8 32 272
use FILL  FILL_1__2140_
timestamp 1701859473
transform 1 0 2770 0 1 4430
box -12 -8 32 272
use FILL  FILL_1__2141_
timestamp 1701859473
transform -1 0 3010 0 1 4430
box -12 -8 32 272
use FILL  FILL_1__2142_
timestamp 1701859473
transform 1 0 2890 0 1 3390
box -12 -8 32 272
use FILL  FILL_1__2143_
timestamp 1701859473
transform -1 0 7390 0 -1 3390
box -12 -8 32 272
use FILL  FILL_1__2144_
timestamp 1701859473
transform 1 0 2030 0 1 2870
box -12 -8 32 272
use FILL  FILL_1__2145_
timestamp 1701859473
transform -1 0 10010 0 -1 2870
box -12 -8 32 272
use FILL  FILL_1__2146_
timestamp 1701859473
transform -1 0 7590 0 -1 3390
box -12 -8 32 272
use FILL  FILL_1__2147_
timestamp 1701859473
transform 1 0 7550 0 -1 3910
box -12 -8 32 272
use FILL  FILL_1__2148_
timestamp 1701859473
transform 1 0 7390 0 1 3390
box -12 -8 32 272
use FILL  FILL_1__2149_
timestamp 1701859473
transform 1 0 7590 0 1 3390
box -12 -8 32 272
use FILL  FILL_1__2150_
timestamp 1701859473
transform -1 0 7850 0 1 3390
box -12 -8 32 272
use FILL  FILL_1__2151_
timestamp 1701859473
transform 1 0 7130 0 -1 3390
box -12 -8 32 272
use FILL  FILL_1__2152_
timestamp 1701859473
transform 1 0 6890 0 -1 3390
box -12 -8 32 272
use FILL  FILL_1__2153_
timestamp 1701859473
transform -1 0 6030 0 -1 3390
box -12 -8 32 272
use FILL  FILL_1__2154_
timestamp 1701859473
transform 1 0 2790 0 -1 7030
box -12 -8 32 272
use FILL  FILL_1__2155_
timestamp 1701859473
transform 1 0 6350 0 1 5990
box -12 -8 32 272
use FILL  FILL_1__2156_
timestamp 1701859473
transform -1 0 4570 0 1 3910
box -12 -8 32 272
use FILL  FILL_1__2157_
timestamp 1701859473
transform -1 0 4710 0 -1 4430
box -12 -8 32 272
use FILL  FILL_1__2158_
timestamp 1701859473
transform -1 0 2570 0 1 2350
box -12 -8 32 272
use FILL  FILL_1__2159_
timestamp 1701859473
transform 1 0 3470 0 1 3910
box -12 -8 32 272
use FILL  FILL_1__2160_
timestamp 1701859473
transform -1 0 3790 0 -1 4430
box -12 -8 32 272
use FILL  FILL_1__2161_
timestamp 1701859473
transform -1 0 3930 0 1 3910
box -12 -8 32 272
use FILL  FILL_1__2162_
timestamp 1701859473
transform -1 0 4370 0 1 3910
box -12 -8 32 272
use FILL  FILL_1__2163_
timestamp 1701859473
transform 1 0 3690 0 -1 3910
box -12 -8 32 272
use FILL  FILL_1__2164_
timestamp 1701859473
transform -1 0 510 0 -1 4950
box -12 -8 32 272
use FILL  FILL_1__2165_
timestamp 1701859473
transform -1 0 3210 0 -1 3910
box -12 -8 32 272
use FILL  FILL_1__2166_
timestamp 1701859473
transform 1 0 3910 0 -1 3910
box -12 -8 32 272
use FILL  FILL_1__2167_
timestamp 1701859473
transform 1 0 4110 0 1 3910
box -12 -8 32 272
use FILL  FILL_1__2168_
timestamp 1701859473
transform 1 0 3030 0 1 3910
box -12 -8 32 272
use FILL  FILL_1__2169_
timestamp 1701859473
transform 1 0 2390 0 -1 4430
box -12 -8 32 272
use FILL  FILL_1__2170_
timestamp 1701859473
transform -1 0 2650 0 -1 4430
box -12 -8 32 272
use FILL  FILL_1__2171_
timestamp 1701859473
transform 1 0 3990 0 -1 4430
box -12 -8 32 272
use FILL  FILL_1__2172_
timestamp 1701859473
transform 1 0 4230 0 -1 4430
box -12 -8 32 272
use FILL  FILL_1__2173_
timestamp 1701859473
transform -1 0 4470 0 -1 4430
box -12 -8 32 272
use FILL  FILL_1__2174_
timestamp 1701859473
transform 1 0 5970 0 1 7030
box -12 -8 32 272
use FILL  FILL_1__2175_
timestamp 1701859473
transform -1 0 2470 0 1 8070
box -12 -8 32 272
use FILL  FILL_1__2176_
timestamp 1701859473
transform -1 0 6390 0 -1 8070
box -12 -8 32 272
use FILL  FILL_1__2177_
timestamp 1701859473
transform 1 0 4910 0 1 8070
box -12 -8 32 272
use FILL  FILL_1__2178_
timestamp 1701859473
transform -1 0 4090 0 -1 8590
box -12 -8 32 272
use FILL  FILL_1__2179_
timestamp 1701859473
transform -1 0 5910 0 -1 8070
box -12 -8 32 272
use FILL  FILL_1__2180_
timestamp 1701859473
transform -1 0 2930 0 -1 9630
box -12 -8 32 272
use FILL  FILL_1__2181_
timestamp 1701859473
transform 1 0 4990 0 1 7550
box -12 -8 32 272
use FILL  FILL_1__2182_
timestamp 1701859473
transform 1 0 5510 0 -1 10150
box -12 -8 32 272
use FILL  FILL_1__2183_
timestamp 1701859473
transform -1 0 3490 0 1 10150
box -12 -8 32 272
use FILL  FILL_1__2184_
timestamp 1701859473
transform 1 0 4310 0 1 8070
box -12 -8 32 272
use FILL  FILL_1__2185_
timestamp 1701859473
transform 1 0 5910 0 1 10150
box -12 -8 32 272
use FILL  FILL_1__2186_
timestamp 1701859473
transform 1 0 3470 0 1 10670
box -12 -8 32 272
use FILL  FILL_1__2187_
timestamp 1701859473
transform -1 0 5390 0 -1 10670
box -12 -8 32 272
use FILL  FILL_1__2188_
timestamp 1701859473
transform 1 0 2070 0 -1 10670
box -12 -8 32 272
use FILL  FILL_1__2189_
timestamp 1701859473
transform 1 0 5630 0 -1 10670
box -12 -8 32 272
use FILL  FILL_1__2190_
timestamp 1701859473
transform -1 0 2790 0 1 10150
box -12 -8 32 272
use FILL  FILL_1__2191_
timestamp 1701859473
transform -1 0 5270 0 -1 10150
box -12 -8 32 272
use FILL  FILL_1__2192_
timestamp 1701859473
transform -1 0 11070 0 1 3910
box -12 -8 32 272
use FILL  FILL_1__2193_
timestamp 1701859473
transform 1 0 1190 0 -1 3910
box -12 -8 32 272
use FILL  FILL_1__2194_
timestamp 1701859473
transform 1 0 990 0 -1 3910
box -12 -8 32 272
use FILL  FILL_1__2195_
timestamp 1701859473
transform 1 0 2570 0 1 3910
box -12 -8 32 272
use FILL  FILL_1__2196_
timestamp 1701859473
transform 1 0 2810 0 1 3910
box -12 -8 32 272
use FILL  FILL_1__2197_
timestamp 1701859473
transform 1 0 5290 0 1 3910
box -12 -8 32 272
use FILL  FILL_1__2198_
timestamp 1701859473
transform 1 0 230 0 1 1830
box -12 -8 32 272
use FILL  FILL_1__2199_
timestamp 1701859473
transform -1 0 2790 0 -1 3910
box -12 -8 32 272
use FILL  FILL_1__2200_
timestamp 1701859473
transform 1 0 5310 0 -1 3910
box -12 -8 32 272
use FILL  FILL_1__2201_
timestamp 1701859473
transform -1 0 5550 0 1 3910
box -12 -8 32 272
use FILL  FILL_1__2202_
timestamp 1701859473
transform -1 0 8130 0 -1 4430
box -12 -8 32 272
use FILL  FILL_1__2203_
timestamp 1701859473
transform -1 0 4850 0 -1 3910
box -12 -8 32 272
use FILL  FILL_1__2204_
timestamp 1701859473
transform 1 0 5070 0 -1 3910
box -12 -8 32 272
use FILL  FILL_1__2205_
timestamp 1701859473
transform -1 0 8930 0 -1 3910
box -12 -8 32 272
use FILL  FILL_1__2206_
timestamp 1701859473
transform 1 0 9010 0 1 3910
box -12 -8 32 272
use FILL  FILL_1__2207_
timestamp 1701859473
transform 1 0 9470 0 -1 3910
box -12 -8 32 272
use FILL  FILL_1__2208_
timestamp 1701859473
transform -1 0 9730 0 -1 3910
box -12 -8 32 272
use FILL  FILL_1__2209_
timestamp 1701859473
transform -1 0 9530 0 1 4430
box -12 -8 32 272
use FILL  FILL_1__2210_
timestamp 1701859473
transform -1 0 10530 0 -1 4950
box -12 -8 32 272
use FILL  FILL_1__2211_
timestamp 1701859473
transform 1 0 9230 0 -1 3910
box -12 -8 32 272
use FILL  FILL_1__2212_
timestamp 1701859473
transform -1 0 8810 0 1 3910
box -12 -8 32 272
use FILL  FILL_1__2213_
timestamp 1701859473
transform -1 0 9250 0 1 3910
box -12 -8 32 272
use FILL  FILL_1__2214_
timestamp 1701859473
transform -1 0 9450 0 -1 4430
box -12 -8 32 272
use FILL  FILL_1__2215_
timestamp 1701859473
transform 1 0 9650 0 -1 4430
box -12 -8 32 272
use FILL  FILL_1__2216_
timestamp 1701859473
transform -1 0 9410 0 -1 7030
box -12 -8 32 272
use FILL  FILL_1__2217_
timestamp 1701859473
transform 1 0 9190 0 -1 4430
box -12 -8 32 272
use FILL  FILL_1__2218_
timestamp 1701859473
transform -1 0 9710 0 1 3910
box -12 -8 32 272
use FILL  FILL_1__2219_
timestamp 1701859473
transform 1 0 9890 0 1 3910
box -12 -8 32 272
use FILL  FILL_1__2220_
timestamp 1701859473
transform 1 0 10270 0 -1 4950
box -12 -8 32 272
use FILL  FILL_1__2221_
timestamp 1701859473
transform -1 0 9650 0 -1 7030
box -12 -8 32 272
use FILL  FILL_1__2222_
timestamp 1701859473
transform 1 0 10010 0 1 4430
box -12 -8 32 272
use FILL  FILL_1__2223_
timestamp 1701859473
transform -1 0 9910 0 -1 4430
box -12 -8 32 272
use FILL  FILL_1__2224_
timestamp 1701859473
transform -1 0 9770 0 1 4430
box -12 -8 32 272
use FILL  FILL_1__2225_
timestamp 1701859473
transform 1 0 10010 0 -1 4950
box -12 -8 32 272
use FILL  FILL_1__2226_
timestamp 1701859473
transform 1 0 8890 0 -1 7030
box -12 -8 32 272
use FILL  FILL_1__2227_
timestamp 1701859473
transform -1 0 9170 0 -1 7030
box -12 -8 32 272
use FILL  FILL_1__2228_
timestamp 1701859473
transform -1 0 5710 0 -1 7030
box -12 -8 32 272
use FILL  FILL_1__2229_
timestamp 1701859473
transform 1 0 4270 0 1 3390
box -12 -8 32 272
use FILL  FILL_1__2230_
timestamp 1701859473
transform -1 0 4370 0 -1 3910
box -12 -8 32 272
use FILL  FILL_1__2231_
timestamp 1701859473
transform -1 0 4150 0 -1 3910
box -12 -8 32 272
use FILL  FILL_1__2232_
timestamp 1701859473
transform 1 0 1550 0 1 2870
box -12 -8 32 272
use FILL  FILL_1__2233_
timestamp 1701859473
transform 1 0 2270 0 1 2870
box -12 -8 32 272
use FILL  FILL_1__2234_
timestamp 1701859473
transform -1 0 2530 0 1 2870
box -12 -8 32 272
use FILL  FILL_1__2235_
timestamp 1701859473
transform 1 0 6290 0 1 3390
box -12 -8 32 272
use FILL  FILL_1__2236_
timestamp 1701859473
transform -1 0 5570 0 -1 3910
box -12 -8 32 272
use FILL  FILL_1__2237_
timestamp 1701859473
transform -1 0 4610 0 -1 3910
box -12 -8 32 272
use FILL  FILL_1__2238_
timestamp 1701859473
transform 1 0 4670 0 -1 4950
box -12 -8 32 272
use FILL  FILL_1__2239_
timestamp 1701859473
transform 1 0 2790 0 1 4950
box -12 -8 32 272
use FILL  FILL_1__2240_
timestamp 1701859473
transform 1 0 2350 0 1 3910
box -12 -8 32 272
use FILL  FILL_1__2241_
timestamp 1701859473
transform -1 0 2370 0 1 4950
box -12 -8 32 272
use FILL  FILL_1__2242_
timestamp 1701859473
transform 1 0 2410 0 -1 4950
box -12 -8 32 272
use FILL  FILL_1__2243_
timestamp 1701859473
transform 1 0 2590 0 1 4950
box -12 -8 32 272
use FILL  FILL_1__2244_
timestamp 1701859473
transform 1 0 3010 0 1 4950
box -12 -8 32 272
use FILL  FILL_1__2245_
timestamp 1701859473
transform 1 0 2850 0 1 5990
box -12 -8 32 272
use FILL  FILL_1__2246_
timestamp 1701859473
transform 1 0 2870 0 -1 4950
box -12 -8 32 272
use FILL  FILL_1__2247_
timestamp 1701859473
transform -1 0 2990 0 -1 6510
box -12 -8 32 272
use FILL  FILL_1__2248_
timestamp 1701859473
transform 1 0 3450 0 -1 7030
box -12 -8 32 272
use FILL  FILL_1__2249_
timestamp 1701859473
transform 1 0 6230 0 1 7030
box -12 -8 32 272
use FILL  FILL_1__2250_
timestamp 1701859473
transform -1 0 10530 0 -1 7550
box -12 -8 32 272
use FILL  FILL_1__2251_
timestamp 1701859473
transform -1 0 10590 0 1 8070
box -12 -8 32 272
use FILL  FILL_1__2252_
timestamp 1701859473
transform -1 0 10890 0 -1 8070
box -12 -8 32 272
use FILL  FILL_1__2253_
timestamp 1701859473
transform -1 0 10650 0 -1 8070
box -12 -8 32 272
use FILL  FILL_1__2254_
timestamp 1701859473
transform 1 0 5350 0 1 8070
box -12 -8 32 272
use FILL  FILL_1__2255_
timestamp 1701859473
transform 1 0 2970 0 1 7030
box -12 -8 32 272
use FILL  FILL_1__2256_
timestamp 1701859473
transform -1 0 5090 0 1 7030
box -12 -8 32 272
use FILL  FILL_1__2257_
timestamp 1701859473
transform 1 0 5030 0 -1 7550
box -12 -8 32 272
use FILL  FILL_1__2258_
timestamp 1701859473
transform 1 0 5670 0 -1 8590
box -12 -8 32 272
use FILL  FILL_1__2259_
timestamp 1701859473
transform 1 0 10290 0 -1 7550
box -12 -8 32 272
use FILL  FILL_1__2260_
timestamp 1701859473
transform 1 0 9870 0 1 8070
box -12 -8 32 272
use FILL  FILL_1__2261_
timestamp 1701859473
transform -1 0 10170 0 1 7550
box -12 -8 32 272
use FILL  FILL_1__2262_
timestamp 1701859473
transform -1 0 9930 0 1 7550
box -12 -8 32 272
use FILL  FILL_1__2263_
timestamp 1701859473
transform 1 0 5430 0 1 7550
box -12 -8 32 272
use FILL  FILL_1__2264_
timestamp 1701859473
transform 1 0 1590 0 -1 6510
box -12 -8 32 272
use FILL  FILL_1__2265_
timestamp 1701859473
transform 1 0 1770 0 -1 6510
box -12 -8 32 272
use FILL  FILL_1__2266_
timestamp 1701859473
transform 1 0 3870 0 1 6510
box -12 -8 32 272
use FILL  FILL_1__2267_
timestamp 1701859473
transform -1 0 3630 0 -1 7550
box -12 -8 32 272
use FILL  FILL_1__2268_
timestamp 1701859473
transform 1 0 4310 0 -1 7550
box -12 -8 32 272
use FILL  FILL_1__2269_
timestamp 1701859473
transform 1 0 5630 0 1 7550
box -12 -8 32 272
use FILL  FILL_1__2270_
timestamp 1701859473
transform 1 0 8550 0 1 7550
box -12 -8 32 272
use FILL  FILL_1__2271_
timestamp 1701859473
transform -1 0 8830 0 -1 8070
box -12 -8 32 272
use FILL  FILL_1__2272_
timestamp 1701859473
transform -1 0 9090 0 -1 8070
box -12 -8 32 272
use FILL  FILL_1__2273_
timestamp 1701859473
transform -1 0 8590 0 -1 8070
box -12 -8 32 272
use FILL  FILL_1__2274_
timestamp 1701859473
transform -1 0 5950 0 -1 9630
box -12 -8 32 272
use FILL  FILL_1__2275_
timestamp 1701859473
transform -1 0 2250 0 1 8070
box -12 -8 32 272
use FILL  FILL_1__2276_
timestamp 1701859473
transform -1 0 3130 0 1 8070
box -12 -8 32 272
use FILL  FILL_1__2277_
timestamp 1701859473
transform -1 0 3610 0 -1 8590
box -12 -8 32 272
use FILL  FILL_1__2278_
timestamp 1701859473
transform 1 0 6510 0 1 9110
box -12 -8 32 272
use FILL  FILL_1__2279_
timestamp 1701859473
transform -1 0 10210 0 1 5990
box -12 -8 32 272
use FILL  FILL_1__2280_
timestamp 1701859473
transform 1 0 10390 0 1 5990
box -12 -8 32 272
use FILL  FILL_1__2281_
timestamp 1701859473
transform -1 0 10670 0 -1 5990
box -12 -8 32 272
use FILL  FILL_1__2282_
timestamp 1701859473
transform -1 0 10450 0 -1 6510
box -12 -8 32 272
use FILL  FILL_1__2283_
timestamp 1701859473
transform 1 0 5910 0 -1 8590
box -12 -8 32 272
use FILL  FILL_1__2284_
timestamp 1701859473
transform -1 0 2030 0 1 8070
box -12 -8 32 272
use FILL  FILL_1__2285_
timestamp 1701859473
transform -1 0 4090 0 1 8070
box -12 -8 32 272
use FILL  FILL_1__2286_
timestamp 1701859473
transform 1 0 4990 0 -1 8590
box -12 -8 32 272
use FILL  FILL_1__2287_
timestamp 1701859473
transform -1 0 6070 0 1 8590
box -12 -8 32 272
use FILL  FILL_1__2288_
timestamp 1701859473
transform -1 0 8790 0 1 7550
box -12 -8 32 272
use FILL  FILL_1__2289_
timestamp 1701859473
transform 1 0 8450 0 1 8070
box -12 -8 32 272
use FILL  FILL_1__2290_
timestamp 1701859473
transform -1 0 9950 0 -1 8070
box -12 -8 32 272
use FILL  FILL_1__2291_
timestamp 1701859473
transform -1 0 8730 0 1 8070
box -12 -8 32 272
use FILL  FILL_1__2292_
timestamp 1701859473
transform -1 0 6170 0 -1 9110
box -12 -8 32 272
use FILL  FILL_1__2293_
timestamp 1701859473
transform -1 0 2490 0 -1 8590
box -12 -8 32 272
use FILL  FILL_1__2294_
timestamp 1701859473
transform -1 0 3970 0 1 8590
box -12 -8 32 272
use FILL  FILL_1__2295_
timestamp 1701859473
transform 1 0 4890 0 1 8590
box -12 -8 32 272
use FILL  FILL_1__2296_
timestamp 1701859473
transform 1 0 6610 0 -1 9110
box -12 -8 32 272
use FILL  FILL_1__2297_
timestamp 1701859473
transform -1 0 9510 0 -1 5990
box -12 -8 32 272
use FILL  FILL_1__2298_
timestamp 1701859473
transform -1 0 9950 0 -1 5470
box -12 -8 32 272
use FILL  FILL_1__2299_
timestamp 1701859473
transform -1 0 9290 0 -1 6510
box -12 -8 32 272
use FILL  FILL_1__2300_
timestamp 1701859473
transform 1 0 9490 0 1 5990
box -12 -8 32 272
use FILL  FILL_1__2301_
timestamp 1701859473
transform 1 0 5530 0 1 9630
box -12 -8 32 272
use FILL  FILL_1__2302_
timestamp 1701859473
transform -1 0 3430 0 -1 9110
box -12 -8 32 272
use FILL  FILL_1__2303_
timestamp 1701859473
transform 1 0 2550 0 1 9110
box -12 -8 32 272
use FILL  FILL_1__2304_
timestamp 1701859473
transform 1 0 2750 0 -1 9110
box -12 -8 32 272
use FILL  FILL_1__2305_
timestamp 1701859473
transform -1 0 3730 0 1 8590
box -12 -8 32 272
use FILL  FILL_1__2306_
timestamp 1701859473
transform 1 0 4410 0 1 8590
box -12 -8 32 272
use FILL  FILL_1__2307_
timestamp 1701859473
transform 1 0 6270 0 1 9110
box -12 -8 32 272
use FILL  FILL_1__2308_
timestamp 1701859473
transform -1 0 8850 0 -1 6510
box -12 -8 32 272
use FILL  FILL_1__2309_
timestamp 1701859473
transform -1 0 8550 0 1 5990
box -12 -8 32 272
use FILL  FILL_1__2310_
timestamp 1701859473
transform -1 0 9050 0 -1 6510
box -12 -8 32 272
use FILL  FILL_1__2311_
timestamp 1701859473
transform -1 0 8610 0 -1 6510
box -12 -8 32 272
use FILL  FILL_1__2312_
timestamp 1701859473
transform -1 0 5510 0 -1 9630
box -12 -8 32 272
use FILL  FILL_1__2313_
timestamp 1701859473
transform -1 0 1790 0 1 8590
box -12 -8 32 272
use FILL  FILL_1__2314_
timestamp 1701859473
transform 1 0 1390 0 -1 8590
box -12 -8 32 272
use FILL  FILL_1__2315_
timestamp 1701859473
transform 1 0 1830 0 -1 8590
box -12 -8 32 272
use FILL  FILL_1__2316_
timestamp 1701859473
transform -1 0 4190 0 1 8590
box -12 -8 32 272
use FILL  FILL_1__2317_
timestamp 1701859473
transform 1 0 4650 0 1 8590
box -12 -8 32 272
use FILL  FILL_1__2318_
timestamp 1701859473
transform 1 0 6750 0 1 9110
box -12 -8 32 272
use FILL  FILL_1__2319_
timestamp 1701859473
transform -1 0 11070 0 1 4430
box -12 -8 32 272
use FILL  FILL_1__2320_
timestamp 1701859473
transform 1 0 5050 0 1 3910
box -12 -8 32 272
use FILL  FILL_1__2321_
timestamp 1701859473
transform 1 0 6470 0 1 3910
box -12 -8 32 272
use FILL  FILL_1__2322_
timestamp 1701859473
transform -1 0 7850 0 1 3910
box -12 -8 32 272
use FILL  FILL_1__2323_
timestamp 1701859473
transform 1 0 7890 0 -1 4430
box -12 -8 32 272
use FILL  FILL_1__2324_
timestamp 1701859473
transform -1 0 11110 0 -1 2870
box -12 -8 32 272
use FILL  FILL_1__2325_
timestamp 1701859473
transform -1 0 8090 0 1 3910
box -12 -8 32 272
use FILL  FILL_1__2326_
timestamp 1701859473
transform -1 0 3130 0 -1 4950
box -12 -8 32 272
use FILL  FILL_1__2327_
timestamp 1701859473
transform -1 0 3330 0 -1 4950
box -12 -8 32 272
use FILL  FILL_1__2328_
timestamp 1701859473
transform 1 0 3810 0 -1 5470
box -12 -8 32 272
use FILL  FILL_1__2329_
timestamp 1701859473
transform 1 0 3570 0 -1 5470
box -12 -8 32 272
use FILL  FILL_1__2330_
timestamp 1701859473
transform 1 0 3710 0 1 4950
box -12 -8 32 272
use FILL  FILL_1__2331_
timestamp 1701859473
transform 1 0 4790 0 1 3910
box -12 -8 32 272
use FILL  FILL_1__2332_
timestamp 1701859473
transform -1 0 4130 0 1 4950
box -12 -8 32 272
use FILL  FILL_1__2333_
timestamp 1701859473
transform -1 0 11090 0 -1 4430
box -12 -8 32 272
use FILL  FILL_1__2334_
timestamp 1701859473
transform 1 0 8970 0 -1 4430
box -12 -8 32 272
use FILL  FILL_1__2335_
timestamp 1701859473
transform 1 0 5150 0 -1 5470
box -12 -8 32 272
use FILL  FILL_1__2336_
timestamp 1701859473
transform -1 0 5010 0 1 5990
box -12 -8 32 272
use FILL  FILL_1__2337_
timestamp 1701859473
transform 1 0 4510 0 1 3390
box -12 -8 32 272
use FILL  FILL_1__2338_
timestamp 1701859473
transform 1 0 3110 0 1 3390
box -12 -8 32 272
use FILL  FILL_1__2339_
timestamp 1701859473
transform 1 0 4690 0 1 3390
box -12 -8 32 272
use FILL  FILL_1__2340_
timestamp 1701859473
transform 1 0 4930 0 1 3390
box -12 -8 32 272
use FILL  FILL_1__2341_
timestamp 1701859473
transform -1 0 510 0 1 5990
box -12 -8 32 272
use FILL  FILL_1__2342_
timestamp 1701859473
transform 1 0 2610 0 1 5470
box -12 -8 32 272
use FILL  FILL_1__2343_
timestamp 1701859473
transform -1 0 4550 0 1 6510
box -12 -8 32 272
use FILL  FILL_1__2344_
timestamp 1701859473
transform -1 0 4830 0 1 5470
box -12 -8 32 272
use FILL  FILL_1__2345_
timestamp 1701859473
transform -1 0 4630 0 1 5470
box -12 -8 32 272
use FILL  FILL_1__2346_
timestamp 1701859473
transform -1 0 4790 0 -1 5990
box -12 -8 32 272
use FILL  FILL_1__2347_
timestamp 1701859473
transform -1 0 5650 0 -1 5990
box -12 -8 32 272
use FILL  FILL_1__2348_
timestamp 1701859473
transform 1 0 5210 0 -1 6510
box -12 -8 32 272
use FILL  FILL_1__2349_
timestamp 1701859473
transform -1 0 4990 0 -1 6510
box -12 -8 32 272
use FILL  FILL_1__2350_
timestamp 1701859473
transform -1 0 4410 0 -1 6510
box -12 -8 32 272
use FILL  FILL_1__2351_
timestamp 1701859473
transform 1 0 5550 0 1 7030
box -12 -8 32 272
use FILL  FILL_1__2352_
timestamp 1701859473
transform -1 0 5770 0 1 7030
box -12 -8 32 272
use FILL  FILL_1__2353_
timestamp 1701859473
transform -1 0 710 0 1 7030
box -12 -8 32 272
use FILL  FILL_1__2354_
timestamp 1701859473
transform 1 0 5410 0 -1 5990
box -12 -8 32 272
use FILL  FILL_1__2355_
timestamp 1701859473
transform 1 0 5310 0 1 7030
box -12 -8 32 272
use FILL  FILL_1__2356_
timestamp 1701859473
transform -1 0 4810 0 -1 7550
box -12 -8 32 272
use FILL  FILL_1__2357_
timestamp 1701859473
transform 1 0 4670 0 1 8070
box -12 -8 32 272
use FILL  FILL_1__2358_
timestamp 1701859473
transform 1 0 5150 0 1 8070
box -12 -8 32 272
use FILL  FILL_1__2359_
timestamp 1701859473
transform -1 0 5470 0 -1 8590
box -12 -8 32 272
use FILL  FILL_1__2360_
timestamp 1701859473
transform -1 0 710 0 -1 6510
box -12 -8 32 272
use FILL  FILL_1__2361_
timestamp 1701859473
transform -1 0 5210 0 1 5990
box -12 -8 32 272
use FILL  FILL_1__2362_
timestamp 1701859473
transform 1 0 5210 0 1 6510
box -12 -8 32 272
use FILL  FILL_1__2363_
timestamp 1701859473
transform 1 0 5230 0 -1 7030
box -12 -8 32 272
use FILL  FILL_1__2364_
timestamp 1701859473
transform 1 0 5230 0 -1 8070
box -12 -8 32 272
use FILL  FILL_1__2365_
timestamp 1701859473
transform 1 0 5470 0 -1 8070
box -12 -8 32 272
use FILL  FILL_1__2366_
timestamp 1701859473
transform -1 0 5690 0 -1 8070
box -12 -8 32 272
use FILL  FILL_1__2367_
timestamp 1701859473
transform 1 0 2650 0 -1 7550
box -12 -8 32 272
use FILL  FILL_1__2368_
timestamp 1701859473
transform -1 0 5490 0 -1 7030
box -12 -8 32 272
use FILL  FILL_1__2369_
timestamp 1701859473
transform 1 0 5190 0 1 7550
box -12 -8 32 272
use FILL  FILL_1__2370_
timestamp 1701859473
transform -1 0 5230 0 -1 8590
box -12 -8 32 272
use FILL  FILL_1__2371_
timestamp 1701859473
transform 1 0 5910 0 -1 9110
box -12 -8 32 272
use FILL  FILL_1__2372_
timestamp 1701859473
transform 1 0 6070 0 1 9110
box -12 -8 32 272
use FILL  FILL_1__2373_
timestamp 1701859473
transform -1 0 6150 0 -1 9630
box -12 -8 32 272
use FILL  FILL_1__2374_
timestamp 1701859473
transform 1 0 30 0 -1 9110
box -12 -8 32 272
use FILL  FILL_1__2375_
timestamp 1701859473
transform -1 0 4170 0 1 5470
box -12 -8 32 272
use FILL  FILL_1__2376_
timestamp 1701859473
transform 1 0 4510 0 -1 5990
box -12 -8 32 272
use FILL  FILL_1__2377_
timestamp 1701859473
transform -1 0 3930 0 -1 6510
box -12 -8 32 272
use FILL  FILL_1__2378_
timestamp 1701859473
transform 1 0 3670 0 -1 6510
box -12 -8 32 272
use FILL  FILL_1__2379_
timestamp 1701859473
transform -1 0 4990 0 1 6510
box -12 -8 32 272
use FILL  FILL_1__2380_
timestamp 1701859473
transform -1 0 4770 0 -1 8590
box -12 -8 32 272
use FILL  FILL_1__2381_
timestamp 1701859473
transform 1 0 3830 0 -1 8590
box -12 -8 32 272
use FILL  FILL_1__2382_
timestamp 1701859473
transform -1 0 4530 0 -1 8590
box -12 -8 32 272
use FILL  FILL_1__2383_
timestamp 1701859473
transform -1 0 5610 0 1 8590
box -12 -8 32 272
use FILL  FILL_1__2384_
timestamp 1701859473
transform -1 0 5830 0 1 8590
box -12 -8 32 272
use FILL  FILL_1__2385_
timestamp 1701859473
transform 1 0 1210 0 -1 10150
box -12 -8 32 272
use FILL  FILL_1__2386_
timestamp 1701859473
transform 1 0 5470 0 -1 7550
box -12 -8 32 272
use FILL  FILL_1__2387_
timestamp 1701859473
transform 1 0 5450 0 -1 9110
box -12 -8 32 272
use FILL  FILL_1__2388_
timestamp 1701859473
transform -1 0 5250 0 -1 9110
box -12 -8 32 272
use FILL  FILL_1__2389_
timestamp 1701859473
transform -1 0 5030 0 -1 9630
box -12 -8 32 272
use FILL  FILL_1__2390_
timestamp 1701859473
transform 1 0 5090 0 1 9630
box -12 -8 32 272
use FILL  FILL_1__2391_
timestamp 1701859473
transform -1 0 5310 0 1 9630
box -12 -8 32 272
use FILL  FILL_1__2392_
timestamp 1701859473
transform 1 0 1410 0 -1 10150
box -12 -8 32 272
use FILL  FILL_1__2393_
timestamp 1701859473
transform -1 0 5270 0 -1 7550
box -12 -8 32 272
use FILL  FILL_1__2394_
timestamp 1701859473
transform 1 0 5350 0 1 8590
box -12 -8 32 272
use FILL  FILL_1__2395_
timestamp 1701859473
transform -1 0 5710 0 -1 9110
box -12 -8 32 272
use FILL  FILL_1__2396_
timestamp 1701859473
transform 1 0 5630 0 1 9110
box -12 -8 32 272
use FILL  FILL_1__2397_
timestamp 1701859473
transform 1 0 5870 0 1 9110
box -12 -8 32 272
use FILL  FILL_1__2398_
timestamp 1701859473
transform 1 0 5690 0 -1 9630
box -12 -8 32 272
use FILL  FILL_1__2399_
timestamp 1701859473
transform -1 0 3130 0 -1 5470
box -12 -8 32 272
use FILL  FILL_1__2400_
timestamp 1701859473
transform -1 0 3310 0 1 5990
box -12 -8 32 272
use FILL  FILL_1__2401_
timestamp 1701859473
transform 1 0 3230 0 -1 6510
box -12 -8 32 272
use FILL  FILL_1__2402_
timestamp 1701859473
transform -1 0 2170 0 -1 4430
box -12 -8 32 272
use FILL  FILL_1__2403_
timestamp 1701859473
transform -1 0 2570 0 1 4430
box -12 -8 32 272
use FILL  FILL_1__2404_
timestamp 1701859473
transform -1 0 2890 0 -1 5470
box -12 -8 32 272
use FILL  FILL_1__2405_
timestamp 1701859473
transform 1 0 2270 0 -1 2870
box -12 -8 32 272
use FILL  FILL_1__2406_
timestamp 1701859473
transform 1 0 2970 0 -1 3390
box -12 -8 32 272
use FILL  FILL_1__2407_
timestamp 1701859473
transform -1 0 3110 0 1 5470
box -12 -8 32 272
use FILL  FILL_1__2408_
timestamp 1701859473
transform 1 0 730 0 -1 2870
box -12 -8 32 272
use FILL  FILL_1__2409_
timestamp 1701859473
transform 1 0 750 0 -1 3910
box -12 -8 32 272
use FILL  FILL_1__2410_
timestamp 1701859473
transform 1 0 1150 0 1 4430
box -12 -8 32 272
use FILL  FILL_1__2411_
timestamp 1701859473
transform -1 0 710 0 -1 4950
box -12 -8 32 272
use FILL  FILL_1__2412_
timestamp 1701859473
transform 1 0 2390 0 -1 5990
box -12 -8 32 272
use FILL  FILL_1__2413_
timestamp 1701859473
transform 1 0 2850 0 1 5470
box -12 -8 32 272
use FILL  FILL_1__2414_
timestamp 1701859473
transform 1 0 4010 0 -1 5470
box -12 -8 32 272
use FILL  FILL_1__2415_
timestamp 1701859473
transform -1 0 3950 0 1 7030
box -12 -8 32 272
use FILL  FILL_1__2416_
timestamp 1701859473
transform 1 0 3910 0 1 4950
box -12 -8 32 272
use FILL  FILL_1__2417_
timestamp 1701859473
transform 1 0 4250 0 -1 5470
box -12 -8 32 272
use FILL  FILL_1__2418_
timestamp 1701859473
transform -1 0 1510 0 -1 4950
box -12 -8 32 272
use FILL  FILL_1__2419_
timestamp 1701859473
transform 1 0 2090 0 1 4430
box -12 -8 32 272
use FILL  FILL_1__2420_
timestamp 1701859473
transform 1 0 3750 0 1 5990
box -12 -8 32 272
use FILL  FILL_1__2421_
timestamp 1701859473
transform -1 0 3530 0 1 5990
box -12 -8 32 272
use FILL  FILL_1__2422_
timestamp 1701859473
transform -1 0 3410 0 -1 5990
box -12 -8 32 272
use FILL  FILL_1__2423_
timestamp 1701859473
transform -1 0 3630 0 -1 5990
box -12 -8 32 272
use FILL  FILL_1__2424_
timestamp 1701859473
transform 1 0 3170 0 -1 5990
box -12 -8 32 272
use FILL  FILL_1__2425_
timestamp 1701859473
transform 1 0 4310 0 1 5990
box -12 -8 32 272
use FILL  FILL_1__2426_
timestamp 1701859473
transform 1 0 3910 0 -1 7030
box -12 -8 32 272
use FILL  FILL_1__2427_
timestamp 1701859473
transform 1 0 4730 0 1 5990
box -12 -8 32 272
use FILL  FILL_1__2428_
timestamp 1701859473
transform 1 0 4490 0 1 5990
box -12 -8 32 272
use FILL  FILL_1__2429_
timestamp 1701859473
transform -1 0 4170 0 -1 6510
box -12 -8 32 272
use FILL  FILL_1__2430_
timestamp 1701859473
transform 1 0 4730 0 1 6510
box -12 -8 32 272
use FILL  FILL_1__2431_
timestamp 1701859473
transform -1 0 4830 0 -1 7030
box -12 -8 32 272
use FILL  FILL_1__2432_
timestamp 1701859473
transform 1 0 5050 0 -1 7030
box -12 -8 32 272
use FILL  FILL_1__2433_
timestamp 1701859473
transform -1 0 4310 0 -1 8070
box -12 -8 32 272
use FILL  FILL_1__2434_
timestamp 1701859473
transform 1 0 4790 0 1 7550
box -12 -8 32 272
use FILL  FILL_1__2435_
timestamp 1701859473
transform 1 0 4130 0 1 7030
box -12 -8 32 272
use FILL  FILL_1__2436_
timestamp 1701859473
transform -1 0 4570 0 -1 7550
box -12 -8 32 272
use FILL  FILL_1__2437_
timestamp 1701859473
transform -1 0 4550 0 -1 8070
box -12 -8 32 272
use FILL  FILL_1__2438_
timestamp 1701859473
transform -1 0 4790 0 -1 8070
box -12 -8 32 272
use FILL  FILL_1__2439_
timestamp 1701859473
transform -1 0 5030 0 -1 8070
box -12 -8 32 272
use FILL  FILL_1__2440_
timestamp 1701859473
transform 1 0 4570 0 1 10150
box -12 -8 32 272
use FILL  FILL_1__2441_
timestamp 1701859473
transform 1 0 3850 0 -1 7550
box -12 -8 32 272
use FILL  FILL_1__2442_
timestamp 1701859473
transform -1 0 4070 0 -1 8070
box -12 -8 32 272
use FILL  FILL_1__2443_
timestamp 1701859473
transform -1 0 3850 0 1 8070
box -12 -8 32 272
use FILL  FILL_1__2444_
timestamp 1701859473
transform 1 0 3590 0 1 8070
box -12 -8 32 272
use FILL  FILL_1__2445_
timestamp 1701859473
transform -1 0 4570 0 1 7550
box -12 -8 32 272
use FILL  FILL_1__2446_
timestamp 1701859473
transform 1 0 4490 0 1 8070
box -12 -8 32 272
use FILL  FILL_1__2447_
timestamp 1701859473
transform 1 0 4230 0 1 9110
box -12 -8 32 272
use FILL  FILL_1__2448_
timestamp 1701859473
transform 1 0 4890 0 1 9110
box -12 -8 32 272
use FILL  FILL_1__2449_
timestamp 1701859473
transform 1 0 5150 0 1 9110
box -12 -8 32 272
use FILL  FILL_1__2450_
timestamp 1701859473
transform 1 0 5390 0 1 9110
box -12 -8 32 272
use FILL  FILL_1__2451_
timestamp 1701859473
transform -1 0 5270 0 -1 9630
box -12 -8 32 272
use FILL  FILL_1__2452_
timestamp 1701859473
transform -1 0 5190 0 -1 10670
box -12 -8 32 272
use FILL  FILL_1__2453_
timestamp 1701859473
transform 1 0 3730 0 -1 10150
box -12 -8 32 272
use FILL  FILL_1__2454_
timestamp 1701859473
transform 1 0 3850 0 1 7550
box -12 -8 32 272
use FILL  FILL_1__2455_
timestamp 1701859473
transform 1 0 3810 0 -1 8070
box -12 -8 32 272
use FILL  FILL_1__2456_
timestamp 1701859473
transform -1 0 3590 0 -1 8070
box -12 -8 32 272
use FILL  FILL_1__2457_
timestamp 1701859473
transform 1 0 3350 0 1 8070
box -12 -8 32 272
use FILL  FILL_1__2458_
timestamp 1701859473
transform -1 0 4290 0 -1 8590
box -12 -8 32 272
use FILL  FILL_1__2459_
timestamp 1701859473
transform -1 0 4450 0 -1 11190
box -12 -8 32 272
use FILL  FILL_1__2460_
timestamp 1701859473
transform 1 0 4090 0 -1 10670
box -12 -8 32 272
use FILL  FILL_1__2461_
timestamp 1701859473
transform 1 0 4270 0 -1 9110
box -12 -8 32 272
use FILL  FILL_1__2462_
timestamp 1701859473
transform -1 0 4530 0 -1 9110
box -12 -8 32 272
use FILL  FILL_1__2463_
timestamp 1701859473
transform -1 0 4770 0 -1 9110
box -12 -8 32 272
use FILL  FILL_1__2464_
timestamp 1701859473
transform -1 0 5010 0 -1 9110
box -12 -8 32 272
use FILL  FILL_1__2465_
timestamp 1701859473
transform -1 0 4870 0 -1 11190
box -12 -8 32 272
use FILL  FILL_1__2466_
timestamp 1701859473
transform -1 0 3950 0 -1 10150
box -12 -8 32 272
use FILL  FILL_1__2467_
timestamp 1701859473
transform -1 0 4050 0 -1 9630
box -12 -8 32 272
use FILL  FILL_1__2468_
timestamp 1701859473
transform -1 0 4310 0 -1 9630
box -12 -8 32 272
use FILL  FILL_1__2469_
timestamp 1701859473
transform -1 0 4170 0 1 9630
box -12 -8 32 272
use FILL  FILL_1__2470_
timestamp 1701859473
transform -1 0 4410 0 1 9630
box -12 -8 32 272
use FILL  FILL_1__2471_
timestamp 1701859473
transform -1 0 4990 0 -1 10670
box -12 -8 32 272
use FILL  FILL_1__2472_
timestamp 1701859473
transform 1 0 3950 0 1 9630
box -12 -8 32 272
use FILL  FILL_1__2473_
timestamp 1701859473
transform 1 0 4510 0 -1 9630
box -12 -8 32 272
use FILL  FILL_1__2474_
timestamp 1701859473
transform -1 0 4790 0 -1 9630
box -12 -8 32 272
use FILL  FILL_1__2475_
timestamp 1701859473
transform 1 0 4630 0 1 9630
box -12 -8 32 272
use FILL  FILL_1__2476_
timestamp 1701859473
transform -1 0 4870 0 1 9630
box -12 -8 32 272
use FILL  FILL_1__2477_
timestamp 1701859473
transform 1 0 4810 0 1 10670
box -12 -8 32 272
use FILL  FILL_1__2478_
timestamp 1701859473
transform 1 0 3050 0 1 5990
box -12 -8 32 272
use FILL  FILL_1__2479_
timestamp 1701859473
transform -1 0 2610 0 1 5990
box -12 -8 32 272
use FILL  FILL_1__2480_
timestamp 1701859473
transform -1 0 2630 0 -1 5990
box -12 -8 32 272
use FILL  FILL_1__2481_
timestamp 1701859473
transform -1 0 2870 0 -1 5990
box -12 -8 32 272
use FILL  FILL_1__2482_
timestamp 1701859473
transform 1 0 1450 0 -1 5990
box -12 -8 32 272
use FILL  FILL_1__2483_
timestamp 1701859473
transform 1 0 2270 0 1 6510
box -12 -8 32 272
use FILL  FILL_1__2484_
timestamp 1701859473
transform -1 0 1890 0 1 6510
box -12 -8 32 272
use FILL  FILL_1__2485_
timestamp 1701859473
transform -1 0 2090 0 1 6510
box -12 -8 32 272
use FILL  FILL_1__2486_
timestamp 1701859473
transform 1 0 2290 0 -1 7030
box -12 -8 32 272
use FILL  FILL_1__2487_
timestamp 1701859473
transform 1 0 2050 0 -1 7030
box -12 -8 32 272
use FILL  FILL_1__2488_
timestamp 1701859473
transform -1 0 1850 0 -1 7030
box -12 -8 32 272
use FILL  FILL_1__2489_
timestamp 1701859473
transform 1 0 1350 0 -1 7030
box -12 -8 32 272
use FILL  FILL_1__2490_
timestamp 1701859473
transform -1 0 950 0 1 5470
box -12 -8 32 272
use FILL  FILL_1__2491_
timestamp 1701859473
transform 1 0 1150 0 1 5470
box -12 -8 32 272
use FILL  FILL_1__2492_
timestamp 1701859473
transform -1 0 2010 0 -1 6510
box -12 -8 32 272
use FILL  FILL_1__2493_
timestamp 1701859473
transform 1 0 1890 0 1 5990
box -12 -8 32 272
use FILL  FILL_1__2494_
timestamp 1701859473
transform -1 0 1450 0 1 5990
box -12 -8 32 272
use FILL  FILL_1__2495_
timestamp 1701859473
transform 1 0 1190 0 1 5990
box -12 -8 32 272
use FILL  FILL_1__2496_
timestamp 1701859473
transform 1 0 1590 0 -1 7030
box -12 -8 32 272
use FILL  FILL_1__2497_
timestamp 1701859473
transform -1 0 1790 0 -1 7550
box -12 -8 32 272
use FILL  FILL_1__2498_
timestamp 1701859473
transform 1 0 730 0 1 8070
box -12 -8 32 272
use FILL  FILL_1__2499_
timestamp 1701859473
transform 1 0 2410 0 1 7550
box -12 -8 32 272
use FILL  FILL_1__2500_
timestamp 1701859473
transform 1 0 1830 0 1 7550
box -12 -8 32 272
use FILL  FILL_1__2501_
timestamp 1701859473
transform 1 0 1610 0 1 7550
box -12 -8 32 272
use FILL  FILL_1__2502_
timestamp 1701859473
transform -1 0 1150 0 1 7550
box -12 -8 32 272
use FILL  FILL_1__2503_
timestamp 1701859473
transform -1 0 1390 0 1 8070
box -12 -8 32 272
use FILL  FILL_1__2504_
timestamp 1701859473
transform -1 0 1810 0 1 8070
box -12 -8 32 272
use FILL  FILL_1__2505_
timestamp 1701859473
transform 1 0 1150 0 1 8070
box -12 -8 32 272
use FILL  FILL_1__2506_
timestamp 1701859473
transform -1 0 1670 0 -1 8070
box -12 -8 32 272
use FILL  FILL_1__2507_
timestamp 1701859473
transform 1 0 1410 0 -1 8070
box -12 -8 32 272
use FILL  FILL_1__2508_
timestamp 1701859473
transform 1 0 930 0 1 8070
box -12 -8 32 272
use FILL  FILL_1__2509_
timestamp 1701859473
transform 1 0 490 0 -1 8590
box -12 -8 32 272
use FILL  FILL_1__2510_
timestamp 1701859473
transform -1 0 1430 0 1 9110
box -12 -8 32 272
use FILL  FILL_1__2511_
timestamp 1701859473
transform -1 0 1370 0 -1 9630
box -12 -8 32 272
use FILL  FILL_1__2512_
timestamp 1701859473
transform 1 0 930 0 -1 9630
box -12 -8 32 272
use FILL  FILL_1__2513_
timestamp 1701859473
transform -1 0 930 0 1 8590
box -12 -8 32 272
use FILL  FILL_1__2514_
timestamp 1701859473
transform 1 0 2010 0 -1 8590
box -12 -8 32 272
use FILL  FILL_1__2515_
timestamp 1701859473
transform 1 0 1130 0 -1 9110
box -12 -8 32 272
use FILL  FILL_1__2516_
timestamp 1701859473
transform -1 0 970 0 1 9110
box -12 -8 32 272
use FILL  FILL_1__2517_
timestamp 1701859473
transform -1 0 730 0 1 9110
box -12 -8 32 272
use FILL  FILL_1__2518_
timestamp 1701859473
transform 1 0 1590 0 -1 9630
box -12 -8 32 272
use FILL  FILL_1__2519_
timestamp 1701859473
transform 1 0 1690 0 1 9630
box -12 -8 32 272
use FILL  FILL_1__2520_
timestamp 1701859473
transform -1 0 2530 0 -1 9110
box -12 -8 32 272
use FILL  FILL_1__2521_
timestamp 1701859473
transform 1 0 2270 0 -1 9110
box -12 -8 32 272
use FILL  FILL_1__2522_
timestamp 1701859473
transform -1 0 1890 0 1 9630
box -12 -8 32 272
use FILL  FILL_1__2523_
timestamp 1701859473
transform -1 0 2110 0 1 9630
box -12 -8 32 272
use FILL  FILL_1__2524_
timestamp 1701859473
transform -1 0 1850 0 -1 9110
box -12 -8 32 272
use FILL  FILL_1__2525_
timestamp 1701859473
transform 1 0 730 0 -1 8590
box -12 -8 32 272
use FILL  FILL_1__2526_
timestamp 1701859473
transform -1 0 1630 0 -1 8590
box -12 -8 32 272
use FILL  FILL_1__2527_
timestamp 1701859473
transform -1 0 1170 0 -1 8590
box -12 -8 32 272
use FILL  FILL_1__2528_
timestamp 1701859473
transform -1 0 950 0 -1 8590
box -12 -8 32 272
use FILL  FILL_1__2529_
timestamp 1701859473
transform -1 0 1190 0 1 9110
box -12 -8 32 272
use FILL  FILL_1__2530_
timestamp 1701859473
transform -1 0 7450 0 -1 6510
box -12 -8 32 272
use FILL  FILL_1__2531_
timestamp 1701859473
transform 1 0 7870 0 1 7550
box -12 -8 32 272
use FILL  FILL_1__2532_
timestamp 1701859473
transform -1 0 9770 0 1 2870
box -12 -8 32 272
use FILL  FILL_1__2533_
timestamp 1701859473
transform -1 0 8850 0 1 4430
box -12 -8 32 272
use FILL  FILL_1__2534_
timestamp 1701859473
transform -1 0 9250 0 -1 5470
box -12 -8 32 272
use FILL  FILL_1__2535_
timestamp 1701859473
transform 1 0 30 0 -1 4950
box -12 -8 32 272
use FILL  FILL_1__2536_
timestamp 1701859473
transform 1 0 590 0 1 4950
box -12 -8 32 272
use FILL  FILL_1__2537_
timestamp 1701859473
transform 1 0 730 0 1 3390
box -12 -8 32 272
use FILL  FILL_1__2538_
timestamp 1701859473
transform -1 0 290 0 -1 3910
box -12 -8 32 272
use FILL  FILL_1__2539_
timestamp 1701859473
transform -1 0 50 0 1 4950
box -12 -8 32 272
use FILL  FILL_1__2540_
timestamp 1701859473
transform 1 0 2990 0 1 2350
box -12 -8 32 272
use FILL  FILL_1__2541_
timestamp 1701859473
transform -1 0 3250 0 1 2870
box -12 -8 32 272
use FILL  FILL_1__2542_
timestamp 1701859473
transform -1 0 2250 0 -1 6510
box -12 -8 32 272
use FILL  FILL_1__2543_
timestamp 1701859473
transform 1 0 810 0 1 4950
box -12 -8 32 272
use FILL  FILL_1__2544_
timestamp 1701859473
transform 1 0 1370 0 1 4430
box -12 -8 32 272
use FILL  FILL_1__2545_
timestamp 1701859473
transform 1 0 1230 0 -1 5470
box -12 -8 32 272
use FILL  FILL_1__2546_
timestamp 1701859473
transform -1 0 1970 0 -1 5470
box -12 -8 32 272
use FILL  FILL_1__2547_
timestamp 1701859473
transform 1 0 1910 0 -1 4430
box -12 -8 32 272
use FILL  FILL_1__2548_
timestamp 1701859473
transform 1 0 1030 0 1 4950
box -12 -8 32 272
use FILL  FILL_1__2549_
timestamp 1701859473
transform 1 0 1250 0 1 4950
box -12 -8 32 272
use FILL  FILL_1__2550_
timestamp 1701859473
transform -1 0 1730 0 -1 5470
box -12 -8 32 272
use FILL  FILL_1__2551_
timestamp 1701859473
transform 1 0 2510 0 -1 9630
box -12 -8 32 272
use FILL  FILL_1__2552_
timestamp 1701859473
transform 1 0 3350 0 -1 5470
box -12 -8 32 272
use FILL  FILL_1__2553_
timestamp 1701859473
transform -1 0 2730 0 -1 6510
box -12 -8 32 272
use FILL  FILL_1__2554_
timestamp 1701859473
transform -1 0 3190 0 1 6510
box -12 -8 32 272
use FILL  FILL_1__2555_
timestamp 1701859473
transform -1 0 3430 0 1 6510
box -12 -8 32 272
use FILL  FILL_1__2556_
timestamp 1701859473
transform -1 0 2750 0 1 6510
box -12 -8 32 272
use FILL  FILL_1__2557_
timestamp 1701859473
transform 1 0 2450 0 -1 6510
box -12 -8 32 272
use FILL  FILL_1__2558_
timestamp 1701859473
transform 1 0 3190 0 -1 7550
box -12 -8 32 272
use FILL  FILL_1__2559_
timestamp 1701859473
transform 1 0 3390 0 -1 7550
box -12 -8 32 272
use FILL  FILL_1__2560_
timestamp 1701859473
transform -1 0 3450 0 1 7030
box -12 -8 32 272
use FILL  FILL_1__2561_
timestamp 1701859473
transform -1 0 1470 0 1 4950
box -12 -8 32 272
use FILL  FILL_1__2562_
timestamp 1701859473
transform 1 0 3190 0 1 7030
box -12 -8 32 272
use FILL  FILL_1__2563_
timestamp 1701859473
transform 1 0 3750 0 1 5470
box -12 -8 32 272
use FILL  FILL_1__2564_
timestamp 1701859473
transform -1 0 3630 0 1 6510
box -12 -8 32 272
use FILL  FILL_1__2565_
timestamp 1701859473
transform 1 0 3690 0 1 7030
box -12 -8 32 272
use FILL  FILL_1__2566_
timestamp 1701859473
transform 1 0 3150 0 1 7550
box -12 -8 32 272
use FILL  FILL_1__2567_
timestamp 1701859473
transform 1 0 3110 0 -1 8070
box -12 -8 32 272
use FILL  FILL_1__2568_
timestamp 1701859473
transform -1 0 2930 0 -1 8590
box -12 -8 32 272
use FILL  FILL_1__2569_
timestamp 1701859473
transform 1 0 2690 0 -1 8590
box -12 -8 32 272
use FILL  FILL_1__2570_
timestamp 1701859473
transform 1 0 2870 0 -1 8070
box -12 -8 32 272
use FILL  FILL_1__2571_
timestamp 1701859473
transform -1 0 3830 0 -1 9630
box -12 -8 32 272
use FILL  FILL_1__2572_
timestamp 1701859473
transform -1 0 3850 0 -1 5990
box -12 -8 32 272
use FILL  FILL_1__2573_
timestamp 1701859473
transform -1 0 3710 0 -1 7030
box -12 -8 32 272
use FILL  FILL_1__2574_
timestamp 1701859473
transform 1 0 3430 0 -1 6510
box -12 -8 32 272
use FILL  FILL_1__2575_
timestamp 1701859473
transform 1 0 3330 0 -1 8070
box -12 -8 32 272
use FILL  FILL_1__2576_
timestamp 1701859473
transform -1 0 3370 0 -1 8590
box -12 -8 32 272
use FILL  FILL_1__2577_
timestamp 1701859473
transform 1 0 3250 0 1 9110
box -12 -8 32 272
use FILL  FILL_1__2578_
timestamp 1701859473
transform 1 0 3750 0 1 9110
box -12 -8 32 272
use FILL  FILL_1__2579_
timestamp 1701859473
transform -1 0 2730 0 -1 9630
box -12 -8 32 272
use FILL  FILL_1__2580_
timestamp 1701859473
transform -1 0 4090 0 -1 9110
box -12 -8 32 272
use FILL  FILL_1__2581_
timestamp 1701859473
transform -1 0 4010 0 1 9110
box -12 -8 32 272
use FILL  FILL_1__2582_
timestamp 1701859473
transform 1 0 3510 0 1 9110
box -12 -8 32 272
use FILL  FILL_1__2583_
timestamp 1701859473
transform 1 0 3010 0 1 9110
box -12 -8 32 272
use FILL  FILL_1__2584_
timestamp 1701859473
transform 1 0 2770 0 1 9110
box -12 -8 32 272
use FILL  FILL_1__2585_
timestamp 1701859473
transform 1 0 3870 0 -1 9110
box -12 -8 32 272
use FILL  FILL_1__2586_
timestamp 1701859473
transform 1 0 3030 0 1 9630
box -12 -8 32 272
use FILL  FILL_1__2587_
timestamp 1701859473
transform 1 0 3610 0 -1 9110
box -12 -8 32 272
use FILL  FILL_1__2588_
timestamp 1701859473
transform 1 0 3210 0 1 8590
box -12 -8 32 272
use FILL  FILL_1__2589_
timestamp 1701859473
transform 1 0 3050 0 -1 10150
box -12 -8 32 272
use FILL  FILL_1__2590_
timestamp 1701859473
transform 1 0 2790 0 -1 10150
box -12 -8 32 272
use FILL  FILL_1__2591_
timestamp 1701859473
transform -1 0 3550 0 -1 11190
box -12 -8 32 272
use FILL  FILL_1__2592_
timestamp 1701859473
transform -1 0 3610 0 -1 9630
box -12 -8 32 272
use FILL  FILL_1__2593_
timestamp 1701859473
transform -1 0 3130 0 -1 9630
box -12 -8 32 272
use FILL  FILL_1__2594_
timestamp 1701859473
transform -1 0 3290 0 -1 10150
box -12 -8 32 272
use FILL  FILL_1__2595_
timestamp 1701859473
transform 1 0 3010 0 -1 11190
box -12 -8 32 272
use FILL  FILL_1__2596_
timestamp 1701859473
transform 1 0 3290 0 -1 11190
box -12 -8 32 272
use FILL  FILL_1__2597_
timestamp 1701859473
transform 1 0 2750 0 -1 10670
box -12 -8 32 272
use FILL  FILL_1__2598_
timestamp 1701859473
transform -1 0 3490 0 1 9630
box -12 -8 32 272
use FILL  FILL_1__2599_
timestamp 1701859473
transform -1 0 3270 0 1 9630
box -12 -8 32 272
use FILL  FILL_1__2600_
timestamp 1701859473
transform -1 0 2990 0 1 10150
box -12 -8 32 272
use FILL  FILL_1__2601_
timestamp 1701859473
transform 1 0 2950 0 -1 10670
box -12 -8 32 272
use FILL  FILL_1__2602_
timestamp 1701859473
transform -1 0 3210 0 -1 10670
box -12 -8 32 272
use FILL  FILL_1__2603_
timestamp 1701859473
transform 1 0 3410 0 -1 10670
box -12 -8 32 272
use FILL  FILL_1__2604_
timestamp 1701859473
transform 1 0 3210 0 1 10150
box -12 -8 32 272
use FILL  FILL_1__2605_
timestamp 1701859473
transform 1 0 2330 0 1 10670
box -12 -8 32 272
use FILL  FILL_1__2606_
timestamp 1701859473
transform 1 0 2530 0 1 10670
box -12 -8 32 272
use FILL  FILL_1__2607_
timestamp 1701859473
transform -1 0 2770 0 1 10670
box -12 -8 32 272
use FILL  FILL_1__2608_
timestamp 1701859473
transform -1 0 3730 0 1 9630
box -12 -8 32 272
use FILL  FILL_1__2609_
timestamp 1701859473
transform -1 0 2350 0 1 9630
box -12 -8 32 272
use FILL  FILL_1__2610_
timestamp 1701859473
transform -1 0 2570 0 -1 10150
box -12 -8 32 272
use FILL  FILL_1__2611_
timestamp 1701859473
transform -1 0 2290 0 -1 10670
box -12 -8 32 272
use FILL  FILL_1__2612_
timestamp 1701859473
transform 1 0 2510 0 -1 10670
box -12 -8 32 272
use FILL  FILL_1__2613_
timestamp 1701859473
transform 1 0 1830 0 1 10670
box -12 -8 32 272
use FILL  FILL_1__2614_
timestamp 1701859473
transform 1 0 1830 0 -1 10670
box -12 -8 32 272
use FILL  FILL_1__2615_
timestamp 1701859473
transform -1 0 2350 0 -1 11190
box -12 -8 32 272
use FILL  FILL_1__2616_
timestamp 1701859473
transform -1 0 3370 0 -1 9630
box -12 -8 32 272
use FILL  FILL_1__2617_
timestamp 1701859473
transform 1 0 2270 0 -1 9630
box -12 -8 32 272
use FILL  FILL_1__2618_
timestamp 1701859473
transform -1 0 2550 0 1 10150
box -12 -8 32 272
use FILL  FILL_1__2619_
timestamp 1701859473
transform 1 0 2050 0 1 10670
box -12 -8 32 272
use FILL  FILL_1__2620_
timestamp 1701859473
transform 1 0 2090 0 -1 11190
box -12 -8 32 272
use FILL  FILL_1__2621_
timestamp 1701859473
transform -1 0 1370 0 1 5470
box -12 -8 32 272
use FILL  FILL_1__2622_
timestamp 1701859473
transform -1 0 1210 0 -1 5990
box -12 -8 32 272
use FILL  FILL_1__2623_
timestamp 1701859473
transform 1 0 2430 0 -1 5470
box -12 -8 32 272
use FILL  FILL_1__2624_
timestamp 1701859473
transform -1 0 2390 0 1 5470
box -12 -8 32 272
use FILL  FILL_1__2625_
timestamp 1701859473
transform 1 0 2190 0 -1 5470
box -12 -8 32 272
use FILL  FILL_1__2626_
timestamp 1701859473
transform -1 0 930 0 -1 5470
box -12 -8 32 272
use FILL  FILL_1__2627_
timestamp 1701859473
transform -1 0 1450 0 1 3910
box -12 -8 32 272
use FILL  FILL_1__2628_
timestamp 1701859473
transform 1 0 1130 0 1 3910
box -12 -8 32 272
use FILL  FILL_1__2629_
timestamp 1701859473
transform -1 0 730 0 -1 5470
box -12 -8 32 272
use FILL  FILL_1__2630_
timestamp 1701859473
transform 1 0 710 0 -1 5990
box -12 -8 32 272
use FILL  FILL_1__2631_
timestamp 1701859473
transform -1 0 710 0 1 5990
box -12 -8 32 272
use FILL  FILL_1__2632_
timestamp 1701859473
transform 1 0 2090 0 1 10150
box -12 -8 32 272
use FILL  FILL_1__2633_
timestamp 1701859473
transform -1 0 2330 0 1 10150
box -12 -8 32 272
use FILL  FILL_1__2634_
timestamp 1701859473
transform 1 0 2290 0 -1 10150
box -12 -8 32 272
use FILL  FILL_1__2635_
timestamp 1701859473
transform 1 0 2070 0 -1 10150
box -12 -8 32 272
use FILL  FILL_1__2636_
timestamp 1701859473
transform -1 0 710 0 -1 10150
box -12 -8 32 272
use FILL  FILL_1__2637_
timestamp 1701859473
transform -1 0 510 0 1 6510
box -12 -8 32 272
use FILL  FILL_1__2638_
timestamp 1701859473
transform -1 0 290 0 1 6510
box -12 -8 32 272
use FILL  FILL_1__2639_
timestamp 1701859473
transform -1 0 270 0 -1 6510
box -12 -8 32 272
use FILL  FILL_1__2640_
timestamp 1701859473
transform -1 0 270 0 1 5990
box -12 -8 32 272
use FILL  FILL_1__2641_
timestamp 1701859473
transform 1 0 30 0 -1 7550
box -12 -8 32 272
use FILL  FILL_1__2642_
timestamp 1701859473
transform -1 0 370 0 1 4950
box -12 -8 32 272
use FILL  FILL_1__2643_
timestamp 1701859473
transform -1 0 2510 0 1 6510
box -12 -8 32 272
use FILL  FILL_1__2644_
timestamp 1701859473
transform 1 0 2550 0 -1 7030
box -12 -8 32 272
use FILL  FILL_1__2645_
timestamp 1701859473
transform 1 0 2730 0 1 7030
box -12 -8 32 272
use FILL  FILL_1__2646_
timestamp 1701859473
transform 1 0 2030 0 1 7030
box -12 -8 32 272
use FILL  FILL_1__2647_
timestamp 1701859473
transform 1 0 710 0 1 7550
box -12 -8 32 272
use FILL  FILL_1__2648_
timestamp 1701859473
transform 1 0 250 0 1 7550
box -12 -8 32 272
use FILL  FILL_1__2649_
timestamp 1701859473
transform 1 0 230 0 -1 7550
box -12 -8 32 272
use FILL  FILL_1__2650_
timestamp 1701859473
transform -1 0 710 0 -1 7550
box -12 -8 32 272
use FILL  FILL_1__2651_
timestamp 1701859473
transform 1 0 450 0 -1 7550
box -12 -8 32 272
use FILL  FILL_1__2652_
timestamp 1701859473
transform 1 0 450 0 1 7030
box -12 -8 32 272
use FILL  FILL_1__2653_
timestamp 1701859473
transform 1 0 30 0 1 7550
box -12 -8 32 272
use FILL  FILL_1__2654_
timestamp 1701859473
transform -1 0 510 0 1 7550
box -12 -8 32 272
use FILL  FILL_1__2655_
timestamp 1701859473
transform 1 0 1830 0 1 7030
box -12 -8 32 272
use FILL  FILL_1__2656_
timestamp 1701859473
transform 1 0 1470 0 -1 5470
box -12 -8 32 272
use FILL  FILL_1__2657_
timestamp 1701859473
transform -1 0 1670 0 1 5990
box -12 -8 32 272
use FILL  FILL_1__2658_
timestamp 1701859473
transform -1 0 2150 0 1 5470
box -12 -8 32 272
use FILL  FILL_1__2659_
timestamp 1701859473
transform 1 0 1910 0 -1 5990
box -12 -8 32 272
use FILL  FILL_1__2660_
timestamp 1701859473
transform -1 0 1910 0 1 5470
box -12 -8 32 272
use FILL  FILL_1__2661_
timestamp 1701859473
transform -1 0 1590 0 1 5470
box -12 -8 32 272
use FILL  FILL_1__2662_
timestamp 1701859473
transform 1 0 690 0 1 5470
box -12 -8 32 272
use FILL  FILL_1__2663_
timestamp 1701859473
transform -1 0 970 0 -1 5990
box -12 -8 32 272
use FILL  FILL_1__2664_
timestamp 1701859473
transform 1 0 690 0 -1 7030
box -12 -8 32 272
use FILL  FILL_1__2665_
timestamp 1701859473
transform 1 0 1150 0 -1 7030
box -12 -8 32 272
use FILL  FILL_1__2666_
timestamp 1701859473
transform 1 0 1350 0 1 7030
box -12 -8 32 272
use FILL  FILL_1__2667_
timestamp 1701859473
transform 1 0 890 0 -1 7030
box -12 -8 32 272
use FILL  FILL_1__2668_
timestamp 1701859473
transform -1 0 2690 0 1 7550
box -12 -8 32 272
use FILL  FILL_1__2669_
timestamp 1701859473
transform 1 0 2630 0 -1 8070
box -12 -8 32 272
use FILL  FILL_1__2670_
timestamp 1701859473
transform 1 0 1890 0 -1 8070
box -12 -8 32 272
use FILL  FILL_1__2671_
timestamp 1701859473
transform -1 0 1390 0 1 7550
box -12 -8 32 272
use FILL  FILL_1__2672_
timestamp 1701859473
transform 1 0 1110 0 -1 7550
box -12 -8 32 272
use FILL  FILL_1__2673_
timestamp 1701859473
transform -1 0 1310 0 -1 7550
box -12 -8 32 272
use FILL  FILL_1__2674_
timestamp 1701859473
transform 1 0 1590 0 1 7030
box -12 -8 32 272
use FILL  FILL_1__2675_
timestamp 1701859473
transform 1 0 1530 0 -1 7550
box -12 -8 32 272
use FILL  FILL_1__2676_
timestamp 1701859473
transform -1 0 1970 0 -1 7550
box -12 -8 32 272
use FILL  FILL_1__2677_
timestamp 1701859473
transform 1 0 2370 0 -1 8070
box -12 -8 32 272
use FILL  FILL_1__2678_
timestamp 1701859473
transform -1 0 2150 0 -1 8070
box -12 -8 32 272
use FILL  FILL_1__2679_
timestamp 1701859473
transform -1 0 1590 0 1 8070
box -12 -8 32 272
use FILL  FILL_1__2680_
timestamp 1701859473
transform -1 0 270 0 -1 8590
box -12 -8 32 272
use FILL  FILL_1__2681_
timestamp 1701859473
transform 1 0 890 0 -1 7550
box -12 -8 32 272
use FILL  FILL_1__2682_
timestamp 1701859473
transform -1 0 270 0 -1 8070
box -12 -8 32 272
use FILL  FILL_1__2683_
timestamp 1701859473
transform -1 0 50 0 -1 9630
box -12 -8 32 272
use FILL  FILL_1__2684_
timestamp 1701859473
transform -1 0 50 0 1 10150
box -12 -8 32 272
use FILL  FILL_1__2685_
timestamp 1701859473
transform 1 0 930 0 1 5990
box -12 -8 32 272
use FILL  FILL_1__2686_
timestamp 1701859473
transform 1 0 910 0 1 7550
box -12 -8 32 272
use FILL  FILL_1__2687_
timestamp 1701859473
transform -1 0 910 0 -1 10150
box -12 -8 32 272
use FILL  FILL_1__2688_
timestamp 1701859473
transform 1 0 30 0 -1 10150
box -12 -8 32 272
use FILL  FILL_1__2689_
timestamp 1701859473
transform 1 0 250 0 -1 9630
box -12 -8 32 272
use FILL  FILL_1__2690_
timestamp 1701859473
transform 1 0 250 0 1 9110
box -12 -8 32 272
use FILL  FILL_1__2691_
timestamp 1701859473
transform 1 0 2710 0 1 8590
box -12 -8 32 272
use FILL  FILL_1__2692_
timestamp 1701859473
transform 1 0 2470 0 1 8590
box -12 -8 32 272
use FILL  FILL_1__2693_
timestamp 1701859473
transform -1 0 1130 0 -1 9630
box -12 -8 32 272
use FILL  FILL_1__2694_
timestamp 1701859473
transform 1 0 710 0 -1 9630
box -12 -8 32 272
use FILL  FILL_1__2695_
timestamp 1701859473
transform 1 0 30 0 1 9630
box -12 -8 32 272
use FILL  FILL_1__2696_
timestamp 1701859473
transform -1 0 510 0 -1 10150
box -12 -8 32 272
use FILL  FILL_1__2697_
timestamp 1701859473
transform 1 0 250 0 -1 10150
box -12 -8 32 272
use FILL  FILL_1__2698_
timestamp 1701859473
transform 1 0 270 0 1 9630
box -12 -8 32 272
use FILL  FILL_1__2699_
timestamp 1701859473
transform 1 0 490 0 -1 9630
box -12 -8 32 272
use FILL  FILL_1__2700_
timestamp 1701859473
transform 1 0 510 0 1 9630
box -12 -8 32 272
use FILL  FILL_1__2701_
timestamp 1701859473
transform -1 0 730 0 -1 10670
box -12 -8 32 272
use FILL  FILL_1__2702_
timestamp 1701859473
transform 1 0 3450 0 1 8590
box -12 -8 32 272
use FILL  FILL_1__2703_
timestamp 1701859473
transform -1 0 2990 0 1 8590
box -12 -8 32 272
use FILL  FILL_1__2704_
timestamp 1701859473
transform -1 0 1470 0 1 9630
box -12 -8 32 272
use FILL  FILL_1__2705_
timestamp 1701859473
transform 1 0 1210 0 1 9630
box -12 -8 32 272
use FILL  FILL_1__2706_
timestamp 1701859473
transform 1 0 230 0 1 10150
box -12 -8 32 272
use FILL  FILL_1__2707_
timestamp 1701859473
transform -1 0 470 0 1 10150
box -12 -8 32 272
use FILL  FILL_1__2708_
timestamp 1701859473
transform 1 0 670 0 1 10150
box -12 -8 32 272
use FILL  FILL_1__2709_
timestamp 1701859473
transform -1 0 490 0 -1 10670
box -12 -8 32 272
use FILL  FILL_1__2710_
timestamp 1701859473
transform 1 0 1670 0 1 10150
box -12 -8 32 272
use FILL  FILL_1__2711_
timestamp 1701859473
transform 1 0 2210 0 1 8590
box -12 -8 32 272
use FILL  FILL_1__2712_
timestamp 1701859473
transform -1 0 1990 0 1 8590
box -12 -8 32 272
use FILL  FILL_1__2713_
timestamp 1701859473
transform -1 0 1850 0 -1 9630
box -12 -8 32 272
use FILL  FILL_1__2714_
timestamp 1701859473
transform 1 0 1610 0 -1 10150
box -12 -8 32 272
use FILL  FILL_1__2715_
timestamp 1701859473
transform 1 0 930 0 1 10150
box -12 -8 32 272
use FILL  FILL_1__2716_
timestamp 1701859473
transform 1 0 1170 0 1 10150
box -12 -8 32 272
use FILL  FILL_1__2717_
timestamp 1701859473
transform 1 0 1430 0 1 10150
box -12 -8 32 272
use FILL  FILL_1__2718_
timestamp 1701859473
transform -1 0 10010 0 1 4950
box -12 -8 32 272
use FILL  FILL_1__2719_
timestamp 1701859473
transform -1 0 9770 0 1 4950
box -12 -8 32 272
use FILL  FILL_1__2720_
timestamp 1701859473
transform -1 0 4550 0 1 4950
box -12 -8 32 272
use FILL  FILL_1__2721_
timestamp 1701859473
transform -1 0 7310 0 -1 2350
box -12 -8 32 272
use FILL  FILL_1__2722_
timestamp 1701859473
transform 1 0 9950 0 -1 790
box -12 -8 32 272
use FILL  FILL_1__2723_
timestamp 1701859473
transform -1 0 7070 0 1 1830
box -12 -8 32 272
use FILL  FILL_1__2724_
timestamp 1701859473
transform -1 0 7070 0 -1 2350
box -12 -8 32 272
use FILL  FILL_1__2725_
timestamp 1701859473
transform 1 0 6930 0 1 3390
box -12 -8 32 272
use FILL  FILL_1__2726_
timestamp 1701859473
transform -1 0 7170 0 1 3390
box -12 -8 32 272
use FILL  FILL_1__2727_
timestamp 1701859473
transform -1 0 5390 0 1 3390
box -12 -8 32 272
use FILL  FILL_1__2728_
timestamp 1701859473
transform -1 0 5610 0 1 3390
box -12 -8 32 272
use FILL  FILL_1__2729_
timestamp 1701859473
transform -1 0 6710 0 -1 3910
box -12 -8 32 272
use FILL  FILL_1__2730_
timestamp 1701859473
transform 1 0 8210 0 -1 3910
box -12 -8 32 272
use FILL  FILL_1__2731_
timestamp 1701859473
transform 1 0 9230 0 1 1830
box -12 -8 32 272
use FILL  FILL_1__2732_
timestamp 1701859473
transform 1 0 7670 0 1 1830
box -12 -8 32 272
use FILL  FILL_1__2733_
timestamp 1701859473
transform 1 0 8550 0 1 2350
box -12 -8 32 272
use FILL  FILL_1__2734_
timestamp 1701859473
transform 1 0 7130 0 -1 5470
box -12 -8 32 272
use FILL  FILL_1__2735_
timestamp 1701859473
transform 1 0 7210 0 -1 2870
box -12 -8 32 272
use FILL  FILL_1__2736_
timestamp 1701859473
transform -1 0 7490 0 1 1310
box -12 -8 32 272
use FILL  FILL_1__2737_
timestamp 1701859473
transform 1 0 8550 0 1 1830
box -12 -8 32 272
use FILL  FILL_1__2738_
timestamp 1701859473
transform -1 0 7930 0 -1 2870
box -12 -8 32 272
use FILL  FILL_1__2739_
timestamp 1701859473
transform -1 0 7750 0 1 2870
box -12 -8 32 272
use FILL  FILL_1__2740_
timestamp 1701859473
transform -1 0 6530 0 -1 1830
box -12 -8 32 272
use FILL  FILL_1__2741_
timestamp 1701859473
transform 1 0 6730 0 -1 1830
box -12 -8 32 272
use FILL  FILL_1__2742_
timestamp 1701859473
transform -1 0 8170 0 -1 2870
box -12 -8 32 272
use FILL  FILL_1__2743_
timestamp 1701859473
transform -1 0 8190 0 1 2870
box -12 -8 32 272
use FILL  FILL_1__2744_
timestamp 1701859473
transform -1 0 7310 0 -1 270
box -12 -8 32 272
use FILL  FILL_1__2745_
timestamp 1701859473
transform -1 0 7270 0 1 1830
box -12 -8 32 272
use FILL  FILL_1__2746_
timestamp 1701859473
transform 1 0 7930 0 1 2870
box -12 -8 32 272
use FILL  FILL_1__2747_
timestamp 1701859473
transform -1 0 7730 0 -1 2350
box -12 -8 32 272
use FILL  FILL_1__2748_
timestamp 1701859473
transform 1 0 7910 0 -1 2350
box -12 -8 32 272
use FILL  FILL_1__2749_
timestamp 1701859473
transform 1 0 5870 0 1 1830
box -12 -8 32 272
use FILL  FILL_1__2750_
timestamp 1701859473
transform -1 0 6630 0 -1 1310
box -12 -8 32 272
use FILL  FILL_1__2751_
timestamp 1701859473
transform -1 0 6350 0 1 1830
box -12 -8 32 272
use FILL  FILL_1__2752_
timestamp 1701859473
transform -1 0 7710 0 1 2350
box -12 -8 32 272
use FILL  FILL_1__2753_
timestamp 1701859473
transform -1 0 7450 0 1 2350
box -12 -8 32 272
use FILL  FILL_1__2754_
timestamp 1701859473
transform 1 0 8790 0 -1 4950
box -12 -8 32 272
use FILL  FILL_1__2755_
timestamp 1701859473
transform 1 0 9690 0 1 790
box -12 -8 32 272
use FILL  FILL_1__2756_
timestamp 1701859473
transform -1 0 9930 0 1 790
box -12 -8 32 272
use FILL  FILL_1__2757_
timestamp 1701859473
transform 1 0 10630 0 -1 2870
box -12 -8 32 272
use FILL  FILL_1__2758_
timestamp 1701859473
transform -1 0 9130 0 -1 2870
box -12 -8 32 272
use FILL  FILL_1__2759_
timestamp 1701859473
transform 1 0 9050 0 1 4430
box -12 -8 32 272
use FILL  FILL_1__2760_
timestamp 1701859473
transform 1 0 10390 0 -1 790
box -12 -8 32 272
use FILL  FILL_1__2761_
timestamp 1701859473
transform 1 0 10150 0 -1 790
box -12 -8 32 272
use FILL  FILL_1__2762_
timestamp 1701859473
transform -1 0 10830 0 -1 1830
box -12 -8 32 272
use FILL  FILL_1__2763_
timestamp 1701859473
transform 1 0 6570 0 1 1830
box -12 -8 32 272
use FILL  FILL_1__2764_
timestamp 1701859473
transform -1 0 6830 0 1 1830
box -12 -8 32 272
use FILL  FILL_1__2765_
timestamp 1701859473
transform -1 0 10130 0 1 1830
box -12 -8 32 272
use FILL  FILL_1__2766_
timestamp 1701859473
transform -1 0 9950 0 -1 1830
box -12 -8 32 272
use FILL  FILL_1__2767_
timestamp 1701859473
transform -1 0 10370 0 -1 1830
box -12 -8 32 272
use FILL  FILL_1__2768_
timestamp 1701859473
transform -1 0 10350 0 1 1830
box -12 -8 32 272
use FILL  FILL_1__2769_
timestamp 1701859473
transform -1 0 10810 0 1 2350
box -12 -8 32 272
use FILL  FILL_1__2770_
timestamp 1701859473
transform -1 0 10590 0 -1 1830
box -12 -8 32 272
use FILL  FILL_1__2771_
timestamp 1701859473
transform 1 0 11010 0 1 2350
box -12 -8 32 272
use FILL  FILL_1__2772_
timestamp 1701859473
transform -1 0 10670 0 1 4950
box -12 -8 32 272
use FILL  FILL_1__2773_
timestamp 1701859473
transform 1 0 10410 0 -1 3910
box -12 -8 32 272
use FILL  FILL_1__2774_
timestamp 1701859473
transform -1 0 10710 0 -1 2350
box -12 -8 32 272
use FILL  FILL_1__2775_
timestamp 1701859473
transform -1 0 9070 0 -1 1310
box -12 -8 32 272
use FILL  FILL_1__2776_
timestamp 1701859473
transform 1 0 10610 0 -1 790
box -12 -8 32 272
use FILL  FILL_1__2777_
timestamp 1701859473
transform -1 0 8370 0 -1 270
box -12 -8 32 272
use FILL  FILL_1__2778_
timestamp 1701859473
transform 1 0 10910 0 1 270
box -12 -8 32 272
use FILL  FILL_1__2779_
timestamp 1701859473
transform 1 0 8990 0 -1 1830
box -12 -8 32 272
use FILL  FILL_1__2780_
timestamp 1701859473
transform -1 0 10010 0 1 1310
box -12 -8 32 272
use FILL  FILL_1__2781_
timestamp 1701859473
transform 1 0 10150 0 -1 1310
box -12 -8 32 272
use FILL  FILL_1__2782_
timestamp 1701859473
transform 1 0 8770 0 1 1830
box -12 -8 32 272
use FILL  FILL_1__2783_
timestamp 1701859473
transform 1 0 8330 0 -1 1310
box -12 -8 32 272
use FILL  FILL_1__2784_
timestamp 1701859473
transform 1 0 8570 0 -1 1310
box -12 -8 32 272
use FILL  FILL_1__2785_
timestamp 1701859473
transform 1 0 8790 0 -1 1830
box -12 -8 32 272
use FILL  FILL_1__2786_
timestamp 1701859473
transform -1 0 9270 0 -1 1310
box -12 -8 32 272
use FILL  FILL_1__2787_
timestamp 1701859473
transform -1 0 9470 0 -1 1830
box -12 -8 32 272
use FILL  FILL_1__2788_
timestamp 1701859473
transform 1 0 10150 0 -1 1830
box -12 -8 32 272
use FILL  FILL_1__2789_
timestamp 1701859473
transform 1 0 10230 0 1 1310
box -12 -8 32 272
use FILL  FILL_1__2790_
timestamp 1701859473
transform -1 0 10030 0 -1 2350
box -12 -8 32 272
use FILL  FILL_1__2791_
timestamp 1701859473
transform 1 0 9790 0 -1 2350
box -12 -8 32 272
use FILL  FILL_1__2792_
timestamp 1701859473
transform -1 0 10250 0 -1 2350
box -12 -8 32 272
use FILL  FILL_1__2793_
timestamp 1701859473
transform -1 0 10490 0 -1 2350
box -12 -8 32 272
use FILL  FILL_1__2794_
timestamp 1701859473
transform -1 0 10910 0 -1 2350
box -12 -8 32 272
use FILL  FILL_1__2795_
timestamp 1701859473
transform -1 0 10870 0 -1 2870
box -12 -8 32 272
use FILL  FILL_1__2796_
timestamp 1701859473
transform -1 0 10210 0 -1 2870
box -12 -8 32 272
use FILL  FILL_1__2797_
timestamp 1701859473
transform -1 0 9710 0 -1 1830
box -12 -8 32 272
use FILL  FILL_1__2798_
timestamp 1701859473
transform -1 0 10590 0 1 2350
box -12 -8 32 272
use FILL  FILL_1__2799_
timestamp 1701859473
transform 1 0 10370 0 -1 2870
box -12 -8 32 272
use FILL  FILL_1__2800_
timestamp 1701859473
transform -1 0 10390 0 -1 4430
box -12 -8 32 272
use FILL  FILL_1__2801_
timestamp 1701859473
transform -1 0 9350 0 -1 2870
box -12 -8 32 272
use FILL  FILL_1__2802_
timestamp 1701859473
transform -1 0 7210 0 -1 1830
box -12 -8 32 272
use FILL  FILL_1__2803_
timestamp 1701859473
transform 1 0 8410 0 -1 2870
box -12 -8 32 272
use FILL  FILL_1__2804_
timestamp 1701859473
transform -1 0 9470 0 -1 3390
box -12 -8 32 272
use FILL  FILL_1__2805_
timestamp 1701859473
transform -1 0 9770 0 -1 2870
box -12 -8 32 272
use FILL  FILL_1__2806_
timestamp 1701859473
transform 1 0 9530 0 -1 2870
box -12 -8 32 272
use FILL  FILL_1__2807_
timestamp 1701859473
transform 1 0 8870 0 -1 2350
box -12 -8 32 272
use FILL  FILL_1__2808_
timestamp 1701859473
transform 1 0 8630 0 -1 2350
box -12 -8 32 272
use FILL  FILL_1__2809_
timestamp 1701859473
transform 1 0 10350 0 1 2350
box -12 -8 32 272
use FILL  FILL_1__2810_
timestamp 1701859473
transform -1 0 10130 0 1 2350
box -12 -8 32 272
use FILL  FILL_1__2811_
timestamp 1701859473
transform 1 0 4910 0 -1 4430
box -12 -8 32 272
use FILL  FILL_1__2812_
timestamp 1701859473
transform -1 0 8870 0 1 4950
box -12 -8 32 272
use FILL  FILL_1__2813_
timestamp 1701859473
transform 1 0 8970 0 1 3390
box -12 -8 32 272
use FILL  FILL_1__2814_
timestamp 1701859473
transform -1 0 8790 0 -1 4430
box -12 -8 32 272
use FILL  FILL_1__2815_
timestamp 1701859473
transform -1 0 8570 0 1 3910
box -12 -8 32 272
use FILL  FILL_1__2816_
timestamp 1701859473
transform -1 0 8190 0 1 4950
box -12 -8 32 272
use FILL  FILL_1__2817_
timestamp 1701859473
transform 1 0 8630 0 1 4950
box -12 -8 32 272
use FILL  FILL_1__2818_
timestamp 1701859473
transform 1 0 8330 0 -1 4430
box -12 -8 32 272
use FILL  FILL_1__2819_
timestamp 1701859473
transform 1 0 8530 0 -1 4430
box -12 -8 32 272
use FILL  FILL_1__2820_
timestamp 1701859473
transform -1 0 9490 0 1 2350
box -12 -8 32 272
use FILL  FILL_1__2821_
timestamp 1701859473
transform 1 0 9010 0 1 2350
box -12 -8 32 272
use FILL  FILL_1__2822_
timestamp 1701859473
transform -1 0 9010 0 1 1830
box -12 -8 32 272
use FILL  FILL_1__2823_
timestamp 1701859473
transform -1 0 8790 0 1 2350
box -12 -8 32 272
use FILL  FILL_1__2824_
timestamp 1701859473
transform 1 0 9910 0 -1 3390
box -12 -8 32 272
use FILL  FILL_1__2825_
timestamp 1701859473
transform -1 0 10630 0 -1 3390
box -12 -8 32 272
use FILL  FILL_1__2826_
timestamp 1701859473
transform 1 0 9490 0 1 790
box -12 -8 32 272
use FILL  FILL_1__2827_
timestamp 1701859473
transform -1 0 9230 0 -1 1830
box -12 -8 32 272
use FILL  FILL_1__2828_
timestamp 1701859473
transform 1 0 6950 0 -1 1830
box -12 -8 32 272
use FILL  FILL_1__2829_
timestamp 1701859473
transform -1 0 9970 0 1 2870
box -12 -8 32 272
use FILL  FILL_1__2830_
timestamp 1701859473
transform 1 0 8270 0 -1 3390
box -12 -8 32 272
use FILL  FILL_1__2831_
timestamp 1701859473
transform 1 0 8310 0 1 3910
box -12 -8 32 272
use FILL  FILL_1__2832_
timestamp 1701859473
transform -1 0 9290 0 1 2350
box -12 -8 32 272
use FILL  FILL_1__2833_
timestamp 1701859473
transform -1 0 9230 0 -1 3390
box -12 -8 32 272
use FILL  FILL_1__2834_
timestamp 1701859473
transform -1 0 8990 0 -1 3390
box -12 -8 32 272
use FILL  FILL_1__2835_
timestamp 1701859473
transform -1 0 9290 0 1 790
box -12 -8 32 272
use FILL  FILL_1__2836_
timestamp 1701859473
transform 1 0 8870 0 1 1310
box -12 -8 32 272
use FILL  FILL_1__2837_
timestamp 1701859473
transform -1 0 9550 0 1 1310
box -12 -8 32 272
use FILL  FILL_1__2838_
timestamp 1701859473
transform -1 0 9670 0 1 3390
box -12 -8 32 272
use FILL  FILL_1__2839_
timestamp 1701859473
transform -1 0 9710 0 -1 3390
box -12 -8 32 272
use FILL  FILL_1__2840_
timestamp 1701859473
transform 1 0 9030 0 -1 270
box -12 -8 32 272
use FILL  FILL_1__2841_
timestamp 1701859473
transform -1 0 8830 0 -1 270
box -12 -8 32 272
use FILL  FILL_1__2842_
timestamp 1701859473
transform 1 0 9250 0 -1 270
box -12 -8 32 272
use FILL  FILL_1__2843_
timestamp 1701859473
transform 1 0 9490 0 -1 270
box -12 -8 32 272
use FILL  FILL_1__2844_
timestamp 1701859473
transform 1 0 9290 0 1 270
box -12 -8 32 272
use FILL  FILL_1__2845_
timestamp 1701859473
transform -1 0 9970 0 1 270
box -12 -8 32 272
use FILL  FILL_1__2846_
timestamp 1701859473
transform 1 0 9710 0 1 270
box -12 -8 32 272
use FILL  FILL_1__2847_
timestamp 1701859473
transform -1 0 11110 0 -1 10670
box -12 -8 32 272
use FILL  FILL_1__2848_
timestamp 1701859473
transform -1 0 10590 0 -1 1310
box -12 -8 32 272
use FILL  FILL_1__2849_
timestamp 1701859473
transform -1 0 10930 0 1 1310
box -12 -8 32 272
use FILL  FILL_1__2850_
timestamp 1701859473
transform -1 0 11070 0 -1 1830
box -12 -8 32 272
use FILL  FILL_1__2851_
timestamp 1701859473
transform 1 0 10670 0 -1 3910
box -12 -8 32 272
use FILL  FILL_1__2852_
timestamp 1701859473
transform -1 0 8870 0 1 270
box -12 -8 32 272
use FILL  FILL_1__2853_
timestamp 1701859473
transform -1 0 9090 0 1 270
box -12 -8 32 272
use FILL  FILL_1__2854_
timestamp 1701859473
transform 1 0 10590 0 1 790
box -12 -8 32 272
use FILL  FILL_1__2855_
timestamp 1701859473
transform -1 0 9790 0 1 1310
box -12 -8 32 272
use FILL  FILL_1__2856_
timestamp 1701859473
transform -1 0 10450 0 1 1310
box -12 -8 32 272
use FILL  FILL_1__2857_
timestamp 1701859473
transform -1 0 10690 0 1 1310
box -12 -8 32 272
use FILL  FILL_1__2858_
timestamp 1701859473
transform -1 0 11050 0 1 1830
box -12 -8 32 272
use FILL  FILL_1__2859_
timestamp 1701859473
transform 1 0 10910 0 -1 3910
box -12 -8 32 272
use FILL  FILL_1__2860_
timestamp 1701859473
transform 1 0 10830 0 -1 3390
box -12 -8 32 272
use FILL  FILL_1__2861_
timestamp 1701859473
transform 1 0 9710 0 -1 270
box -12 -8 32 272
use FILL  FILL_1__2862_
timestamp 1701859473
transform 1 0 8570 0 -1 270
box -12 -8 32 272
use FILL  FILL_1__2863_
timestamp 1701859473
transform -1 0 10210 0 1 270
box -12 -8 32 272
use FILL  FILL_1__2864_
timestamp 1701859473
transform 1 0 10450 0 1 270
box -12 -8 32 272
use FILL  FILL_1__2865_
timestamp 1701859473
transform -1 0 10690 0 1 270
box -12 -8 32 272
use FILL  FILL_1__2866_
timestamp 1701859473
transform -1 0 11070 0 -1 790
box -12 -8 32 272
use FILL  FILL_1__2867_
timestamp 1701859473
transform 1 0 11030 0 -1 3390
box -12 -8 32 272
use FILL  FILL_1__2868_
timestamp 1701859473
transform 1 0 11010 0 1 790
box -12 -8 32 272
use FILL  FILL_1__2869_
timestamp 1701859473
transform 1 0 10130 0 1 790
box -12 -8 32 272
use FILL  FILL_1__2870_
timestamp 1701859473
transform -1 0 10350 0 1 790
box -12 -8 32 272
use FILL  FILL_1__2871_
timestamp 1701859473
transform -1 0 10790 0 1 790
box -12 -8 32 272
use FILL  FILL_1__2872_
timestamp 1701859473
transform -1 0 11130 0 1 1310
box -12 -8 32 272
use FILL  FILL_1__2873_
timestamp 1701859473
transform -1 0 9910 0 1 3390
box -12 -8 32 272
use FILL  FILL_1__2874_
timestamp 1701859473
transform -1 0 10150 0 1 3390
box -12 -8 32 272
use FILL  FILL_1__2875_
timestamp 1701859473
transform -1 0 10730 0 -1 4950
box -12 -8 32 272
use FILL  FILL_1__2876_
timestamp 1701859473
transform -1 0 9690 0 1 1830
box -12 -8 32 272
use FILL  FILL_1__2877_
timestamp 1701859473
transform 1 0 9870 0 1 1830
box -12 -8 32 272
use FILL  FILL_1__2878_
timestamp 1701859473
transform 1 0 9690 0 -1 1310
box -12 -8 32 272
use FILL  FILL_1__2879_
timestamp 1701859473
transform -1 0 9930 0 -1 1310
box -12 -8 32 272
use FILL  FILL_1__2880_
timestamp 1701859473
transform 1 0 9430 0 1 1830
box -12 -8 32 272
use FILL  FILL_1__2881_
timestamp 1701859473
transform 1 0 10810 0 -1 790
box -12 -8 32 272
use FILL  FILL_1__2882_
timestamp 1701859473
transform -1 0 9490 0 -1 1310
box -12 -8 32 272
use FILL  FILL_1__2883_
timestamp 1701859473
transform -1 0 10390 0 -1 1310
box -12 -8 32 272
use FILL  FILL_1__2884_
timestamp 1701859473
transform 1 0 11030 0 -1 1310
box -12 -8 32 272
use FILL  FILL_1__2885_
timestamp 1701859473
transform -1 0 10810 0 -1 1310
box -12 -8 32 272
use FILL  FILL_1__2886_
timestamp 1701859473
transform 1 0 10570 0 1 1830
box -12 -8 32 272
use FILL  FILL_1__2887_
timestamp 1701859473
transform 1 0 10130 0 -1 4430
box -12 -8 32 272
use FILL  FILL_1__2888_
timestamp 1701859473
transform -1 0 3950 0 1 5470
box -12 -8 32 272
use FILL  FILL_1__2889_
timestamp 1701859473
transform 1 0 6070 0 1 2350
box -12 -8 32 272
use FILL  FILL_1__2890_
timestamp 1701859473
transform -1 0 8350 0 1 5990
box -12 -8 32 272
use FILL  FILL_1__2891_
timestamp 1701859473
transform -1 0 8150 0 1 5990
box -12 -8 32 272
use FILL  FILL_1__2892_
timestamp 1701859473
transform 1 0 7370 0 -1 5470
box -12 -8 32 272
use FILL  FILL_1__2893_
timestamp 1701859473
transform 1 0 7190 0 1 5470
box -12 -8 32 272
use FILL  FILL_1__2894_
timestamp 1701859473
transform 1 0 6470 0 -1 6510
box -12 -8 32 272
use FILL  FILL_1__2895_
timestamp 1701859473
transform 1 0 6610 0 1 6510
box -12 -8 32 272
use FILL  FILL_1__2896_
timestamp 1701859473
transform -1 0 7870 0 -1 5470
box -12 -8 32 272
use FILL  FILL_1__2897_
timestamp 1701859473
transform 1 0 7670 0 1 5470
box -12 -8 32 272
use FILL  FILL_1__2898_
timestamp 1701859473
transform 1 0 7190 0 -1 6510
box -12 -8 32 272
use FILL  FILL_1__2899_
timestamp 1701859473
transform 1 0 6710 0 -1 6510
box -12 -8 32 272
use FILL  FILL_1__2900_
timestamp 1701859473
transform -1 0 6250 0 -1 6510
box -12 -8 32 272
use FILL  FILL_1__2901_
timestamp 1701859473
transform 1 0 5990 0 -1 6510
box -12 -8 32 272
use FILL  FILL_1__2902_
timestamp 1701859473
transform -1 0 7910 0 1 5990
box -12 -8 32 272
use FILL  FILL_1__2903_
timestamp 1701859473
transform 1 0 7190 0 1 5990
box -12 -8 32 272
use FILL  FILL_1__2904_
timestamp 1701859473
transform 1 0 8310 0 -1 5470
box -12 -8 32 272
use FILL  FILL_1__2905_
timestamp 1701859473
transform 1 0 8330 0 1 5470
box -12 -8 32 272
use FILL  FILL_1__2906_
timestamp 1701859473
transform 1 0 8070 0 -1 5990
box -12 -8 32 272
use FILL  FILL_1__2907_
timestamp 1701859473
transform -1 0 7850 0 -1 5990
box -12 -8 32 272
use FILL  FILL_1__2908_
timestamp 1701859473
transform -1 0 8170 0 -1 4950
box -12 -8 32 272
use FILL  FILL_1__2909_
timestamp 1701859473
transform 1 0 3310 0 -1 4430
box -12 -8 32 272
use FILL  FILL_1__2910_
timestamp 1701859473
transform -1 0 6470 0 -1 4430
box -12 -8 32 272
use FILL  FILL_1__2911_
timestamp 1701859473
transform -1 0 6810 0 1 4430
box -12 -8 32 272
use FILL  FILL_1__2912_
timestamp 1701859473
transform 1 0 8590 0 -1 4950
box -12 -8 32 272
use FILL  FILL_1__2913_
timestamp 1701859473
transform -1 0 6770 0 -1 4950
box -12 -8 32 272
use FILL  FILL_1__2914_
timestamp 1701859473
transform 1 0 7030 0 -1 8070
box -12 -8 32 272
use FILL  FILL_1__2915_
timestamp 1701859473
transform 1 0 7150 0 -1 5990
box -12 -8 32 272
use FILL  FILL_1__2916_
timestamp 1701859473
transform 1 0 6910 0 -1 5990
box -12 -8 32 272
use FILL  FILL_1__2917_
timestamp 1701859473
transform -1 0 6290 0 -1 5990
box -12 -8 32 272
use FILL  FILL_1__2918_
timestamp 1701859473
transform 1 0 6210 0 1 5470
box -12 -8 32 272
use FILL  FILL_1__2919_
timestamp 1701859473
transform 1 0 6130 0 1 4950
box -12 -8 32 272
use FILL  FILL_1__2920_
timestamp 1701859473
transform 1 0 5890 0 1 4950
box -12 -8 32 272
use FILL  FILL_1__2921_
timestamp 1701859473
transform -1 0 7350 0 -1 3910
box -12 -8 32 272
use FILL  FILL_1__2922_
timestamp 1701859473
transform -1 0 7390 0 1 3910
box -12 -8 32 272
use FILL  FILL_1__2923_
timestamp 1701859473
transform -1 0 6710 0 -1 4430
box -12 -8 32 272
use FILL  FILL_1__2924_
timestamp 1701859473
transform 1 0 6330 0 1 4950
box -12 -8 32 272
use FILL  FILL_1__2925_
timestamp 1701859473
transform 1 0 7230 0 1 7550
box -12 -8 32 272
use FILL  FILL_1__2926_
timestamp 1701859473
transform -1 0 7470 0 1 4430
box -12 -8 32 272
use FILL  FILL_1__2927_
timestamp 1701859473
transform 1 0 7250 0 -1 4950
box -12 -8 32 272
use FILL  FILL_1__2928_
timestamp 1701859473
transform 1 0 6990 0 -1 4950
box -12 -8 32 272
use FILL  FILL_1__2929_
timestamp 1701859473
transform -1 0 6570 0 1 4950
box -12 -8 32 272
use FILL  FILL_1__2930_
timestamp 1701859473
transform 1 0 6110 0 1 1830
box -12 -8 32 272
use FILL  FILL_1__2931_
timestamp 1701859473
transform 1 0 6990 0 -1 2870
box -12 -8 32 272
use FILL  FILL_1__2932_
timestamp 1701859473
transform 1 0 5150 0 -1 4430
box -12 -8 32 272
use FILL  FILL_1__2933_
timestamp 1701859473
transform 1 0 5350 0 -1 4430
box -12 -8 32 272
use FILL  FILL_1__2934_
timestamp 1701859473
transform 1 0 5590 0 -1 4430
box -12 -8 32 272
use FILL  FILL_1__2935_
timestamp 1701859473
transform 1 0 6410 0 1 6510
box -12 -8 32 272
use FILL  FILL_1__2936_
timestamp 1701859473
transform 1 0 6290 0 -1 4950
box -12 -8 32 272
use FILL  FILL_1__2937_
timestamp 1701859473
transform 1 0 6510 0 -1 4950
box -12 -8 32 272
use FILL  FILL_1__2938_
timestamp 1701859473
transform 1 0 4990 0 1 4950
box -12 -8 32 272
use FILL  FILL_1__2939_
timestamp 1701859473
transform 1 0 4770 0 1 4950
box -12 -8 32 272
use FILL  FILL_1__2940_
timestamp 1701859473
transform -1 0 5830 0 -1 5470
box -12 -8 32 272
use FILL  FILL_1__2941_
timestamp 1701859473
transform 1 0 5590 0 -1 5470
box -12 -8 32 272
use FILL  FILL_1__2942_
timestamp 1701859473
transform -1 0 9290 0 1 4430
box -12 -8 32 272
use FILL  FILL_1__2943_
timestamp 1701859473
transform 1 0 6250 0 -1 4430
box -12 -8 32 272
use FILL  FILL_1__2944_
timestamp 1701859473
transform -1 0 6270 0 1 3910
box -12 -8 32 272
use FILL  FILL_1__2945_
timestamp 1701859473
transform -1 0 6350 0 1 4430
box -12 -8 32 272
use FILL  FILL_1__2946_
timestamp 1701859473
transform 1 0 6110 0 1 4430
box -12 -8 32 272
use FILL  FILL_1__2947_
timestamp 1701859473
transform -1 0 6510 0 -1 5990
box -12 -8 32 272
use FILL  FILL_1__2948_
timestamp 1701859473
transform 1 0 6050 0 -1 5990
box -12 -8 32 272
use FILL  FILL_1__2949_
timestamp 1701859473
transform -1 0 5870 0 -1 5990
box -12 -8 32 272
use FILL  FILL_1__2950_
timestamp 1701859473
transform 1 0 5730 0 1 5470
box -12 -8 32 272
use FILL  FILL_1__2951_
timestamp 1701859473
transform -1 0 5990 0 1 5470
box -12 -8 32 272
use FILL  FILL_1__2952_
timestamp 1701859473
transform -1 0 6070 0 -1 4950
box -12 -8 32 272
use FILL  FILL_1__2953_
timestamp 1701859473
transform -1 0 4350 0 1 4950
box -12 -8 32 272
use FILL  FILL_1__2954_
timestamp 1701859473
transform -1 0 6610 0 1 4430
box -12 -8 32 272
use FILL  FILL_1__2955_
timestamp 1701859473
transform -1 0 5890 0 1 4430
box -12 -8 32 272
use FILL  FILL_1__2956_
timestamp 1701859473
transform 1 0 5170 0 1 4430
box -12 -8 32 272
use FILL  FILL_1__2957_
timestamp 1701859473
transform 1 0 5110 0 -1 4950
box -12 -8 32 272
use FILL  FILL_1__2958_
timestamp 1701859473
transform -1 0 5430 0 1 4430
box -12 -8 32 272
use FILL  FILL_1__2959_
timestamp 1701859473
transform 1 0 6930 0 -1 5470
box -12 -8 32 272
use FILL  FILL_1__2960_
timestamp 1701859473
transform -1 0 6470 0 1 5470
box -12 -8 32 272
use FILL  FILL_1__2961_
timestamp 1701859473
transform 1 0 6230 0 -1 5470
box -12 -8 32 272
use FILL  FILL_1__2962_
timestamp 1701859473
transform -1 0 6490 0 -1 5470
box -12 -8 32 272
use FILL  FILL_1__2963_
timestamp 1701859473
transform -1 0 6730 0 -1 5470
box -12 -8 32 272
use FILL  FILL_1__2964_
timestamp 1701859473
transform -1 0 5370 0 -1 4950
box -12 -8 32 272
use FILL  FILL_1__2965_
timestamp 1701859473
transform 1 0 4870 0 -1 4950
box -12 -8 32 272
use FILL  FILL_1__2966_
timestamp 1701859473
transform -1 0 6330 0 1 2350
box -12 -8 32 272
use FILL  FILL_1__2967_
timestamp 1701859473
transform 1 0 7590 0 1 3910
box -12 -8 32 272
use FILL  FILL_1__2968_
timestamp 1701859473
transform -1 0 6910 0 -1 3910
box -12 -8 32 272
use FILL  FILL_1__2969_
timestamp 1701859473
transform -1 0 7130 0 -1 3910
box -12 -8 32 272
use FILL  FILL_1__2970_
timestamp 1701859473
transform -1 0 7170 0 1 3910
box -12 -8 32 272
use FILL  FILL_1__2971_
timestamp 1701859473
transform -1 0 6690 0 1 3910
box -12 -8 32 272
use FILL  FILL_1__2972_
timestamp 1701859473
transform 1 0 6910 0 1 3910
box -12 -8 32 272
use FILL  FILL_1__2973_
timestamp 1701859473
transform -1 0 7030 0 1 4430
box -12 -8 32 272
use FILL  FILL_1__2974_
timestamp 1701859473
transform 1 0 6930 0 -1 4430
box -12 -8 32 272
use FILL  FILL_1__2975_
timestamp 1701859473
transform -1 0 7690 0 -1 4430
box -12 -8 32 272
use FILL  FILL_1__2976_
timestamp 1701859473
transform -1 0 7450 0 -1 4430
box -12 -8 32 272
use FILL  FILL_1__2977_
timestamp 1701859473
transform 1 0 7170 0 -1 4430
box -12 -8 32 272
use FILL  FILL_1__2978_
timestamp 1701859473
transform 1 0 7230 0 1 4430
box -12 -8 32 272
use FILL  FILL_1__2979_
timestamp 1701859473
transform -1 0 3570 0 -1 4950
box -12 -8 32 272
use FILL  FILL_1__2980_
timestamp 1701859473
transform -1 0 2950 0 1 7550
box -12 -8 32 272
use FILL  FILL_1__2981_
timestamp 1701859473
transform 1 0 3470 0 1 4950
box -12 -8 32 272
use FILL  FILL_1__2982_
timestamp 1701859473
transform 1 0 9530 0 1 6510
box -12 -8 32 272
use FILL  FILL_1__2983_
timestamp 1701859473
transform 1 0 1850 0 1 4430
box -12 -8 32 272
use FILL  FILL_1__2984_
timestamp 1701859473
transform -1 0 3470 0 -1 3910
box -12 -8 32 272
use FILL  FILL_1__2985_
timestamp 1701859473
transform 1 0 3630 0 1 4430
box -12 -8 32 272
use FILL  FILL_1__2986_
timestamp 1701859473
transform -1 0 5830 0 -1 4430
box -12 -8 32 272
use FILL  FILL_1__2987_
timestamp 1701859473
transform -1 0 5650 0 1 4430
box -12 -8 32 272
use FILL  FILL_1__2988_
timestamp 1701859473
transform 1 0 9310 0 1 6510
box -12 -8 32 272
use FILL  FILL_1__2989_
timestamp 1701859473
transform 1 0 5930 0 1 6510
box -12 -8 32 272
use FILL  FILL_1__2990_
timestamp 1701859473
transform -1 0 6190 0 1 6510
box -12 -8 32 272
use FILL  FILL_1__2991_
timestamp 1701859473
transform 1 0 7090 0 1 6510
box -12 -8 32 272
use FILL  FILL_1__2992_
timestamp 1701859473
transform 1 0 9610 0 1 7030
box -12 -8 32 272
use FILL  FILL_1__2993_
timestamp 1701859473
transform 1 0 9810 0 1 7030
box -12 -8 32 272
use FILL  FILL_1__2994_
timestamp 1701859473
transform -1 0 10730 0 -1 7550
box -12 -8 32 272
use FILL  FILL_1__2995_
timestamp 1701859473
transform -1 0 7530 0 -1 7550
box -12 -8 32 272
use FILL  FILL_1__2996_
timestamp 1701859473
transform 1 0 7430 0 1 7550
box -12 -8 32 272
use FILL  FILL_1__2997_
timestamp 1701859473
transform -1 0 7310 0 -1 7550
box -12 -8 32 272
use FILL  FILL_1__2998_
timestamp 1701859473
transform -1 0 6370 0 -1 7550
box -12 -8 32 272
use FILL  FILL_1__2999_
timestamp 1701859473
transform 1 0 6090 0 1 7550
box -12 -8 32 272
use FILL  FILL_1__3000_
timestamp 1701859473
transform -1 0 5930 0 -1 7550
box -12 -8 32 272
use FILL  FILL_1__3001_
timestamp 1701859473
transform -1 0 5710 0 -1 7550
box -12 -8 32 272
use FILL  FILL_1__3002_
timestamp 1701859473
transform -1 0 6130 0 -1 7550
box -12 -8 32 272
use FILL  FILL_1__3003_
timestamp 1701859473
transform -1 0 6310 0 1 7550
box -12 -8 32 272
use FILL  FILL_1__3004_
timestamp 1701859473
transform 1 0 8110 0 1 7550
box -12 -8 32 272
use FILL  FILL_1__3005_
timestamp 1701859473
transform 1 0 10930 0 -1 7550
box -12 -8 32 272
use FILL  FILL_1__3006_
timestamp 1701859473
transform -1 0 10410 0 1 7550
box -12 -8 32 272
use FILL  FILL_1__3007_
timestamp 1701859473
transform 1 0 6930 0 1 7030
box -12 -8 32 272
use FILL  FILL_1__3008_
timestamp 1701859473
transform -1 0 6490 0 1 7030
box -12 -8 32 272
use FILL  FILL_1__3009_
timestamp 1701859473
transform -1 0 5890 0 -1 7030
box -12 -8 32 272
use FILL  FILL_1__3010_
timestamp 1701859473
transform 1 0 6110 0 -1 7030
box -12 -8 32 272
use FILL  FILL_1__3011_
timestamp 1701859473
transform 1 0 6690 0 1 7030
box -12 -8 32 272
use FILL  FILL_1__3012_
timestamp 1701859473
transform -1 0 7810 0 -1 7030
box -12 -8 32 272
use FILL  FILL_1__3013_
timestamp 1701859473
transform 1 0 8250 0 -1 7030
box -12 -8 32 272
use FILL  FILL_1__3014_
timestamp 1701859473
transform 1 0 10610 0 1 7550
box -12 -8 32 272
use FILL  FILL_1__3015_
timestamp 1701859473
transform -1 0 6330 0 -1 7030
box -12 -8 32 272
use FILL  FILL_1__3016_
timestamp 1701859473
transform -1 0 7210 0 1 7030
box -12 -8 32 272
use FILL  FILL_1__3017_
timestamp 1701859473
transform 1 0 6550 0 -1 7030
box -12 -8 32 272
use FILL  FILL_1__3018_
timestamp 1701859473
transform -1 0 6850 0 -1 7030
box -12 -8 32 272
use FILL  FILL_1__3019_
timestamp 1701859473
transform -1 0 7090 0 -1 7030
box -12 -8 32 272
use FILL  FILL_1__3020_
timestamp 1701859473
transform 1 0 8250 0 1 7030
box -12 -8 32 272
use FILL  FILL_1__3021_
timestamp 1701859473
transform -1 0 9310 0 -1 8070
box -12 -8 32 272
use FILL  FILL_1__3022_
timestamp 1701859473
transform 1 0 9490 0 -1 8070
box -12 -8 32 272
use FILL  FILL_1__3023_
timestamp 1701859473
transform -1 0 5710 0 1 6510
box -12 -8 32 272
use FILL  FILL_1__3024_
timestamp 1701859473
transform 1 0 5450 0 1 6510
box -12 -8 32 272
use FILL  FILL_1__3025_
timestamp 1701859473
transform -1 0 5470 0 -1 6510
box -12 -8 32 272
use FILL  FILL_1__3026_
timestamp 1701859473
transform 1 0 10890 0 -1 5990
box -12 -8 32 272
use FILL  FILL_1__3027_
timestamp 1701859473
transform -1 0 11130 0 -1 5990
box -12 -8 32 272
use FILL  FILL_1__3028_
timestamp 1701859473
transform -1 0 9750 0 -1 8070
box -12 -8 32 272
use FILL  FILL_1__3029_
timestamp 1701859473
transform -1 0 7070 0 -1 7550
box -12 -8 32 272
use FILL  FILL_1__3030_
timestamp 1701859473
transform -1 0 8050 0 -1 7030
box -12 -8 32 272
use FILL  FILL_1__3031_
timestamp 1701859473
transform 1 0 8030 0 1 7030
box -12 -8 32 272
use FILL  FILL_1__3032_
timestamp 1701859473
transform 1 0 7650 0 1 7550
box -12 -8 32 272
use FILL  FILL_1__3033_
timestamp 1701859473
transform -1 0 6730 0 1 8070
box -12 -8 32 272
use FILL  FILL_1__3034_
timestamp 1701859473
transform -1 0 7710 0 -1 8070
box -12 -8 32 272
use FILL  FILL_1__3035_
timestamp 1701859473
transform 1 0 7450 0 -1 8070
box -12 -8 32 272
use FILL  FILL_1__3036_
timestamp 1701859473
transform -1 0 6930 0 1 8070
box -12 -8 32 272
use FILL  FILL_1__3037_
timestamp 1701859473
transform -1 0 6490 0 1 8070
box -12 -8 32 272
use FILL  FILL_1__3038_
timestamp 1701859473
transform -1 0 7110 0 1 8070
box -12 -8 32 272
use FILL  FILL_1__3039_
timestamp 1701859473
transform 1 0 7330 0 1 8070
box -12 -8 32 272
use FILL  FILL_1__3040_
timestamp 1701859473
transform 1 0 9670 0 1 7550
box -12 -8 32 272
use FILL  FILL_1__3041_
timestamp 1701859473
transform -1 0 9530 0 -1 6510
box -12 -8 32 272
use FILL  FILL_1__3042_
timestamp 1701859473
transform 1 0 7230 0 -1 8070
box -12 -8 32 272
use FILL  FILL_1__3043_
timestamp 1701859473
transform -1 0 6550 0 1 7550
box -12 -8 32 272
use FILL  FILL_1__3044_
timestamp 1701859473
transform -1 0 6590 0 -1 7550
box -12 -8 32 272
use FILL  FILL_1__3045_
timestamp 1701859473
transform 1 0 6810 0 -1 7550
box -12 -8 32 272
use FILL  FILL_1__3046_
timestamp 1701859473
transform -1 0 7770 0 1 6510
box -12 -8 32 272
use FILL  FILL_1__3047_
timestamp 1701859473
transform 1 0 9110 0 1 6510
box -12 -8 32 272
use FILL  FILL_1__3048_
timestamp 1701859473
transform 1 0 9730 0 -1 6510
box -12 -8 32 272
use FILL  FILL_1__3049_
timestamp 1701859473
transform -1 0 6810 0 1 7550
box -12 -8 32 272
use FILL  FILL_1__3050_
timestamp 1701859473
transform -1 0 7030 0 1 7550
box -12 -8 32 272
use FILL  FILL_1__3051_
timestamp 1701859473
transform -1 0 7770 0 1 7030
box -12 -8 32 272
use FILL  FILL_1__3052_
timestamp 1701859473
transform 1 0 7470 0 1 7030
box -12 -8 32 272
use FILL  FILL_1__3053_
timestamp 1701859473
transform 1 0 7310 0 -1 7030
box -12 -8 32 272
use FILL  FILL_1__3054_
timestamp 1701859473
transform -1 0 7570 0 -1 7030
box -12 -8 32 272
use FILL  FILL_1__3055_
timestamp 1701859473
transform 1 0 7990 0 1 6510
box -12 -8 32 272
use FILL  FILL_1__3056_
timestamp 1701859473
transform -1 0 9510 0 1 5470
box -12 -8 32 272
use FILL  FILL_1__3057_
timestamp 1701859473
transform -1 0 9270 0 1 5470
box -12 -8 32 272
use FILL  FILL_1__3058_
timestamp 1701859473
transform 1 0 8690 0 -1 7550
box -12 -8 32 272
use FILL  FILL_1__3059_
timestamp 1701859473
transform -1 0 8570 0 -1 5990
box -12 -8 32 272
use FILL  FILL_1__3060_
timestamp 1701859473
transform 1 0 9750 0 1 6510
box -12 -8 32 272
use FILL  FILL_1__3061_
timestamp 1701859473
transform 1 0 9990 0 1 6510
box -12 -8 32 272
use FILL  FILL_1__3062_
timestamp 1701859473
transform -1 0 9610 0 -1 7550
box -12 -8 32 272
use FILL  FILL_1__3063_
timestamp 1701859473
transform 1 0 9350 0 -1 7550
box -12 -8 32 272
use FILL  FILL_1__3064_
timestamp 1701859473
transform -1 0 10310 0 -1 7030
box -12 -8 32 272
use FILL  FILL_1__3065_
timestamp 1701859473
transform -1 0 10550 0 -1 7030
box -12 -8 32 272
use FILL  FILL_1__3066_
timestamp 1701859473
transform -1 0 8470 0 -1 7550
box -12 -8 32 272
use FILL  FILL_1__3067_
timestamp 1701859473
transform 1 0 8210 0 -1 7550
box -12 -8 32 272
use FILL  FILL_1__3068_
timestamp 1701859473
transform 1 0 10170 0 -1 5990
box -12 -8 32 272
use FILL  FILL_1__3069_
timestamp 1701859473
transform 1 0 10410 0 -1 5990
box -12 -8 32 272
use FILL  FILL_1__3070_
timestamp 1701859473
transform 1 0 8870 0 -1 7550
box -12 -8 32 272
use FILL  FILL_1__3071_
timestamp 1701859473
transform -1 0 9130 0 -1 7550
box -12 -8 32 272
use FILL  FILL_1__3072_
timestamp 1701859473
transform -1 0 9750 0 1 5990
box -12 -8 32 272
use FILL  FILL_1__3073_
timestamp 1701859473
transform -1 0 9970 0 1 5990
box -12 -8 32 272
use FILL  FILL_1__3074_
timestamp 1701859473
transform 1 0 8790 0 1 5990
box -12 -8 32 272
use FILL  FILL_1__3075_
timestamp 1701859473
transform 1 0 8790 0 -1 5990
box -12 -8 32 272
use FILL  FILL_1__3076_
timestamp 1701859473
transform 1 0 10690 0 1 6510
box -12 -8 32 272
use FILL  FILL_1__3077_
timestamp 1701859473
transform 1 0 10890 0 1 6510
box -12 -8 32 272
use FILL  FILL_1__3078_
timestamp 1701859473
transform -1 0 8690 0 -1 7030
box -12 -8 32 272
use FILL  FILL_1__3079_
timestamp 1701859473
transform -1 0 8470 0 -1 7030
box -12 -8 32 272
use FILL  FILL_1__3080_
timestamp 1701859473
transform 1 0 10950 0 -1 8590
box -12 -8 32 272
use FILL  FILL_1__3081_
timestamp 1701859473
transform -1 0 10950 0 -1 270
box -12 -8 32 272
use FILL  FILL_1__3082_
timestamp 1701859473
transform 1 0 10050 0 -1 8590
box -12 -8 32 272
use FILL  FILL_1__3083_
timestamp 1701859473
transform -1 0 9830 0 -1 8590
box -12 -8 32 272
use FILL  FILL_1__3084_
timestamp 1701859473
transform -1 0 9010 0 1 7550
box -12 -8 32 272
use FILL  FILL_1__3085_
timestamp 1701859473
transform 1 0 8910 0 1 7030
box -12 -8 32 272
use FILL  FILL_1__3086_
timestamp 1701859473
transform -1 0 10670 0 1 5990
box -12 -8 32 272
use FILL  FILL_1__3087_
timestamp 1701859473
transform 1 0 10870 0 1 5990
box -12 -8 32 272
use FILL  FILL_1__3088_
timestamp 1701859473
transform 1 0 8230 0 1 8070
box -12 -8 32 272
use FILL  FILL_1__3089_
timestamp 1701859473
transform -1 0 8010 0 1 8070
box -12 -8 32 272
use FILL  FILL_1__3090_
timestamp 1701859473
transform -1 0 11110 0 1 4950
box -12 -8 32 272
use FILL  FILL_1__3091_
timestamp 1701859473
transform 1 0 10850 0 1 4950
box -12 -8 32 272
use FILL  FILL_1__3092_
timestamp 1701859473
transform 1 0 8770 0 -1 5470
box -12 -8 32 272
use FILL  FILL_1__3093_
timestamp 1701859473
transform -1 0 9010 0 -1 5470
box -12 -8 32 272
use FILL  FILL_1__3094_
timestamp 1701859473
transform -1 0 10210 0 -1 5470
box -12 -8 32 272
use FILL  FILL_1__3095_
timestamp 1701859473
transform 1 0 10150 0 1 5470
box -12 -8 32 272
use FILL  FILL_1__3096_
timestamp 1701859473
transform 1 0 8890 0 1 6510
box -12 -8 32 272
use FILL  FILL_1__3097_
timestamp 1701859473
transform -1 0 8670 0 1 6510
box -12 -8 32 272
use FILL  FILL_1__3098_
timestamp 1701859473
transform -1 0 10370 0 1 8070
box -12 -8 32 272
use FILL  FILL_1__3099_
timestamp 1701859473
transform -1 0 11130 0 -1 8070
box -12 -8 32 272
use FILL  FILL_1__3100_
timestamp 1701859473
transform 1 0 10130 0 1 8070
box -12 -8 32 272
use FILL  FILL_1__3101_
timestamp 1701859473
transform 1 0 10270 0 -1 8590
box -12 -8 32 272
use FILL  FILL_1__3102_
timestamp 1701859473
transform 1 0 8350 0 -1 8070
box -12 -8 32 272
use FILL  FILL_1__3103_
timestamp 1701859473
transform -1 0 8330 0 1 7550
box -12 -8 32 272
use FILL  FILL_1__3104_
timestamp 1701859473
transform -1 0 11130 0 1 6510
box -12 -8 32 272
use FILL  FILL_1__3105_
timestamp 1701859473
transform -1 0 10930 0 -1 4950
box -12 -8 32 272
use FILL  FILL_1__3106_
timestamp 1701859473
transform 1 0 9350 0 -1 8590
box -12 -8 32 272
use FILL  FILL_1__3107_
timestamp 1701859473
transform -1 0 9590 0 -1 8590
box -12 -8 32 272
use FILL  FILL_1__3108_
timestamp 1701859473
transform 1 0 9950 0 1 5470
box -12 -8 32 272
use FILL  FILL_1__3109_
timestamp 1701859473
transform -1 0 9730 0 1 5470
box -12 -8 32 272
use FILL  FILL_1__3110_
timestamp 1701859473
transform 1 0 8370 0 -1 6510
box -12 -8 32 272
use FILL  FILL_1__3111_
timestamp 1701859473
transform -1 0 8150 0 -1 6510
box -12 -8 32 272
use FILL  FILL_1__3112_
timestamp 1701859473
transform 1 0 490 0 -1 2870
box -12 -8 32 272
use FILL  FILL_1__3113_
timestamp 1701859473
transform 1 0 30 0 -1 2870
box -12 -8 32 272
use FILL  FILL_1__3114_
timestamp 1701859473
transform -1 0 290 0 -1 2870
box -12 -8 32 272
use FILL  FILL_1__3115_
timestamp 1701859473
transform -1 0 1170 0 1 2350
box -12 -8 32 272
use FILL  FILL_1__3116_
timestamp 1701859473
transform 1 0 930 0 -1 2350
box -12 -8 32 272
use FILL  FILL_1__3117_
timestamp 1701859473
transform 1 0 2010 0 -1 1310
box -12 -8 32 272
use FILL  FILL_1__3118_
timestamp 1701859473
transform -1 0 1390 0 -1 2350
box -12 -8 32 272
use FILL  FILL_1__3119_
timestamp 1701859473
transform -1 0 1150 0 -1 2350
box -12 -8 32 272
use FILL  FILL_1__3120_
timestamp 1701859473
transform -1 0 450 0 1 2350
box -12 -8 32 272
use FILL  FILL_1__3121_
timestamp 1701859473
transform 1 0 230 0 1 2870
box -12 -8 32 272
use FILL  FILL_1__3122_
timestamp 1701859473
transform 1 0 2490 0 -1 3390
box -12 -8 32 272
use FILL  FILL_1__3123_
timestamp 1701859473
transform 1 0 510 0 1 3390
box -12 -8 32 272
use FILL  FILL_1__3124_
timestamp 1701859473
transform -1 0 290 0 1 3390
box -12 -8 32 272
use FILL  FILL_1__3125_
timestamp 1701859473
transform -1 0 710 0 -1 2350
box -12 -8 32 272
use FILL  FILL_1__3126_
timestamp 1701859473
transform -1 0 1410 0 1 2350
box -12 -8 32 272
use FILL  FILL_1__3127_
timestamp 1701859473
transform -1 0 930 0 1 2350
box -12 -8 32 272
use FILL  FILL_1__3128_
timestamp 1701859473
transform -1 0 1870 0 1 2350
box -12 -8 32 272
use FILL  FILL_1__3129_
timestamp 1701859473
transform -1 0 1630 0 -1 2350
box -12 -8 32 272
use FILL  FILL_1__3130_
timestamp 1701859473
transform -1 0 1650 0 1 2350
box -12 -8 32 272
use FILL  FILL_1__3131_
timestamp 1701859473
transform -1 0 690 0 1 2350
box -12 -8 32 272
use FILL  FILL_1__3132_
timestamp 1701859473
transform 1 0 450 0 1 2870
box -12 -8 32 272
use FILL  FILL_1__3133_
timestamp 1701859473
transform 1 0 510 0 -1 3910
box -12 -8 32 272
use FILL  FILL_1__3134_
timestamp 1701859473
transform -1 0 1190 0 1 3390
box -12 -8 32 272
use FILL  FILL_1__3135_
timestamp 1701859473
transform 1 0 950 0 1 3390
box -12 -8 32 272
use FILL  FILL_1__3136_
timestamp 1701859473
transform -1 0 530 0 -1 3390
box -12 -8 32 272
use FILL  FILL_1__3137_
timestamp 1701859473
transform 1 0 250 0 -1 3390
box -12 -8 32 272
use FILL  FILL_1__3138_
timestamp 1701859473
transform -1 0 1650 0 1 4430
box -12 -8 32 272
use FILL  FILL_1__3139_
timestamp 1701859473
transform -1 0 1850 0 -1 3390
box -12 -8 32 272
use FILL  FILL_1__3140_
timestamp 1701859473
transform -1 0 270 0 1 3910
box -12 -8 32 272
use FILL  FILL_1__3141_
timestamp 1701859473
transform 1 0 710 0 1 4430
box -12 -8 32 272
use FILL  FILL_1__3142_
timestamp 1701859473
transform 1 0 950 0 1 4430
box -12 -8 32 272
use FILL  FILL_1__3143_
timestamp 1701859473
transform 1 0 970 0 -1 4430
box -12 -8 32 272
use FILL  FILL_1__3144_
timestamp 1701859473
transform -1 0 1210 0 -1 4430
box -12 -8 32 272
use FILL  FILL_1__3145_
timestamp 1701859473
transform -1 0 490 0 1 3910
box -12 -8 32 272
use FILL  FILL_1__3146_
timestamp 1701859473
transform -1 0 710 0 1 3910
box -12 -8 32 272
use FILL  FILL_1__3147_
timestamp 1701859473
transform 1 0 490 0 -1 4430
box -12 -8 32 272
use FILL  FILL_1__3148_
timestamp 1701859473
transform -1 0 750 0 -1 4430
box -12 -8 32 272
use FILL  FILL_1__3149_
timestamp 1701859473
transform -1 0 50 0 -1 3910
box -12 -8 32 272
use FILL  FILL_1__3150_
timestamp 1701859473
transform -1 0 910 0 1 3910
box -12 -8 32 272
use FILL  FILL_1__3151_
timestamp 1701859473
transform 1 0 30 0 1 3910
box -12 -8 32 272
use FILL  FILL_1__3152_
timestamp 1701859473
transform 1 0 30 0 -1 4430
box -12 -8 32 272
use FILL  FILL_1__3153_
timestamp 1701859473
transform -1 0 270 0 -1 4430
box -12 -8 32 272
use FILL  FILL_1__3154_
timestamp 1701859473
transform -1 0 770 0 -1 3390
box -12 -8 32 272
use FILL  FILL_1__3155_
timestamp 1701859473
transform -1 0 50 0 1 2870
box -12 -8 32 272
use FILL  FILL_1__3156_
timestamp 1701859473
transform 1 0 30 0 -1 3390
box -12 -8 32 272
use FILL  FILL_1__3157_
timestamp 1701859473
transform -1 0 50 0 1 3390
box -12 -8 32 272
use FILL  FILL_1__3158_
timestamp 1701859473
transform 1 0 30 0 1 4430
box -12 -8 32 272
use FILL  FILL_1__3159_
timestamp 1701859473
transform 1 0 250 0 1 4430
box -12 -8 32 272
use FILL  FILL_1__3160_
timestamp 1701859473
transform -1 0 490 0 1 4430
box -12 -8 32 272
use FILL  FILL_1__3161_
timestamp 1701859473
transform 1 0 4130 0 -1 7030
box -12 -8 32 272
use FILL  FILL_1__3162_
timestamp 1701859473
transform -1 0 4370 0 -1 7030
box -12 -8 32 272
use FILL  FILL_1__3163_
timestamp 1701859473
transform 1 0 4590 0 -1 7030
box -12 -8 32 272
use FILL  FILL_1__3164_
timestamp 1701859473
transform 1 0 4830 0 1 7030
box -12 -8 32 272
use FILL  FILL_1__3165_
timestamp 1701859473
transform 1 0 4090 0 1 7550
box -12 -8 32 272
use FILL  FILL_1__3166_
timestamp 1701859473
transform -1 0 4330 0 1 7550
box -12 -8 32 272
use FILL  FILL_1__3167_
timestamp 1701859473
transform 1 0 4810 0 -1 10150
box -12 -8 32 272
use FILL  FILL_1__3168_
timestamp 1701859473
transform 1 0 5010 0 -1 10150
box -12 -8 32 272
use FILL  FILL_1__3169_
timestamp 1701859473
transform -1 0 3650 0 -1 10670
box -12 -8 32 272
use FILL  FILL_1__3170_
timestamp 1701859473
transform -1 0 3870 0 -1 10670
box -12 -8 32 272
use FILL  FILL_1__3171_
timestamp 1701859473
transform 1 0 4290 0 -1 10670
box -12 -8 32 272
use FILL  FILL_1__3172_
timestamp 1701859473
transform -1 0 4530 0 -1 10670
box -12 -8 32 272
use FILL  FILL_1__3173_
timestamp 1701859473
transform 1 0 4130 0 1 10150
box -12 -8 32 272
use FILL  FILL_1__3174_
timestamp 1701859473
transform -1 0 4370 0 1 10150
box -12 -8 32 272
use FILL  FILL_1__3175_
timestamp 1701859473
transform 1 0 5470 0 1 10150
box -12 -8 32 272
use FILL  FILL_1__3176_
timestamp 1701859473
transform 1 0 5230 0 1 10150
box -12 -8 32 272
use FILL  FILL_1__3177_
timestamp 1701859473
transform -1 0 1710 0 -1 5990
box -12 -8 32 272
use FILL  FILL_1__3178_
timestamp 1701859473
transform 1 0 2150 0 -1 5990
box -12 -8 32 272
use FILL  FILL_1__3179_
timestamp 1701859473
transform -1 0 1430 0 1 6510
box -12 -8 32 272
use FILL  FILL_1__3180_
timestamp 1701859473
transform -1 0 1650 0 1 6510
box -12 -8 32 272
use FILL  FILL_1__3181_
timestamp 1701859473
transform -1 0 510 0 -1 6510
box -12 -8 32 272
use FILL  FILL_1__3182_
timestamp 1701859473
transform -1 0 910 0 -1 6510
box -12 -8 32 272
use FILL  FILL_1__3183_
timestamp 1701859473
transform 1 0 270 0 1 8070
box -12 -8 32 272
use FILL  FILL_1__3184_
timestamp 1701859473
transform -1 0 510 0 1 8070
box -12 -8 32 272
use FILL  FILL_1__3185_
timestamp 1701859473
transform -1 0 50 0 -1 8590
box -12 -8 32 272
use FILL  FILL_1__3186_
timestamp 1701859473
transform -1 0 50 0 1 8070
box -12 -8 32 272
use FILL  FILL_1__3187_
timestamp 1701859473
transform 1 0 670 0 -1 9110
box -12 -8 32 272
use FILL  FILL_1__3188_
timestamp 1701859473
transform 1 0 890 0 -1 9110
box -12 -8 32 272
use FILL  FILL_1__3189_
timestamp 1701859473
transform 1 0 2070 0 -1 9630
box -12 -8 32 272
use FILL  FILL_1__3190_
timestamp 1701859473
transform 1 0 2310 0 1 9110
box -12 -8 32 272
use FILL  FILL_1__3191_
timestamp 1701859473
transform 1 0 1370 0 -1 9110
box -12 -8 32 272
use FILL  FILL_1__3192_
timestamp 1701859473
transform -1 0 1610 0 -1 9110
box -12 -8 32 272
use FILL  FILL_1__3324_
timestamp 1701859473
transform 1 0 5550 0 1 8070
box -12 -8 32 272
use FILL  FILL_1__3325_
timestamp 1701859473
transform -1 0 6270 0 1 8070
box -12 -8 32 272
use FILL  FILL_1__3326_
timestamp 1701859473
transform -1 0 6170 0 -1 8070
box -12 -8 32 272
use FILL  FILL_1__3327_
timestamp 1701859473
transform -1 0 6130 0 -1 8590
box -12 -8 32 272
use FILL  FILL_1__3328_
timestamp 1701859473
transform -1 0 6030 0 1 8070
box -12 -8 32 272
use FILL  FILL_1__3329_
timestamp 1701859473
transform 1 0 5790 0 1 8070
box -12 -8 32 272
use FILL  FILL_1__3330_
timestamp 1701859473
transform -1 0 6970 0 1 8590
box -12 -8 32 272
use FILL  FILL_1__3331_
timestamp 1701859473
transform 1 0 7250 0 -1 8590
box -12 -8 32 272
use FILL  FILL_1__3332_
timestamp 1701859473
transform 1 0 6970 0 -1 8590
box -12 -8 32 272
use FILL  FILL_1__3333_
timestamp 1701859473
transform 1 0 10170 0 1 8590
box -12 -8 32 272
use FILL  FILL_1__3334_
timestamp 1701859473
transform 1 0 9290 0 1 8590
box -12 -8 32 272
use FILL  FILL_1__3335_
timestamp 1701859473
transform 1 0 7830 0 -1 10150
box -12 -8 32 272
use FILL  FILL_1__3336_
timestamp 1701859473
transform -1 0 6670 0 1 9630
box -12 -8 32 272
use FILL  FILL_1__3337_
timestamp 1701859473
transform -1 0 6190 0 1 9630
box -12 -8 32 272
use FILL  FILL_1__3338_
timestamp 1701859473
transform 1 0 7150 0 -1 10150
box -12 -8 32 272
use FILL  FILL_1__3339_
timestamp 1701859473
transform -1 0 8030 0 1 10150
box -12 -8 32 272
use FILL  FILL_1__3340_
timestamp 1701859473
transform 1 0 7790 0 1 10150
box -12 -8 32 272
use FILL  FILL_1__3341_
timestamp 1701859473
transform 1 0 7550 0 1 10150
box -12 -8 32 272
use FILL  FILL_1__3342_
timestamp 1701859473
transform 1 0 6770 0 -1 11190
box -12 -8 32 272
use FILL  FILL_1__3343_
timestamp 1701859473
transform -1 0 7370 0 -1 10150
box -12 -8 32 272
use FILL  FILL_1__3344_
timestamp 1701859473
transform 1 0 7590 0 -1 10150
box -12 -8 32 272
use FILL  FILL_1__3345_
timestamp 1701859473
transform -1 0 8970 0 1 9630
box -12 -8 32 272
use FILL  FILL_1__3346_
timestamp 1701859473
transform 1 0 8490 0 1 10150
box -12 -8 32 272
use FILL  FILL_1__3347_
timestamp 1701859473
transform -1 0 8270 0 1 10150
box -12 -8 32 272
use FILL  FILL_1__3348_
timestamp 1701859473
transform 1 0 9090 0 -1 10670
box -12 -8 32 272
use FILL  FILL_1__3349_
timestamp 1701859473
transform 1 0 7830 0 1 9630
box -12 -8 32 272
use FILL  FILL_1__3350_
timestamp 1701859473
transform 1 0 7530 0 -1 8590
box -12 -8 32 272
use FILL  FILL_1__3351_
timestamp 1701859473
transform -1 0 7710 0 1 8590
box -12 -8 32 272
use FILL  FILL_1__3352_
timestamp 1701859473
transform -1 0 8170 0 -1 9110
box -12 -8 32 272
use FILL  FILL_1__3353_
timestamp 1701859473
transform 1 0 8050 0 -1 10150
box -12 -8 32 272
use FILL  FILL_1__3354_
timestamp 1701859473
transform 1 0 7730 0 -1 10670
box -12 -8 32 272
use FILL  FILL_1__3355_
timestamp 1701859473
transform -1 0 7510 0 -1 10670
box -12 -8 32 272
use FILL  FILL_1__3356_
timestamp 1701859473
transform 1 0 7290 0 -1 10670
box -12 -8 32 272
use FILL  FILL_1__3357_
timestamp 1701859473
transform 1 0 7110 0 1 10670
box -12 -8 32 272
use FILL  FILL_1__3358_
timestamp 1701859473
transform 1 0 7370 0 1 10670
box -12 -8 32 272
use FILL  FILL_1__3359_
timestamp 1701859473
transform 1 0 7610 0 1 10670
box -12 -8 32 272
use FILL  FILL_1__3360_
timestamp 1701859473
transform -1 0 7870 0 1 10670
box -12 -8 32 272
use FILL  FILL_1__3361_
timestamp 1701859473
transform 1 0 8890 0 -1 10670
box -12 -8 32 272
use FILL  FILL_1__3362_
timestamp 1701859473
transform 1 0 7950 0 -1 10670
box -12 -8 32 272
use FILL  FILL_1__3363_
timestamp 1701859473
transform 1 0 8070 0 1 10670
box -12 -8 32 272
use FILL  FILL_1__3364_
timestamp 1701859473
transform 1 0 7910 0 -1 11190
box -12 -8 32 272
use FILL  FILL_1__3365_
timestamp 1701859473
transform -1 0 7450 0 -1 11190
box -12 -8 32 272
use FILL  FILL_1__3366_
timestamp 1701859473
transform 1 0 6970 0 -1 11190
box -12 -8 32 272
use FILL  FILL_1__3367_
timestamp 1701859473
transform 1 0 6850 0 1 10670
box -12 -8 32 272
use FILL  FILL_1__3368_
timestamp 1701859473
transform 1 0 7190 0 -1 11190
box -12 -8 32 272
use FILL  FILL_1__3369_
timestamp 1701859473
transform 1 0 7670 0 -1 11190
box -12 -8 32 272
use FILL  FILL_1__3370_
timestamp 1701859473
transform 1 0 8190 0 -1 10670
box -12 -8 32 272
use FILL  FILL_1__3371_
timestamp 1701859473
transform 1 0 8290 0 1 10670
box -12 -8 32 272
use FILL  FILL_1__3372_
timestamp 1701859473
transform 1 0 9470 0 1 10670
box -12 -8 32 272
use FILL  FILL_1__3373_
timestamp 1701859473
transform -1 0 6570 0 -1 11190
box -12 -8 32 272
use FILL  FILL_1__3374_
timestamp 1701859473
transform 1 0 5670 0 1 10670
box -12 -8 32 272
use FILL  FILL_1__3375_
timestamp 1701859473
transform -1 0 5930 0 1 10670
box -12 -8 32 272
use FILL  FILL_1__3376_
timestamp 1701859473
transform -1 0 6150 0 1 10670
box -12 -8 32 272
use FILL  FILL_1__3377_
timestamp 1701859473
transform 1 0 6390 0 1 10670
box -12 -8 32 272
use FILL  FILL_1__3378_
timestamp 1701859473
transform 1 0 6330 0 -1 11190
box -12 -8 32 272
use FILL  FILL_1__3379_
timestamp 1701859473
transform 1 0 8650 0 -1 10670
box -12 -8 32 272
use FILL  FILL_1__3380_
timestamp 1701859473
transform 1 0 8770 0 1 10670
box -12 -8 32 272
use FILL  FILL_1__3381_
timestamp 1701859473
transform -1 0 6650 0 1 10670
box -12 -8 32 272
use FILL  FILL_1__3382_
timestamp 1701859473
transform 1 0 6110 0 -1 10670
box -12 -8 32 272
use FILL  FILL_1__3383_
timestamp 1701859473
transform -1 0 6370 0 -1 10670
box -12 -8 32 272
use FILL  FILL_1__3384_
timestamp 1701859473
transform -1 0 6810 0 -1 10670
box -12 -8 32 272
use FILL  FILL_1__3385_
timestamp 1701859473
transform 1 0 6570 0 -1 10670
box -12 -8 32 272
use FILL  FILL_1__3386_
timestamp 1701859473
transform 1 0 7050 0 -1 10670
box -12 -8 32 272
use FILL  FILL_1__3387_
timestamp 1701859473
transform 1 0 8410 0 -1 10670
box -12 -8 32 272
use FILL  FILL_1__3388_
timestamp 1701859473
transform 1 0 8530 0 1 10670
box -12 -8 32 272
use FILL  FILL_1__3389_
timestamp 1701859473
transform 1 0 10190 0 -1 10670
box -12 -8 32 272
use FILL  FILL_1__3390_
timestamp 1701859473
transform 1 0 9750 0 -1 10670
box -12 -8 32 272
use FILL  FILL_1__3391_
timestamp 1701859473
transform 1 0 9950 0 -1 10670
box -12 -8 32 272
use FILL  FILL_1__3392_
timestamp 1701859473
transform 1 0 10410 0 -1 10670
box -12 -8 32 272
use FILL  FILL_1__3393_
timestamp 1701859473
transform -1 0 11150 0 -1 10150
box -12 -8 32 272
use FILL  FILL_1__3394_
timestamp 1701859473
transform 1 0 7330 0 1 10150
box -12 -8 32 272
use FILL  FILL_1__3395_
timestamp 1701859473
transform 1 0 6390 0 1 10150
box -12 -8 32 272
use FILL  FILL_1__3396_
timestamp 1701859473
transform -1 0 6650 0 1 10150
box -12 -8 32 272
use FILL  FILL_1__3397_
timestamp 1701859473
transform -1 0 6970 0 -1 10150
box -12 -8 32 272
use FILL  FILL_1__3398_
timestamp 1701859473
transform 1 0 6250 0 -1 10150
box -12 -8 32 272
use FILL  FILL_1__3399_
timestamp 1701859473
transform -1 0 6730 0 -1 10150
box -12 -8 32 272
use FILL  FILL_1__3400_
timestamp 1701859473
transform -1 0 6910 0 1 10150
box -12 -8 32 272
use FILL  FILL_1__3401_
timestamp 1701859473
transform 1 0 7090 0 1 10150
box -12 -8 32 272
use FILL  FILL_1__3402_
timestamp 1701859473
transform -1 0 9030 0 1 10150
box -12 -8 32 272
use FILL  FILL_1__3403_
timestamp 1701859473
transform 1 0 9470 0 1 10150
box -12 -8 32 272
use FILL  FILL_1__3404_
timestamp 1701859473
transform -1 0 5730 0 1 9630
box -12 -8 32 272
use FILL  FILL_1__3405_
timestamp 1701859473
transform -1 0 6010 0 -1 10150
box -12 -8 32 272
use FILL  FILL_1__3406_
timestamp 1701859473
transform 1 0 6370 0 -1 9630
box -12 -8 32 272
use FILL  FILL_1__3407_
timestamp 1701859473
transform -1 0 6590 0 -1 9630
box -12 -8 32 272
use FILL  FILL_1__3408_
timestamp 1701859473
transform 1 0 6850 0 1 9630
box -12 -8 32 272
use FILL  FILL_1__3409_
timestamp 1701859473
transform -1 0 6470 0 -1 10150
box -12 -8 32 272
use FILL  FILL_1__3410_
timestamp 1701859473
transform 1 0 9210 0 -1 10150
box -12 -8 32 272
use FILL  FILL_1__3411_
timestamp 1701859473
transform 1 0 9230 0 1 10150
box -12 -8 32 272
use FILL  FILL_1__3412_
timestamp 1701859473
transform 1 0 9950 0 1 10150
box -12 -8 32 272
use FILL  FILL_1__3413_
timestamp 1701859473
transform -1 0 5970 0 1 9630
box -12 -8 32 272
use FILL  FILL_1__3414_
timestamp 1701859473
transform 1 0 8110 0 1 9110
box -12 -8 32 272
use FILL  FILL_1__3415_
timestamp 1701859473
transform 1 0 6390 0 1 9630
box -12 -8 32 272
use FILL  FILL_1__3416_
timestamp 1701859473
transform 1 0 7230 0 1 8590
box -12 -8 32 272
use FILL  FILL_1__3417_
timestamp 1701859473
transform 1 0 7310 0 -1 9110
box -12 -8 32 272
use FILL  FILL_1__3418_
timestamp 1701859473
transform -1 0 7450 0 -1 9630
box -12 -8 32 272
use FILL  FILL_1__3419_
timestamp 1701859473
transform 1 0 7210 0 -1 9630
box -12 -8 32 272
use FILL  FILL_1__3420_
timestamp 1701859473
transform -1 0 6790 0 -1 9630
box -12 -8 32 272
use FILL  FILL_1__3421_
timestamp 1701859473
transform -1 0 7010 0 -1 9630
box -12 -8 32 272
use FILL  FILL_1__3422_
timestamp 1701859473
transform -1 0 7110 0 1 9630
box -12 -8 32 272
use FILL  FILL_1__3423_
timestamp 1701859473
transform -1 0 8170 0 -1 9630
box -12 -8 32 272
use FILL  FILL_1__3424_
timestamp 1701859473
transform -1 0 7690 0 -1 9630
box -12 -8 32 272
use FILL  FILL_1__3425_
timestamp 1701859473
transform -1 0 7350 0 1 9630
box -12 -8 32 272
use FILL  FILL_1__3426_
timestamp 1701859473
transform -1 0 8990 0 -1 10150
box -12 -8 32 272
use FILL  FILL_1__3427_
timestamp 1701859473
transform 1 0 8750 0 -1 10150
box -12 -8 32 272
use FILL  FILL_1__3428_
timestamp 1701859473
transform 1 0 7430 0 1 8590
box -12 -8 32 272
use FILL  FILL_1__3429_
timestamp 1701859473
transform 1 0 7510 0 -1 9110
box -12 -8 32 272
use FILL  FILL_1__3430_
timestamp 1701859473
transform -1 0 7730 0 -1 9110
box -12 -8 32 272
use FILL  FILL_1__3431_
timestamp 1701859473
transform 1 0 7650 0 1 9110
box -12 -8 32 272
use FILL  FILL_1__3432_
timestamp 1701859473
transform 1 0 7890 0 1 9110
box -12 -8 32 272
use FILL  FILL_1__3433_
timestamp 1701859473
transform -1 0 7930 0 -1 9630
box -12 -8 32 272
use FILL  FILL_1__3434_
timestamp 1701859473
transform 1 0 7570 0 1 9630
box -12 -8 32 272
use FILL  FILL_1__3435_
timestamp 1701859473
transform 1 0 10190 0 1 10150
box -12 -8 32 272
use FILL  FILL_1__3436_
timestamp 1701859473
transform -1 0 10190 0 -1 10150
box -12 -8 32 272
use FILL  FILL_1__3437_
timestamp 1701859473
transform 1 0 10630 0 1 10150
box -12 -8 32 272
use FILL  FILL_1__3438_
timestamp 1701859473
transform 1 0 10410 0 1 10150
box -12 -8 32 272
use FILL  FILL_1__3439_
timestamp 1701859473
transform 1 0 10850 0 1 10150
box -12 -8 32 272
use FILL  FILL_1__3440_
timestamp 1701859473
transform -1 0 10670 0 -1 10150
box -12 -8 32 272
use FILL  FILL_1__3441_
timestamp 1701859473
transform -1 0 10530 0 1 9630
box -12 -8 32 272
use FILL  FILL_1__3442_
timestamp 1701859473
transform -1 0 10410 0 -1 10150
box -12 -8 32 272
use FILL  FILL_1__3443_
timestamp 1701859473
transform -1 0 10970 0 1 9630
box -12 -8 32 272
use FILL  FILL_1__3444_
timestamp 1701859473
transform -1 0 8370 0 -1 9630
box -12 -8 32 272
use FILL  FILL_1__3445_
timestamp 1701859473
transform -1 0 8070 0 1 9630
box -12 -8 32 272
use FILL  FILL_1__3446_
timestamp 1701859473
transform 1 0 8510 0 1 9630
box -12 -8 32 272
use FILL  FILL_1__3447_
timestamp 1701859473
transform 1 0 8290 0 1 9630
box -12 -8 32 272
use FILL  FILL_1__3448_
timestamp 1701859473
transform -1 0 8730 0 1 9630
box -12 -8 32 272
use FILL  FILL_1__3449_
timestamp 1701859473
transform -1 0 9770 0 1 10150
box -12 -8 32 272
use FILL  FILL_1__3450_
timestamp 1701859473
transform -1 0 9730 0 -1 10150
box -12 -8 32 272
use FILL  FILL_1__3451_
timestamp 1701859473
transform 1 0 9450 0 -1 10150
box -12 -8 32 272
use FILL  FILL_1__3452_
timestamp 1701859473
transform -1 0 9190 0 1 9630
box -12 -8 32 272
use FILL  FILL_1__3453_
timestamp 1701859473
transform -1 0 9950 0 -1 10150
box -12 -8 32 272
use FILL  FILL_1__3454_
timestamp 1701859473
transform 1 0 9390 0 1 9630
box -12 -8 32 272
use FILL  FILL_1__3455_
timestamp 1701859473
transform 1 0 9610 0 1 9630
box -12 -8 32 272
use FILL  FILL_1__3456_
timestamp 1701859473
transform -1 0 10310 0 1 9630
box -12 -8 32 272
use FILL  FILL_1__3457_
timestamp 1701859473
transform -1 0 9850 0 1 9630
box -12 -8 32 272
use FILL  FILL_1__3458_
timestamp 1701859473
transform -1 0 10090 0 1 9630
box -12 -8 32 272
use FILL  FILL_1__3459_
timestamp 1701859473
transform -1 0 10230 0 -1 9630
box -12 -8 32 272
use FILL  FILL_1__3460_
timestamp 1701859473
transform 1 0 10890 0 -1 10150
box -12 -8 32 272
use FILL  FILL_1__3461_
timestamp 1701859473
transform -1 0 11130 0 -1 9630
box -12 -8 32 272
use FILL  FILL_1__3462_
timestamp 1701859473
transform -1 0 10670 0 -1 9630
box -12 -8 32 272
use FILL  FILL_1__3463_
timestamp 1701859473
transform 1 0 10350 0 -1 11190
box -12 -8 32 272
use FILL  FILL_1__3464_
timestamp 1701859473
transform 1 0 9690 0 -1 11190
box -12 -8 32 272
use FILL  FILL_1__3465_
timestamp 1701859473
transform 1 0 9930 0 -1 11190
box -12 -8 32 272
use FILL  FILL_1__3466_
timestamp 1701859473
transform 1 0 10110 0 -1 11190
box -12 -8 32 272
use FILL  FILL_1__3467_
timestamp 1701859473
transform -1 0 11090 0 1 10670
box -12 -8 32 272
use FILL  FILL_1__3468_
timestamp 1701859473
transform 1 0 10590 0 1 10670
box -12 -8 32 272
use FILL  FILL_1__3469_
timestamp 1701859473
transform 1 0 9310 0 -1 10670
box -12 -8 32 272
use FILL  FILL_1__3470_
timestamp 1701859473
transform 1 0 9550 0 -1 10670
box -12 -8 32 272
use FILL  FILL_1__3471_
timestamp 1701859473
transform 1 0 9690 0 1 10670
box -12 -8 32 272
use FILL  FILL_1__3472_
timestamp 1701859473
transform -1 0 9950 0 1 10670
box -12 -8 32 272
use FILL  FILL_1__3473_
timestamp 1701859473
transform 1 0 8570 0 -1 11190
box -12 -8 32 272
use FILL  FILL_1__3474_
timestamp 1701859473
transform 1 0 8130 0 -1 11190
box -12 -8 32 272
use FILL  FILL_1__3475_
timestamp 1701859473
transform 1 0 8370 0 -1 11190
box -12 -8 32 272
use FILL  FILL_1__3476_
timestamp 1701859473
transform -1 0 8810 0 -1 11190
box -12 -8 32 272
use FILL  FILL_1__3477_
timestamp 1701859473
transform 1 0 9030 0 -1 11190
box -12 -8 32 272
use FILL  FILL_1__3478_
timestamp 1701859473
transform 1 0 9010 0 1 10670
box -12 -8 32 272
use FILL  FILL_1__3479_
timestamp 1701859473
transform 1 0 8290 0 -1 10150
box -12 -8 32 272
use FILL  FILL_1__3480_
timestamp 1701859473
transform -1 0 8550 0 -1 10150
box -12 -8 32 272
use FILL  FILL_1__3481_
timestamp 1701859473
transform -1 0 8330 0 1 9110
box -12 -8 32 272
use FILL  FILL_1__3482_
timestamp 1701859473
transform -1 0 8550 0 1 9110
box -12 -8 32 272
use FILL  FILL_1__3483_
timestamp 1701859473
transform 1 0 8730 0 1 10150
box -12 -8 32 272
use FILL  FILL_1__3484_
timestamp 1701859473
transform -1 0 10030 0 -1 9630
box -12 -8 32 272
use FILL  FILL_1__3485_
timestamp 1701859473
transform 1 0 11050 0 1 10150
box -12 -8 32 272
use FILL  FILL_1__3486_
timestamp 1701859473
transform 1 0 10390 0 1 9110
box -12 -8 32 272
use FILL  FILL_1__3487_
timestamp 1701859473
transform 1 0 10430 0 -1 9630
box -12 -8 32 272
use FILL  FILL_1__3488_
timestamp 1701859473
transform -1 0 10730 0 1 9630
box -12 -8 32 272
use FILL  FILL_1__3489_
timestamp 1701859473
transform 1 0 10570 0 -1 11190
box -12 -8 32 272
use FILL  FILL_1__3490_
timestamp 1701859473
transform 1 0 11030 0 -1 11190
box -12 -8 32 272
use FILL  FILL_1__3491_
timestamp 1701859473
transform -1 0 10830 0 -1 11190
box -12 -8 32 272
use FILL  FILL_1__3492_
timestamp 1701859473
transform -1 0 10390 0 1 10670
box -12 -8 32 272
use FILL  FILL_1__3493_
timestamp 1701859473
transform -1 0 10170 0 1 10670
box -12 -8 32 272
use FILL  FILL_1__3494_
timestamp 1701859473
transform 1 0 9270 0 1 10670
box -12 -8 32 272
use FILL  FILL_1__3495_
timestamp 1701859473
transform -1 0 9470 0 -1 11190
box -12 -8 32 272
use FILL  FILL_1__3496_
timestamp 1701859473
transform 1 0 9230 0 -1 11190
box -12 -8 32 272
use FILL  FILL_1__3497_
timestamp 1701859473
transform -1 0 9330 0 -1 9630
box -12 -8 32 272
use FILL  FILL_1__3498_
timestamp 1701859473
transform -1 0 8830 0 1 9110
box -12 -8 32 272
use FILL  FILL_1__3499_
timestamp 1701859473
transform 1 0 8350 0 -1 9110
box -12 -8 32 272
use FILL  FILL_1__3500_
timestamp 1701859473
transform 1 0 9730 0 1 9110
box -12 -8 32 272
use FILL  FILL_1__3501_
timestamp 1701859473
transform -1 0 9970 0 1 9110
box -12 -8 32 272
use FILL  FILL_1__3502_
timestamp 1701859473
transform -1 0 8230 0 -1 8590
box -12 -8 32 272
use FILL  FILL_1__3503_
timestamp 1701859473
transform -1 0 8610 0 -1 9630
box -12 -8 32 272
use FILL  FILL_1__3504_
timestamp 1701859473
transform 1 0 8830 0 -1 9630
box -12 -8 32 272
use FILL  FILL_1__3505_
timestamp 1701859473
transform -1 0 9090 0 -1 9630
box -12 -8 32 272
use FILL  FILL_1__3506_
timestamp 1701859473
transform -1 0 8610 0 1 8590
box -12 -8 32 272
use FILL  FILL_1__3507_
timestamp 1701859473
transform 1 0 10690 0 -1 9110
box -12 -8 32 272
use FILL  FILL_1__3508_
timestamp 1701859473
transform 1 0 10450 0 -1 9110
box -12 -8 32 272
use FILL  FILL_1__3509_
timestamp 1701859473
transform 1 0 8390 0 1 8590
box -12 -8 32 272
use FILL  FILL_1__3510_
timestamp 1701859473
transform -1 0 8850 0 1 8590
box -12 -8 32 272
use FILL  FILL_1__3511_
timestamp 1701859473
transform 1 0 9910 0 -1 270
box -12 -8 32 272
use FILL  FILL_1__3512_
timestamp 1701859473
transform 1 0 10910 0 -1 9110
box -12 -8 32 272
use FILL  FILL_1__3513_
timestamp 1701859473
transform 1 0 10890 0 -1 9630
box -12 -8 32 272
use FILL  FILL_1__3514_
timestamp 1701859473
transform 1 0 10850 0 1 10670
box -12 -8 32 272
use FILL  FILL_1__3515_
timestamp 1701859473
transform -1 0 10650 0 -1 10670
box -12 -8 32 272
use FILL  FILL_1__3516_
timestamp 1701859473
transform 1 0 10870 0 -1 10670
box -12 -8 32 272
use FILL  FILL_1__3517_
timestamp 1701859473
transform 1 0 9550 0 -1 9630
box -12 -8 32 272
use FILL  FILL_1__3518_
timestamp 1701859473
transform 1 0 9770 0 -1 9630
box -12 -8 32 272
use FILL  FILL_1__3519_
timestamp 1701859473
transform 1 0 9050 0 1 9110
box -12 -8 32 272
use FILL  FILL_1__3520_
timestamp 1701859473
transform -1 0 9290 0 1 9110
box -12 -8 32 272
use FILL  FILL_1__3521_
timestamp 1701859473
transform 1 0 6530 0 1 8590
box -12 -8 32 272
use FILL  FILL_1__3522_
timestamp 1701859473
transform 1 0 7930 0 -1 9110
box -12 -8 32 272
use FILL  FILL_1__3523_
timestamp 1701859473
transform 1 0 6730 0 1 8590
box -12 -8 32 272
use FILL  FILL_1__3524_
timestamp 1701859473
transform 1 0 7450 0 1 9110
box -12 -8 32 272
use FILL  FILL_1__3525_
timestamp 1701859473
transform 1 0 6990 0 1 9110
box -12 -8 32 272
use FILL  FILL_1__3526_
timestamp 1701859473
transform -1 0 7230 0 1 9110
box -12 -8 32 272
use FILL  FILL_1__3539_
timestamp 1701859473
transform 1 0 11090 0 -1 7030
box -12 -8 32 272
use FILL  FILL_1__3540_
timestamp 1701859473
transform 1 0 4590 0 1 10670
box -12 -8 32 272
use FILL  FILL_1__3541_
timestamp 1701859473
transform -1 0 50 0 1 5990
box -12 -8 32 272
use FILL  FILL_1__3542_
timestamp 1701859473
transform -1 0 50 0 -1 8070
box -12 -8 32 272
use FILL  FILL_1__3543_
timestamp 1701859473
transform -1 0 50 0 1 8590
box -12 -8 32 272
use FILL  FILL_1__3544_
timestamp 1701859473
transform -1 0 50 0 1 9110
box -12 -8 32 272
use FILL  FILL_1__3545_
timestamp 1701859473
transform -1 0 1890 0 -1 11190
box -12 -8 32 272
use FILL  FILL_1__3546_
timestamp 1701859473
transform -1 0 510 0 1 9110
box -12 -8 32 272
use FILL  FILL_1__3547_
timestamp 1701859473
transform 1 0 4630 0 -1 11190
box -12 -8 32 272
use FILL  FILL_1__3548_
timestamp 1701859473
transform 1 0 5230 0 1 10670
box -12 -8 32 272
use FILL  FILL_1__3549_
timestamp 1701859473
transform -1 0 4230 0 -1 11190
box -12 -8 32 272
use FILL  FILL_1__3550_
timestamp 1701859473
transform -1 0 5070 0 -1 11190
box -12 -8 32 272
use FILL  FILL_1__3551_
timestamp 1701859473
transform 1 0 5470 0 -1 11190
box -12 -8 32 272
use FILL  FILL_1__3552_
timestamp 1701859473
transform 1 0 5250 0 -1 11190
box -12 -8 32 272
use FILL  FILL_1__3553_
timestamp 1701859473
transform -1 0 50 0 -1 5990
box -12 -8 32 272
use FILL  FILL_1__3554_
timestamp 1701859473
transform -1 0 250 0 1 7030
box -12 -8 32 272
use FILL  FILL_1__3555_
timestamp 1701859473
transform -1 0 5030 0 1 10670
box -12 -8 32 272
use FILL  FILL_1__3556_
timestamp 1701859473
transform 1 0 6170 0 1 10150
box -12 -8 32 272
use FILL  FILL_1__3557_
timestamp 1701859473
transform -1 0 5710 0 -1 11190
box -12 -8 32 272
use FILL  FILL_1__3558_
timestamp 1701859473
transform 1 0 6110 0 -1 11190
box -12 -8 32 272
use FILL  FILL_1__3559_
timestamp 1701859473
transform -1 0 4770 0 -1 10670
box -12 -8 32 272
use FILL  FILL_1__3560_
timestamp 1701859473
transform 1 0 5450 0 1 10670
box -12 -8 32 272
use FILL  FILL_1__3561_
timestamp 1701859473
transform 1 0 5890 0 -1 11190
box -12 -8 32 272
use FILL  FILL_1__3562_
timestamp 1701859473
transform 1 0 5690 0 1 10150
box -12 -8 32 272
use FILL  FILL_1__3563_
timestamp 1701859473
transform 1 0 5150 0 1 3390
box -12 -8 32 272
use FILL  FILL_1_BUFX2_insert0
timestamp 1701859473
transform 1 0 5770 0 -1 10150
box -12 -8 32 272
use FILL  FILL_1_BUFX2_insert1
timestamp 1701859473
transform 1 0 6530 0 1 2350
box -12 -8 32 272
use FILL  FILL_1_BUFX2_insert2
timestamp 1701859473
transform 1 0 5370 0 -1 1830
box -12 -8 32 272
use FILL  FILL_1_BUFX2_insert3
timestamp 1701859473
transform -1 0 510 0 -1 5470
box -12 -8 32 272
use FILL  FILL_1_BUFX2_insert4
timestamp 1701859473
transform 1 0 3250 0 1 4950
box -12 -8 32 272
use FILL  FILL_1_BUFX2_insert5
timestamp 1701859473
transform 1 0 1310 0 -1 1830
box -12 -8 32 272
use FILL  FILL_1_BUFX2_insert6
timestamp 1701859473
transform -1 0 50 0 -1 11190
box -12 -8 32 272
use FILL  FILL_1_BUFX2_insert7
timestamp 1701859473
transform 1 0 1610 0 1 10670
box -12 -8 32 272
use FILL  FILL_1_BUFX2_insert8
timestamp 1701859473
transform 1 0 1570 0 1 1830
box -12 -8 32 272
use FILL  FILL_1_BUFX2_insert9
timestamp 1701859473
transform 1 0 1870 0 -1 3910
box -12 -8 32 272
use FILL  FILL_1_BUFX2_insert10
timestamp 1701859473
transform 1 0 1690 0 -1 4430
box -12 -8 32 272
use FILL  FILL_1_BUFX2_insert11
timestamp 1701859473
transform -1 0 1670 0 -1 3910
box -12 -8 32 272
use FILL  FILL_1_BUFX2_insert12
timestamp 1701859473
transform -1 0 1450 0 -1 3910
box -12 -8 32 272
use FILL  FILL_1_BUFX2_insert13
timestamp 1701859473
transform -1 0 1350 0 -1 1310
box -12 -8 32 272
use FILL  FILL_1_BUFX2_insert14
timestamp 1701859473
transform -1 0 3590 0 1 3390
box -12 -8 32 272
use FILL  FILL_1_BUFX2_insert15
timestamp 1701859473
transform 1 0 4470 0 -1 5470
box -12 -8 32 272
use FILL  FILL_1_BUFX2_insert16
timestamp 1701859473
transform 1 0 1270 0 -1 4950
box -12 -8 32 272
use FILL  FILL_1_BUFX2_insert17
timestamp 1701859473
transform 1 0 3550 0 1 1310
box -12 -8 32 272
use FILL  FILL_1_BUFX2_insert18
timestamp 1701859473
transform -1 0 9690 0 1 2350
box -12 -8 32 272
use FILL  FILL_1_BUFX2_insert19
timestamp 1701859473
transform -1 0 8430 0 -1 790
box -12 -8 32 272
use FILL  FILL_1_BUFX2_insert20
timestamp 1701859473
transform 1 0 9890 0 1 2350
box -12 -8 32 272
use FILL  FILL_1_BUFX2_insert21
timestamp 1701859473
transform -1 0 7730 0 -1 1310
box -12 -8 32 272
use FILL  FILL_1_BUFX2_insert22
timestamp 1701859473
transform -1 0 3130 0 -1 2870
box -12 -8 32 272
use FILL  FILL_1_BUFX2_insert23
timestamp 1701859473
transform -1 0 2670 0 -1 4950
box -12 -8 32 272
use FILL  FILL_1_BUFX2_insert24
timestamp 1701859473
transform -1 0 3570 0 -1 4430
box -12 -8 32 272
use FILL  FILL_1_BUFX2_insert25
timestamp 1701859473
transform 1 0 4310 0 1 4430
box -12 -8 32 272
use FILL  FILL_1_BUFX2_insert26
timestamp 1701859473
transform 1 0 4130 0 1 2870
box -12 -8 32 272
use FILL  FILL_1_BUFX2_insert27
timestamp 1701859473
transform 1 0 9530 0 1 4950
box -12 -8 32 272
use FILL  FILL_1_BUFX2_insert28
timestamp 1701859473
transform -1 0 7410 0 -1 5990
box -12 -8 32 272
use FILL  FILL_1_BUFX2_insert29
timestamp 1701859473
transform -1 0 1210 0 1 6510
box -12 -8 32 272
use FILL  FILL_1_BUFX2_insert30
timestamp 1701859473
transform -1 0 8710 0 -1 3910
box -12 -8 32 272
use FILL  FILL_1_BUFX2_insert31
timestamp 1701859473
transform -1 0 9490 0 1 3910
box -12 -8 32 272
use FILL  FILL_1_BUFX2_insert32
timestamp 1701859473
transform 1 0 5790 0 -1 3910
box -12 -8 32 272
use FILL  FILL_1_BUFX2_insert33
timestamp 1701859473
transform -1 0 9470 0 -1 4950
box -12 -8 32 272
use FILL  FILL_1_BUFX2_insert34
timestamp 1701859473
transform 1 0 5130 0 1 8590
box -12 -8 32 272
use FILL  FILL_1_BUFX2_insert35
timestamp 1701859473
transform -1 0 5890 0 1 7550
box -12 -8 32 272
use FILL  FILL_1_BUFX2_insert36
timestamp 1701859473
transform -1 0 1130 0 1 8590
box -12 -8 32 272
use FILL  FILL_1_BUFX2_insert37
timestamp 1701859473
transform -1 0 9510 0 1 8590
box -12 -8 32 272
use FILL  FILL_1_BUFX2_insert49
timestamp 1701859473
transform -1 0 2970 0 1 6510
box -12 -8 32 272
use FILL  FILL_1_BUFX2_insert50
timestamp 1701859473
transform 1 0 2270 0 -1 8590
box -12 -8 32 272
use FILL  FILL_1_BUFX2_insert51
timestamp 1701859473
transform 1 0 3130 0 -1 8590
box -12 -8 32 272
use FILL  FILL_1_BUFX2_insert52
timestamp 1701859473
transform 1 0 3310 0 1 5470
box -12 -8 32 272
use FILL  FILL_1_BUFX2_insert53
timestamp 1701859473
transform -1 0 11150 0 1 9110
box -12 -8 32 272
use FILL  FILL_1_BUFX2_insert54
timestamp 1701859473
transform -1 0 9090 0 1 8590
box -12 -8 32 272
use FILL  FILL_1_BUFX2_insert55
timestamp 1701859473
transform -1 0 9530 0 1 9110
box -12 -8 32 272
use FILL  FILL_1_BUFX2_insert56
timestamp 1701859473
transform -1 0 10190 0 1 9110
box -12 -8 32 272
use FILL  FILL_1_BUFX2_insert57
timestamp 1701859473
transform -1 0 11150 0 -1 2350
box -12 -8 32 272
use FILL  FILL_1_BUFX2_insert58
timestamp 1701859473
transform -1 0 8890 0 1 2870
box -12 -8 32 272
use FILL  FILL_1_BUFX2_insert59
timestamp 1701859473
transform -1 0 7470 0 1 1830
box -12 -8 32 272
use FILL  FILL_1_BUFX2_insert60
timestamp 1701859473
transform 1 0 10810 0 1 1830
box -12 -8 32 272
use FILL  FILL_1_BUFX2_insert61
timestamp 1701859473
transform -1 0 11090 0 1 2870
box -12 -8 32 272
use FILL  FILL_1_BUFX2_insert62
timestamp 1701859473
transform 1 0 2130 0 1 3910
box -12 -8 32 272
use FILL  FILL_1_BUFX2_insert63
timestamp 1701859473
transform 1 0 2050 0 1 3390
box -12 -8 32 272
use FILL  FILL_1_BUFX2_insert64
timestamp 1701859473
transform -1 0 1710 0 1 3910
box -12 -8 32 272
use FILL  FILL_1_BUFX2_insert65
timestamp 1701859473
transform -1 0 1650 0 1 3390
box -12 -8 32 272
use FILL  FILL_1_BUFX2_insert66
timestamp 1701859473
transform -1 0 4230 0 1 1310
box -12 -8 32 272
use FILL  FILL_1_BUFX2_insert67
timestamp 1701859473
transform -1 0 3530 0 -1 10150
box -12 -8 32 272
use FILL  FILL_1_BUFX2_insert68
timestamp 1701859473
transform -1 0 7090 0 1 2870
box -12 -8 32 272
use FILL  FILL_1_BUFX2_insert69
timestamp 1701859473
transform -1 0 5570 0 -1 3390
box -12 -8 32 272
use FILL  FILL_1_BUFX2_insert70
timestamp 1701859473
transform -1 0 3590 0 -1 1830
box -12 -8 32 272
use FILL  FILL_1_BUFX2_insert71
timestamp 1701859473
transform -1 0 7230 0 1 2350
box -12 -8 32 272
use FILL  FILL_1_BUFX2_insert72
timestamp 1701859473
transform -1 0 6410 0 1 1310
box -12 -8 32 272
use FILL  FILL_1_BUFX2_insert73
timestamp 1701859473
transform 1 0 3530 0 1 5470
box -12 -8 32 272
use FILL  FILL_1_BUFX2_insert74
timestamp 1701859473
transform 1 0 7490 0 -1 2350
box -12 -8 32 272
use FILL  FILL_1_BUFX2_insert75
timestamp 1701859473
transform 1 0 7510 0 1 2870
box -12 -8 32 272
use FILL  FILL_1_BUFX2_insert76
timestamp 1701859473
transform 1 0 7290 0 1 2870
box -12 -8 32 272
use FILL  FILL_1_BUFX2_insert77
timestamp 1701859473
transform -1 0 3350 0 -1 2870
box -12 -8 32 272
use FILL  FILL_1_BUFX2_insert78
timestamp 1701859473
transform 1 0 1850 0 -1 2870
box -12 -8 32 272
use FILL  FILL_1_BUFX2_insert79
timestamp 1701859473
transform -1 0 2090 0 -1 2870
box -12 -8 32 272
use FILL  FILL_1_BUFX2_insert80
timestamp 1701859473
transform 1 0 2330 0 1 4430
box -12 -8 32 272
use FILL  FILL_1_BUFX2_insert81
timestamp 1701859473
transform -1 0 1930 0 1 3910
box -12 -8 32 272
use FILL  FILL_1_BUFX2_insert82
timestamp 1701859473
transform -1 0 250 0 1 8590
box -12 -8 32 272
use FILL  FILL_1_BUFX2_insert83
timestamp 1701859473
transform 1 0 4130 0 -1 10150
box -12 -8 32 272
use FILL  FILL_1_BUFX2_insert84
timestamp 1701859473
transform 1 0 4090 0 -1 7550
box -12 -8 32 272
use FILL  FILL_1_BUFX2_insert85
timestamp 1701859473
transform -1 0 50 0 -1 6510
box -12 -8 32 272
use FILL  FILL_1_BUFX2_insert86
timestamp 1701859473
transform 1 0 1850 0 -1 10150
box -12 -8 32 272
use FILL  FILL_1_CLKBUF1_insert38
timestamp 1701859473
transform 1 0 2850 0 -1 7550
box -12 -8 32 272
use FILL  FILL_1_CLKBUF1_insert39
timestamp 1701859473
transform -1 0 4650 0 -1 6510
box -12 -8 32 272
use FILL  FILL_1_CLKBUF1_insert40
timestamp 1701859473
transform -1 0 950 0 -1 4950
box -12 -8 32 272
use FILL  FILL_1_CLKBUF1_insert41
timestamp 1701859473
transform -1 0 10610 0 -1 270
box -12 -8 32 272
use FILL  FILL_1_CLKBUF1_insert42
timestamp 1701859473
transform 1 0 9670 0 -1 4950
box -12 -8 32 272
use FILL  FILL_1_CLKBUF1_insert43
timestamp 1701859473
transform -1 0 10990 0 1 7030
box -12 -8 32 272
use FILL  FILL_1_CLKBUF1_insert44
timestamp 1701859473
transform -1 0 10730 0 1 4430
box -12 -8 32 272
use FILL  FILL_1_CLKBUF1_insert45
timestamp 1701859473
transform 1 0 5650 0 -1 6510
box -12 -8 32 272
use FILL  FILL_1_CLKBUF1_insert46
timestamp 1701859473
transform 1 0 3970 0 1 5990
box -12 -8 32 272
use FILL  FILL_1_CLKBUF1_insert47
timestamp 1701859473
transform -1 0 2090 0 1 7550
box -12 -8 32 272
use FILL  FILL_1_CLKBUF1_insert48
timestamp 1701859473
transform -1 0 10770 0 -1 7030
box -12 -8 32 272
use FILL  FILL_2__1668_
timestamp 1701859473
transform 1 0 6730 0 -1 3390
box -12 -8 32 272
use FILL  FILL_2__1669_
timestamp 1701859473
transform -1 0 6770 0 -1 790
box -12 -8 32 272
use FILL  FILL_2__1670_
timestamp 1701859473
transform 1 0 6550 0 -1 2870
box -12 -8 32 272
use FILL  FILL_2__1671_
timestamp 1701859473
transform -1 0 6350 0 -1 8590
box -12 -8 32 272
use FILL  FILL_2__1672_
timestamp 1701859473
transform 1 0 5910 0 -1 10670
box -12 -8 32 272
use FILL  FILL_2__1673_
timestamp 1701859473
transform 1 0 6310 0 1 8590
box -12 -8 32 272
use FILL  FILL_2__1674_
timestamp 1701859473
transform -1 0 6390 0 -1 9110
box -12 -8 32 272
use FILL  FILL_2__1675_
timestamp 1701859473
transform 1 0 50 0 -1 5470
box -12 -8 32 272
use FILL  FILL_2__1676_
timestamp 1701859473
transform -1 0 290 0 -1 5470
box -12 -8 32 272
use FILL  FILL_2__1677_
timestamp 1701859473
transform -1 0 530 0 1 5470
box -12 -8 32 272
use FILL  FILL_2__1678_
timestamp 1701859473
transform 1 0 50 0 -1 10670
box -12 -8 32 272
use FILL  FILL_2__1679_
timestamp 1701859473
transform -1 0 270 0 -1 11190
box -12 -8 32 272
use FILL  FILL_2__1680_
timestamp 1701859473
transform 1 0 250 0 -1 10670
box -12 -8 32 272
use FILL  FILL_2__1681_
timestamp 1701859473
transform -1 0 70 0 -1 7030
box -12 -8 32 272
use FILL  FILL_2__1682_
timestamp 1701859473
transform -1 0 70 0 1 7030
box -12 -8 32 272
use FILL  FILL_2__1683_
timestamp 1701859473
transform 1 0 50 0 1 6510
box -12 -8 32 272
use FILL  FILL_2__1684_
timestamp 1701859473
transform 1 0 930 0 -1 11190
box -12 -8 32 272
use FILL  FILL_2__1685_
timestamp 1701859473
transform -1 0 1190 0 -1 11190
box -12 -8 32 272
use FILL  FILL_2__1686_
timestamp 1701859473
transform -1 0 990 0 1 10670
box -12 -8 32 272
use FILL  FILL_2__1687_
timestamp 1701859473
transform 1 0 1410 0 -1 11190
box -12 -8 32 272
use FILL  FILL_2__1688_
timestamp 1701859473
transform -1 0 1670 0 -1 11190
box -12 -8 32 272
use FILL  FILL_2__1689_
timestamp 1701859473
transform -1 0 1930 0 1 10150
box -12 -8 32 272
use FILL  FILL_2__1690_
timestamp 1701859473
transform 1 0 2090 0 1 9110
box -12 -8 32 272
use FILL  FILL_2__1691_
timestamp 1701859473
transform -1 0 2110 0 -1 9110
box -12 -8 32 272
use FILL  FILL_2__1692_
timestamp 1701859473
transform 1 0 50 0 1 790
box -12 -8 32 272
use FILL  FILL_2__1693_
timestamp 1701859473
transform 1 0 50 0 -1 1310
box -12 -8 32 272
use FILL  FILL_2__1694_
timestamp 1701859473
transform 1 0 470 0 -1 270
box -12 -8 32 272
use FILL  FILL_2__1695_
timestamp 1701859473
transform -1 0 690 0 -1 270
box -12 -8 32 272
use FILL  FILL_2__1696_
timestamp 1701859473
transform 1 0 1110 0 1 2870
box -12 -8 32 272
use FILL  FILL_2__1697_
timestamp 1701859473
transform -1 0 2770 0 -1 2870
box -12 -8 32 272
use FILL  FILL_2__1698_
timestamp 1701859473
transform -1 0 1870 0 1 3390
box -12 -8 32 272
use FILL  FILL_2__1699_
timestamp 1701859473
transform 1 0 3790 0 1 3390
box -12 -8 32 272
use FILL  FILL_2__1700_
timestamp 1701859473
transform -1 0 2590 0 -1 3910
box -12 -8 32 272
use FILL  FILL_2__1701_
timestamp 1701859473
transform -1 0 1130 0 1 270
box -12 -8 32 272
use FILL  FILL_2__1702_
timestamp 1701859473
transform 1 0 890 0 1 270
box -12 -8 32 272
use FILL  FILL_2__1703_
timestamp 1701859473
transform -1 0 1370 0 1 1830
box -12 -8 32 272
use FILL  FILL_2__1704_
timestamp 1701859473
transform -1 0 9130 0 1 2870
box -12 -8 32 272
use FILL  FILL_2__1705_
timestamp 1701859473
transform 1 0 9750 0 -1 790
box -12 -8 32 272
use FILL  FILL_2__1706_
timestamp 1701859473
transform -1 0 7970 0 -1 4950
box -12 -8 32 272
use FILL  FILL_2__1707_
timestamp 1701859473
transform 1 0 8410 0 -1 4950
box -12 -8 32 272
use FILL  FILL_2__1708_
timestamp 1701859473
transform 1 0 5030 0 -1 5990
box -12 -8 32 272
use FILL  FILL_2__1709_
timestamp 1701859473
transform -1 0 11130 0 1 5990
box -12 -8 32 272
use FILL  FILL_2__1710_
timestamp 1701859473
transform 1 0 5410 0 -1 5470
box -12 -8 32 272
use FILL  FILL_2__1711_
timestamp 1701859473
transform -1 0 5250 0 -1 5990
box -12 -8 32 272
use FILL  FILL_2__1712_
timestamp 1701859473
transform -1 0 5070 0 1 5470
box -12 -8 32 272
use FILL  FILL_2__1713_
timestamp 1701859473
transform 1 0 7930 0 1 4430
box -12 -8 32 272
use FILL  FILL_2__1714_
timestamp 1701859473
transform 1 0 7730 0 1 4950
box -12 -8 32 272
use FILL  FILL_2__1715_
timestamp 1701859473
transform -1 0 7970 0 1 4950
box -12 -8 32 272
use FILL  FILL_2__1716_
timestamp 1701859473
transform -1 0 8190 0 1 4430
box -12 -8 32 272
use FILL  FILL_2__1717_
timestamp 1701859473
transform -1 0 7970 0 1 1310
box -12 -8 32 272
use FILL  FILL_2__1718_
timestamp 1701859473
transform -1 0 5910 0 1 5990
box -12 -8 32 272
use FILL  FILL_2__1719_
timestamp 1701859473
transform -1 0 6770 0 -1 5990
box -12 -8 32 272
use FILL  FILL_2__1720_
timestamp 1701859473
transform -1 0 6750 0 1 5470
box -12 -8 32 272
use FILL  FILL_2__1721_
timestamp 1701859473
transform -1 0 6990 0 1 5470
box -12 -8 32 272
use FILL  FILL_2__1722_
timestamp 1701859473
transform -1 0 7690 0 1 4430
box -12 -8 32 272
use FILL  FILL_2__1723_
timestamp 1701859473
transform 1 0 7910 0 1 1830
box -12 -8 32 272
use FILL  FILL_2__1724_
timestamp 1701859473
transform -1 0 7950 0 -1 1310
box -12 -8 32 272
use FILL  FILL_2__1725_
timestamp 1701859473
transform 1 0 6550 0 1 5990
box -12 -8 32 272
use FILL  FILL_2__1726_
timestamp 1701859473
transform 1 0 6750 0 1 5990
box -12 -8 32 272
use FILL  FILL_2__1727_
timestamp 1701859473
transform -1 0 6990 0 1 5990
box -12 -8 32 272
use FILL  FILL_2__1728_
timestamp 1701859473
transform 1 0 7690 0 1 5990
box -12 -8 32 272
use FILL  FILL_2__1729_
timestamp 1701859473
transform -1 0 7630 0 -1 5990
box -12 -8 32 272
use FILL  FILL_2__1730_
timestamp 1701859473
transform -1 0 8110 0 1 3390
box -12 -8 32 272
use FILL  FILL_2__1731_
timestamp 1701859473
transform -1 0 7970 0 -1 270
box -12 -8 32 272
use FILL  FILL_2__1732_
timestamp 1701859473
transform -1 0 7930 0 1 5470
box -12 -8 32 272
use FILL  FILL_2__1733_
timestamp 1701859473
transform -1 0 8150 0 1 5470
box -12 -8 32 272
use FILL  FILL_2__1734_
timestamp 1701859473
transform 1 0 8110 0 -1 5470
box -12 -8 32 272
use FILL  FILL_2__1735_
timestamp 1701859473
transform 1 0 8570 0 -1 5470
box -12 -8 32 272
use FILL  FILL_2__1736_
timestamp 1701859473
transform 1 0 8410 0 1 4950
box -12 -8 32 272
use FILL  FILL_2__1737_
timestamp 1701859473
transform -1 0 8490 0 -1 3910
box -12 -8 32 272
use FILL  FILL_2__1738_
timestamp 1701859473
transform 1 0 8890 0 1 790
box -12 -8 32 272
use FILL  FILL_2__1739_
timestamp 1701859473
transform -1 0 9110 0 -1 790
box -12 -8 32 272
use FILL  FILL_2__1740_
timestamp 1701859473
transform 1 0 6470 0 1 270
box -12 -8 32 272
use FILL  FILL_2__1741_
timestamp 1701859473
transform 1 0 6370 0 1 790
box -12 -8 32 272
use FILL  FILL_2__1742_
timestamp 1701859473
transform -1 0 6310 0 -1 790
box -12 -8 32 272
use FILL  FILL_2__1743_
timestamp 1701859473
transform -1 0 2310 0 -1 3390
box -12 -8 32 272
use FILL  FILL_2__1744_
timestamp 1701859473
transform 1 0 290 0 -1 4950
box -12 -8 32 272
use FILL  FILL_2__1745_
timestamp 1701859473
transform 1 0 2110 0 -1 3910
box -12 -8 32 272
use FILL  FILL_2__1746_
timestamp 1701859473
transform -1 0 5130 0 -1 3390
box -12 -8 32 272
use FILL  FILL_2__1747_
timestamp 1701859473
transform -1 0 290 0 -1 270
box -12 -8 32 272
use FILL  FILL_2__1748_
timestamp 1701859473
transform -1 0 490 0 1 270
box -12 -8 32 272
use FILL  FILL_2__1749_
timestamp 1701859473
transform -1 0 930 0 1 1310
box -12 -8 32 272
use FILL  FILL_2__1750_
timestamp 1701859473
transform -1 0 1150 0 1 1310
box -12 -8 32 272
use FILL  FILL_2__1751_
timestamp 1701859473
transform -1 0 4510 0 -1 2870
box -12 -8 32 272
use FILL  FILL_2__1752_
timestamp 1701859473
transform 1 0 4710 0 -1 2870
box -12 -8 32 272
use FILL  FILL_2__1753_
timestamp 1701859473
transform -1 0 4330 0 1 790
box -12 -8 32 272
use FILL  FILL_2__1754_
timestamp 1701859473
transform 1 0 270 0 -1 790
box -12 -8 32 272
use FILL  FILL_2__1755_
timestamp 1701859473
transform -1 0 490 0 -1 790
box -12 -8 32 272
use FILL  FILL_2__1756_
timestamp 1701859473
transform -1 0 70 0 -1 270
box -12 -8 32 272
use FILL  FILL_2__1757_
timestamp 1701859473
transform 1 0 670 0 -1 790
box -12 -8 32 272
use FILL  FILL_2__1758_
timestamp 1701859473
transform 1 0 50 0 1 2350
box -12 -8 32 272
use FILL  FILL_2__1759_
timestamp 1701859473
transform -1 0 2550 0 -1 2870
box -12 -8 32 272
use FILL  FILL_2__1760_
timestamp 1701859473
transform 1 0 2930 0 -1 2870
box -12 -8 32 272
use FILL  FILL_2__1761_
timestamp 1701859473
transform -1 0 3250 0 -1 3390
box -12 -8 32 272
use FILL  FILL_2__1762_
timestamp 1701859473
transform -1 0 70 0 1 270
box -12 -8 32 272
use FILL  FILL_2__1763_
timestamp 1701859473
transform 1 0 50 0 -1 790
box -12 -8 32 272
use FILL  FILL_2__1764_
timestamp 1701859473
transform 1 0 490 0 1 1310
box -12 -8 32 272
use FILL  FILL_2__1765_
timestamp 1701859473
transform 1 0 1350 0 1 1310
box -12 -8 32 272
use FILL  FILL_2__1766_
timestamp 1701859473
transform -1 0 3150 0 -1 1830
box -12 -8 32 272
use FILL  FILL_2__1767_
timestamp 1701859473
transform 1 0 1450 0 -1 4430
box -12 -8 32 272
use FILL  FILL_2__1768_
timestamp 1701859473
transform 1 0 270 0 -1 1310
box -12 -8 32 272
use FILL  FILL_2__1769_
timestamp 1701859473
transform -1 0 490 0 1 1830
box -12 -8 32 272
use FILL  FILL_2__1770_
timestamp 1701859473
transform 1 0 2090 0 -1 3390
box -12 -8 32 272
use FILL  FILL_2__1771_
timestamp 1701859473
transform -1 0 2350 0 -1 3910
box -12 -8 32 272
use FILL  FILL_2__1772_
timestamp 1701859473
transform -1 0 3010 0 -1 3910
box -12 -8 32 272
use FILL  FILL_2__1773_
timestamp 1701859473
transform 1 0 3910 0 1 2870
box -12 -8 32 272
use FILL  FILL_2__1774_
timestamp 1701859473
transform -1 0 5290 0 -1 2350
box -12 -8 32 272
use FILL  FILL_2__1775_
timestamp 1701859473
transform 1 0 250 0 1 790
box -12 -8 32 272
use FILL  FILL_2__1776_
timestamp 1701859473
transform -1 0 290 0 1 1310
box -12 -8 32 272
use FILL  FILL_2__1777_
timestamp 1701859473
transform 1 0 710 0 -1 1830
box -12 -8 32 272
use FILL  FILL_2__1778_
timestamp 1701859473
transform -1 0 4430 0 1 5470
box -12 -8 32 272
use FILL  FILL_2__1779_
timestamp 1701859473
transform -1 0 6070 0 -1 5470
box -12 -8 32 272
use FILL  FILL_2__1780_
timestamp 1701859473
transform 1 0 4790 0 1 2870
box -12 -8 32 272
use FILL  FILL_2__1781_
timestamp 1701859473
transform 1 0 4370 0 1 2870
box -12 -8 32 272
use FILL  FILL_2__1782_
timestamp 1701859473
transform -1 0 70 0 1 1310
box -12 -8 32 272
use FILL  FILL_2__1783_
timestamp 1701859473
transform -1 0 1350 0 1 2870
box -12 -8 32 272
use FILL  FILL_2__1784_
timestamp 1701859473
transform -1 0 5050 0 1 2870
box -12 -8 32 272
use FILL  FILL_2__1785_
timestamp 1701859473
transform 1 0 4970 0 -1 2870
box -12 -8 32 272
use FILL  FILL_2__1786_
timestamp 1701859473
transform -1 0 5050 0 -1 2350
box -12 -8 32 272
use FILL  FILL_2__1787_
timestamp 1701859473
transform 1 0 5030 0 1 2350
box -12 -8 32 272
use FILL  FILL_2__1788_
timestamp 1701859473
transform -1 0 4830 0 -1 2350
box -12 -8 32 272
use FILL  FILL_2__1789_
timestamp 1701859473
transform 1 0 50 0 1 1830
box -12 -8 32 272
use FILL  FILL_2__1790_
timestamp 1701859473
transform -1 0 290 0 -1 2350
box -12 -8 32 272
use FILL  FILL_2__1791_
timestamp 1701859473
transform -1 0 2090 0 -1 2350
box -12 -8 32 272
use FILL  FILL_2__1792_
timestamp 1701859473
transform -1 0 3470 0 -1 2350
box -12 -8 32 272
use FILL  FILL_2__1793_
timestamp 1701859473
transform -1 0 4570 0 1 1830
box -12 -8 32 272
use FILL  FILL_2__1794_
timestamp 1701859473
transform 1 0 890 0 1 1830
box -12 -8 32 272
use FILL  FILL_2__1795_
timestamp 1701859473
transform -1 0 2150 0 1 2350
box -12 -8 32 272
use FILL  FILL_2__1796_
timestamp 1701859473
transform -1 0 1770 0 -1 1830
box -12 -8 32 272
use FILL  FILL_2__1797_
timestamp 1701859473
transform 1 0 1990 0 -1 1830
box -12 -8 32 272
use FILL  FILL_2__1798_
timestamp 1701859473
transform 1 0 910 0 -1 1310
box -12 -8 32 272
use FILL  FILL_2__1799_
timestamp 1701859473
transform 1 0 3730 0 1 3910
box -12 -8 32 272
use FILL  FILL_2__1800_
timestamp 1701859473
transform 1 0 3410 0 1 1830
box -12 -8 32 272
use FILL  FILL_2__1801_
timestamp 1701859473
transform -1 0 1150 0 1 1830
box -12 -8 32 272
use FILL  FILL_2__1802_
timestamp 1701859473
transform -1 0 3690 0 1 2350
box -12 -8 32 272
use FILL  FILL_2__1803_
timestamp 1701859473
transform -1 0 3910 0 1 2350
box -12 -8 32 272
use FILL  FILL_2__1804_
timestamp 1701859473
transform -1 0 4150 0 1 2350
box -12 -8 32 272
use FILL  FILL_2__1805_
timestamp 1701859473
transform 1 0 5450 0 1 2350
box -12 -8 32 272
use FILL  FILL_2__1806_
timestamp 1701859473
transform -1 0 4850 0 1 2350
box -12 -8 32 272
use FILL  FILL_2__1807_
timestamp 1701859473
transform -1 0 5250 0 1 2350
box -12 -8 32 272
use FILL  FILL_2__1808_
timestamp 1701859473
transform 1 0 4770 0 1 1830
box -12 -8 32 272
use FILL  FILL_2__1809_
timestamp 1701859473
transform -1 0 7130 0 -1 270
box -12 -8 32 272
use FILL  FILL_2__1810_
timestamp 1701859473
transform -1 0 7110 0 1 1310
box -12 -8 32 272
use FILL  FILL_2__1811_
timestamp 1701859473
transform 1 0 7450 0 -1 1830
box -12 -8 32 272
use FILL  FILL_2__1812_
timestamp 1701859473
transform -1 0 7530 0 -1 1310
box -12 -8 32 272
use FILL  FILL_2__1813_
timestamp 1701859473
transform 1 0 9110 0 1 790
box -12 -8 32 272
use FILL  FILL_2__1814_
timestamp 1701859473
transform -1 0 8150 0 -1 1830
box -12 -8 32 272
use FILL  FILL_2__1815_
timestamp 1701859473
transform 1 0 8350 0 1 2350
box -12 -8 32 272
use FILL  FILL_2__1816_
timestamp 1701859473
transform -1 0 9630 0 -1 2350
box -12 -8 32 272
use FILL  FILL_2__1817_
timestamp 1701859473
transform -1 0 9350 0 1 1310
box -12 -8 32 272
use FILL  FILL_2__1818_
timestamp 1701859473
transform -1 0 9550 0 1 270
box -12 -8 32 272
use FILL  FILL_2__1819_
timestamp 1701859473
transform -1 0 8370 0 -1 1830
box -12 -8 32 272
use FILL  FILL_2__1820_
timestamp 1701859473
transform -1 0 8450 0 1 1310
box -12 -8 32 272
use FILL  FILL_2__1821_
timestamp 1701859473
transform -1 0 4890 0 1 1310
box -12 -8 32 272
use FILL  FILL_2__1822_
timestamp 1701859473
transform -1 0 4690 0 -1 790
box -12 -8 32 272
use FILL  FILL_2__1823_
timestamp 1701859473
transform -1 0 4230 0 -1 790
box -12 -8 32 272
use FILL  FILL_2__1824_
timestamp 1701859473
transform 1 0 4610 0 1 2350
box -12 -8 32 272
use FILL  FILL_2__1825_
timestamp 1701859473
transform 1 0 5670 0 1 1830
box -12 -8 32 272
use FILL  FILL_2__1826_
timestamp 1701859473
transform 1 0 8170 0 -1 270
box -12 -8 32 272
use FILL  FILL_2__1827_
timestamp 1701859473
transform 1 0 9310 0 -1 790
box -12 -8 32 272
use FILL  FILL_2__1828_
timestamp 1701859473
transform 1 0 8470 0 1 270
box -12 -8 32 272
use FILL  FILL_2__1829_
timestamp 1701859473
transform 1 0 5770 0 1 270
box -12 -8 32 272
use FILL  FILL_2__1830_
timestamp 1701859473
transform 1 0 3210 0 1 4430
box -12 -8 32 272
use FILL  FILL_2__1831_
timestamp 1701859473
transform -1 0 7990 0 -1 790
box -12 -8 32 272
use FILL  FILL_2__1832_
timestamp 1701859473
transform 1 0 6490 0 -1 790
box -12 -8 32 272
use FILL  FILL_2__1833_
timestamp 1701859473
transform -1 0 690 0 1 270
box -12 -8 32 272
use FILL  FILL_2__1834_
timestamp 1701859473
transform 1 0 1130 0 -1 1310
box -12 -8 32 272
use FILL  FILL_2__1835_
timestamp 1701859473
transform -1 0 2510 0 -1 1310
box -12 -8 32 272
use FILL  FILL_2__1836_
timestamp 1701859473
transform 1 0 1070 0 1 790
box -12 -8 32 272
use FILL  FILL_2__1837_
timestamp 1701859473
transform -1 0 2470 0 1 790
box -12 -8 32 272
use FILL  FILL_2__1838_
timestamp 1701859473
transform 1 0 2210 0 1 790
box -12 -8 32 272
use FILL  FILL_2__1839_
timestamp 1701859473
transform -1 0 270 0 1 270
box -12 -8 32 272
use FILL  FILL_2__1840_
timestamp 1701859473
transform -1 0 910 0 1 2870
box -12 -8 32 272
use FILL  FILL_2__1841_
timestamp 1701859473
transform 1 0 3690 0 1 2870
box -12 -8 32 272
use FILL  FILL_2__1842_
timestamp 1701859473
transform -1 0 2950 0 -1 1830
box -12 -8 32 272
use FILL  FILL_2__1843_
timestamp 1701859473
transform -1 0 3910 0 -1 2350
box -12 -8 32 272
use FILL  FILL_2__1844_
timestamp 1701859473
transform 1 0 3810 0 -1 2870
box -12 -8 32 272
use FILL  FILL_2__1845_
timestamp 1701859473
transform -1 0 1750 0 -1 4950
box -12 -8 32 272
use FILL  FILL_2__1846_
timestamp 1701859473
transform 1 0 4110 0 1 4430
box -12 -8 32 272
use FILL  FILL_2__1847_
timestamp 1701859473
transform 1 0 3430 0 1 4430
box -12 -8 32 272
use FILL  FILL_2__1848_
timestamp 1701859473
transform 1 0 3870 0 1 4430
box -12 -8 32 272
use FILL  FILL_2__1849_
timestamp 1701859473
transform -1 0 4070 0 -1 2870
box -12 -8 32 272
use FILL  FILL_2__1850_
timestamp 1701859473
transform -1 0 890 0 1 790
box -12 -8 32 272
use FILL  FILL_2__1851_
timestamp 1701859473
transform 1 0 1550 0 -1 1830
box -12 -8 32 272
use FILL  FILL_2__1852_
timestamp 1701859473
transform -1 0 2370 0 1 2350
box -12 -8 32 272
use FILL  FILL_2__1853_
timestamp 1701859473
transform 1 0 50 0 -1 2350
box -12 -8 32 272
use FILL  FILL_2__1854_
timestamp 1701859473
transform 1 0 2290 0 -1 2350
box -12 -8 32 272
use FILL  FILL_2__1855_
timestamp 1701859473
transform -1 0 2550 0 -1 2350
box -12 -8 32 272
use FILL  FILL_2__1856_
timestamp 1701859473
transform 1 0 1450 0 -1 790
box -12 -8 32 272
use FILL  FILL_2__1857_
timestamp 1701859473
transform -1 0 2650 0 -1 790
box -12 -8 32 272
use FILL  FILL_2__1858_
timestamp 1701859473
transform 1 0 2390 0 -1 790
box -12 -8 32 272
use FILL  FILL_2__1859_
timestamp 1701859473
transform 1 0 2170 0 -1 790
box -12 -8 32 272
use FILL  FILL_2__1860_
timestamp 1701859473
transform -1 0 1710 0 -1 790
box -12 -8 32 272
use FILL  FILL_2__1861_
timestamp 1701859473
transform -1 0 1950 0 -1 790
box -12 -8 32 272
use FILL  FILL_2__1862_
timestamp 1701859473
transform -1 0 2030 0 1 270
box -12 -8 32 272
use FILL  FILL_2__1863_
timestamp 1701859473
transform 1 0 2250 0 1 270
box -12 -8 32 272
use FILL  FILL_2__1864_
timestamp 1701859473
transform 1 0 3490 0 1 270
box -12 -8 32 272
use FILL  FILL_2__1865_
timestamp 1701859473
transform 1 0 7290 0 -1 1310
box -12 -8 32 272
use FILL  FILL_2__1866_
timestamp 1701859473
transform 1 0 3650 0 -1 1310
box -12 -8 32 272
use FILL  FILL_2__1867_
timestamp 1701859473
transform 1 0 1110 0 -1 1830
box -12 -8 32 272
use FILL  FILL_2__1868_
timestamp 1701859473
transform 1 0 1550 0 1 1310
box -12 -8 32 272
use FILL  FILL_2__1869_
timestamp 1701859473
transform 1 0 1970 0 1 1310
box -12 -8 32 272
use FILL  FILL_2__1870_
timestamp 1701859473
transform -1 0 1590 0 -1 1310
box -12 -8 32 272
use FILL  FILL_2__1871_
timestamp 1701859473
transform -1 0 2710 0 -1 1310
box -12 -8 32 272
use FILL  FILL_2__1872_
timestamp 1701859473
transform -1 0 490 0 1 790
box -12 -8 32 272
use FILL  FILL_2__1873_
timestamp 1701859473
transform 1 0 670 0 1 790
box -12 -8 32 272
use FILL  FILL_2__1874_
timestamp 1701859473
transform -1 0 1310 0 1 790
box -12 -8 32 272
use FILL  FILL_2__1875_
timestamp 1701859473
transform 1 0 890 0 -1 790
box -12 -8 32 272
use FILL  FILL_2__1876_
timestamp 1701859473
transform 1 0 1210 0 -1 790
box -12 -8 32 272
use FILL  FILL_2__1877_
timestamp 1701859473
transform 1 0 2150 0 1 4950
box -12 -8 32 272
use FILL  FILL_2__1878_
timestamp 1701859473
transform 1 0 490 0 -1 1310
box -12 -8 32 272
use FILL  FILL_2__1879_
timestamp 1701859473
transform 1 0 710 0 1 1310
box -12 -8 32 272
use FILL  FILL_2__1880_
timestamp 1701859473
transform -1 0 1970 0 -1 4950
box -12 -8 32 272
use FILL  FILL_2__1881_
timestamp 1701859473
transform -1 0 2210 0 -1 4950
box -12 -8 32 272
use FILL  FILL_2__1882_
timestamp 1701859473
transform 1 0 1530 0 -1 3390
box -12 -8 32 272
use FILL  FILL_2__1883_
timestamp 1701859473
transform 1 0 1010 0 -1 3390
box -12 -8 32 272
use FILL  FILL_2__1884_
timestamp 1701859473
transform -1 0 4030 0 1 3390
box -12 -8 32 272
use FILL  FILL_2__1885_
timestamp 1701859473
transform -1 0 3750 0 -1 3390
box -12 -8 32 272
use FILL  FILL_2__1886_
timestamp 1701859473
transform 1 0 3490 0 -1 3390
box -12 -8 32 272
use FILL  FILL_2__1887_
timestamp 1701859473
transform -1 0 3470 0 1 2870
box -12 -8 32 272
use FILL  FILL_2__1888_
timestamp 1701859473
transform -1 0 2510 0 1 270
box -12 -8 32 272
use FILL  FILL_2__1889_
timestamp 1701859473
transform 1 0 1650 0 -1 2870
box -12 -8 32 272
use FILL  FILL_2__1890_
timestamp 1701859473
transform -1 0 290 0 -1 1830
box -12 -8 32 272
use FILL  FILL_2__1891_
timestamp 1701859473
transform 1 0 50 0 -1 1830
box -12 -8 32 272
use FILL  FILL_2__1892_
timestamp 1701859473
transform 1 0 4890 0 -1 3390
box -12 -8 32 272
use FILL  FILL_2__1893_
timestamp 1701859473
transform 1 0 3890 0 1 1830
box -12 -8 32 272
use FILL  FILL_2__1894_
timestamp 1701859473
transform 1 0 4090 0 1 1830
box -12 -8 32 272
use FILL  FILL_2__1895_
timestamp 1701859473
transform -1 0 1830 0 1 1830
box -12 -8 32 272
use FILL  FILL_2__1896_
timestamp 1701859473
transform 1 0 1850 0 -1 2350
box -12 -8 32 272
use FILL  FILL_2__1897_
timestamp 1701859473
transform 1 0 3470 0 1 2350
box -12 -8 32 272
use FILL  FILL_2__1898_
timestamp 1701859473
transform 1 0 3250 0 1 2350
box -12 -8 32 272
use FILL  FILL_2__1899_
timestamp 1701859473
transform -1 0 3230 0 -1 2350
box -12 -8 32 272
use FILL  FILL_2__1900_
timestamp 1701859473
transform -1 0 4070 0 -1 1830
box -12 -8 32 272
use FILL  FILL_2__1901_
timestamp 1701859473
transform -1 0 710 0 1 1830
box -12 -8 32 272
use FILL  FILL_2__1902_
timestamp 1701859473
transform 1 0 5010 0 1 1830
box -12 -8 32 272
use FILL  FILL_2__1903_
timestamp 1701859473
transform 1 0 3330 0 1 1310
box -12 -8 32 272
use FILL  FILL_2__1904_
timestamp 1701859473
transform -1 0 3430 0 -1 1310
box -12 -8 32 272
use FILL  FILL_2__1905_
timestamp 1701859473
transform 1 0 2970 0 1 270
box -12 -8 32 272
use FILL  FILL_2__1906_
timestamp 1701859473
transform 1 0 250 0 1 2350
box -12 -8 32 272
use FILL  FILL_2__1907_
timestamp 1701859473
transform -1 0 3010 0 -1 2350
box -12 -8 32 272
use FILL  FILL_2__1908_
timestamp 1701859473
transform 1 0 6430 0 -1 2350
box -12 -8 32 272
use FILL  FILL_2__1909_
timestamp 1701859473
transform -1 0 6030 0 -1 2350
box -12 -8 32 272
use FILL  FILL_2__1910_
timestamp 1701859473
transform -1 0 5530 0 -1 2350
box -12 -8 32 272
use FILL  FILL_2__1911_
timestamp 1701859473
transform -1 0 690 0 1 2870
box -12 -8 32 272
use FILL  FILL_2__1912_
timestamp 1701859473
transform -1 0 3290 0 1 3910
box -12 -8 32 272
use FILL  FILL_2__1913_
timestamp 1701859473
transform -1 0 1010 0 -1 2870
box -12 -8 32 272
use FILL  FILL_2__1914_
timestamp 1701859473
transform -1 0 1450 0 1 3390
box -12 -8 32 272
use FILL  FILL_2__1915_
timestamp 1701859473
transform 1 0 2530 0 1 3390
box -12 -8 32 272
use FILL  FILL_2__1916_
timestamp 1701859473
transform -1 0 3390 0 1 3390
box -12 -8 32 272
use FILL  FILL_2__1917_
timestamp 1701859473
transform -1 0 4670 0 -1 3390
box -12 -8 32 272
use FILL  FILL_2__1918_
timestamp 1701859473
transform 1 0 1710 0 1 4950
box -12 -8 32 272
use FILL  FILL_2__1919_
timestamp 1701859473
transform -1 0 1230 0 -1 2870
box -12 -8 32 272
use FILL  FILL_2__1920_
timestamp 1701859473
transform -1 0 5010 0 1 4430
box -12 -8 32 272
use FILL  FILL_2__1921_
timestamp 1701859473
transform 1 0 4770 0 1 4430
box -12 -8 32 272
use FILL  FILL_2__1922_
timestamp 1701859473
transform -1 0 4570 0 1 4430
box -12 -8 32 272
use FILL  FILL_2__1923_
timestamp 1701859473
transform 1 0 4430 0 -1 3390
box -12 -8 32 272
use FILL  FILL_2__1924_
timestamp 1701859473
transform 1 0 1930 0 1 4950
box -12 -8 32 272
use FILL  FILL_2__1925_
timestamp 1701859473
transform 1 0 6070 0 -1 4430
box -12 -8 32 272
use FILL  FILL_2__1926_
timestamp 1701859473
transform 1 0 690 0 -1 1310
box -12 -8 32 272
use FILL  FILL_2__1927_
timestamp 1701859473
transform 1 0 2930 0 -1 1310
box -12 -8 32 272
use FILL  FILL_2__1928_
timestamp 1701859473
transform -1 0 3190 0 -1 1310
box -12 -8 32 272
use FILL  FILL_2__1929_
timestamp 1701859473
transform 1 0 3370 0 1 790
box -12 -8 32 272
use FILL  FILL_2__1930_
timestamp 1701859473
transform 1 0 3190 0 1 270
box -12 -8 32 272
use FILL  FILL_2__1931_
timestamp 1701859473
transform 1 0 3790 0 1 270
box -12 -8 32 272
use FILL  FILL_2__1932_
timestamp 1701859473
transform -1 0 4030 0 1 270
box -12 -8 32 272
use FILL  FILL_2__1933_
timestamp 1701859473
transform -1 0 1830 0 1 270
box -12 -8 32 272
use FILL  FILL_2__1934_
timestamp 1701859473
transform -1 0 5450 0 1 790
box -12 -8 32 272
use FILL  FILL_2__1935_
timestamp 1701859473
transform 1 0 5570 0 -1 270
box -12 -8 32 272
use FILL  FILL_2__1936_
timestamp 1701859473
transform -1 0 8330 0 1 3390
box -12 -8 32 272
use FILL  FILL_2__1937_
timestamp 1701859473
transform -1 0 7550 0 -1 270
box -12 -8 32 272
use FILL  FILL_2__1938_
timestamp 1701859473
transform -1 0 7750 0 -1 270
box -12 -8 32 272
use FILL  FILL_2__1939_
timestamp 1701859473
transform -1 0 6670 0 -1 270
box -12 -8 32 272
use FILL  FILL_2__1940_
timestamp 1701859473
transform -1 0 5790 0 -1 270
box -12 -8 32 272
use FILL  FILL_2__1941_
timestamp 1701859473
transform 1 0 5810 0 -1 790
box -12 -8 32 272
use FILL  FILL_2__1942_
timestamp 1701859473
transform 1 0 4790 0 -1 1310
box -12 -8 32 272
use FILL  FILL_2__1943_
timestamp 1701859473
transform 1 0 8050 0 1 270
box -12 -8 32 272
use FILL  FILL_2__1944_
timestamp 1701859473
transform -1 0 8290 0 1 270
box -12 -8 32 272
use FILL  FILL_2__1945_
timestamp 1701859473
transform 1 0 7830 0 1 270
box -12 -8 32 272
use FILL  FILL_2__1946_
timestamp 1701859473
transform -1 0 6030 0 1 270
box -12 -8 32 272
use FILL  FILL_2__1947_
timestamp 1701859473
transform -1 0 6050 0 -1 790
box -12 -8 32 272
use FILL  FILL_2__1948_
timestamp 1701859473
transform 1 0 5330 0 -1 790
box -12 -8 32 272
use FILL  FILL_2__1949_
timestamp 1701859473
transform 1 0 4570 0 -1 1310
box -12 -8 32 272
use FILL  FILL_2__1950_
timestamp 1701859473
transform -1 0 8210 0 -1 790
box -12 -8 32 272
use FILL  FILL_2__1951_
timestamp 1701859473
transform 1 0 490 0 -1 2350
box -12 -8 32 272
use FILL  FILL_2__1952_
timestamp 1701859473
transform -1 0 5670 0 1 2350
box -12 -8 32 272
use FILL  FILL_2__1953_
timestamp 1701859473
transform 1 0 5770 0 -1 2350
box -12 -8 32 272
use FILL  FILL_2__1954_
timestamp 1701859473
transform 1 0 8150 0 -1 1310
box -12 -8 32 272
use FILL  FILL_2__1955_
timestamp 1701859473
transform -1 0 8690 0 1 1310
box -12 -8 32 272
use FILL  FILL_2__1956_
timestamp 1701859473
transform -1 0 6230 0 -1 1310
box -12 -8 32 272
use FILL  FILL_2__1957_
timestamp 1701859473
transform -1 0 5990 0 -1 1310
box -12 -8 32 272
use FILL  FILL_2__1958_
timestamp 1701859473
transform 1 0 5250 0 -1 1310
box -12 -8 32 272
use FILL  FILL_2__1959_
timestamp 1701859473
transform 1 0 5690 0 -1 2870
box -12 -8 32 272
use FILL  FILL_2__1960_
timestamp 1701859473
transform -1 0 6130 0 -1 2870
box -12 -8 32 272
use FILL  FILL_2__1961_
timestamp 1701859473
transform -1 0 4390 0 1 2350
box -12 -8 32 272
use FILL  FILL_2__1962_
timestamp 1701859473
transform 1 0 5850 0 1 2350
box -12 -8 32 272
use FILL  FILL_2__1963_
timestamp 1701859473
transform 1 0 5310 0 1 1310
box -12 -8 32 272
use FILL  FILL_2__1964_
timestamp 1701859473
transform 1 0 9130 0 1 1310
box -12 -8 32 272
use FILL  FILL_2__1965_
timestamp 1701859473
transform 1 0 7530 0 1 790
box -12 -8 32 272
use FILL  FILL_2__1966_
timestamp 1701859473
transform -1 0 7650 0 1 270
box -12 -8 32 272
use FILL  FILL_2__1967_
timestamp 1701859473
transform -1 0 6710 0 1 270
box -12 -8 32 272
use FILL  FILL_2__1968_
timestamp 1701859473
transform 1 0 5490 0 -1 1310
box -12 -8 32 272
use FILL  FILL_2__1969_
timestamp 1701859473
transform 1 0 5690 0 1 2870
box -12 -8 32 272
use FILL  FILL_2__1970_
timestamp 1701859473
transform 1 0 5330 0 -1 3390
box -12 -8 32 272
use FILL  FILL_2__1971_
timestamp 1701859473
transform 1 0 5770 0 1 3910
box -12 -8 32 272
use FILL  FILL_2__1972_
timestamp 1701859473
transform 1 0 5710 0 1 4950
box -12 -8 32 272
use FILL  FILL_2__1973_
timestamp 1701859473
transform -1 0 6050 0 -1 3910
box -12 -8 32 272
use FILL  FILL_2__1974_
timestamp 1701859473
transform 1 0 6230 0 -1 3910
box -12 -8 32 272
use FILL  FILL_2__1975_
timestamp 1701859473
transform -1 0 6030 0 1 3910
box -12 -8 32 272
use FILL  FILL_2__1976_
timestamp 1701859473
transform -1 0 6490 0 -1 3910
box -12 -8 32 272
use FILL  FILL_2__1977_
timestamp 1701859473
transform 1 0 6810 0 1 2870
box -12 -8 32 272
use FILL  FILL_2__1978_
timestamp 1701859473
transform -1 0 6350 0 -1 2870
box -12 -8 32 272
use FILL  FILL_2__1979_
timestamp 1701859473
transform 1 0 6390 0 1 2870
box -12 -8 32 272
use FILL  FILL_2__1980_
timestamp 1701859473
transform 1 0 6590 0 1 2870
box -12 -8 32 272
use FILL  FILL_2__1981_
timestamp 1701859473
transform 1 0 6170 0 1 2870
box -12 -8 32 272
use FILL  FILL_2__1982_
timestamp 1701859473
transform -1 0 5630 0 -1 1830
box -12 -8 32 272
use FILL  FILL_2__1983_
timestamp 1701859473
transform -1 0 4730 0 -1 270
box -12 -8 32 272
use FILL  FILL_2__1984_
timestamp 1701859473
transform -1 0 6430 0 -1 1310
box -12 -8 32 272
use FILL  FILL_2__1985_
timestamp 1701859473
transform 1 0 4990 0 -1 1310
box -12 -8 32 272
use FILL  FILL_2__1986_
timestamp 1701859473
transform 1 0 8190 0 1 790
box -12 -8 32 272
use FILL  FILL_2__1987_
timestamp 1701859473
transform 1 0 6870 0 1 1310
box -12 -8 32 272
use FILL  FILL_2__1988_
timestamp 1701859473
transform -1 0 7330 0 1 1310
box -12 -8 32 272
use FILL  FILL_2__1989_
timestamp 1701859473
transform 1 0 2690 0 -1 5470
box -12 -8 32 272
use FILL  FILL_2__1990_
timestamp 1701859473
transform 1 0 2010 0 1 1830
box -12 -8 32 272
use FILL  FILL_2__1991_
timestamp 1701859473
transform -1 0 2730 0 1 1830
box -12 -8 32 272
use FILL  FILL_2__1992_
timestamp 1701859473
transform -1 0 4130 0 -1 2350
box -12 -8 32 272
use FILL  FILL_2__1993_
timestamp 1701859473
transform -1 0 4370 0 -1 2350
box -12 -8 32 272
use FILL  FILL_2__1994_
timestamp 1701859473
transform 1 0 2470 0 1 1830
box -12 -8 32 272
use FILL  FILL_2__1995_
timestamp 1701859473
transform 1 0 2950 0 1 1830
box -12 -8 32 272
use FILL  FILL_2__1996_
timestamp 1701859473
transform -1 0 6630 0 1 790
box -12 -8 32 272
use FILL  FILL_2__1997_
timestamp 1701859473
transform -1 0 4970 0 1 790
box -12 -8 32 272
use FILL  FILL_2__1998_
timestamp 1701859473
transform 1 0 4230 0 1 270
box -12 -8 32 272
use FILL  FILL_2__1999_
timestamp 1701859473
transform -1 0 3830 0 -1 270
box -12 -8 32 272
use FILL  FILL_2__2000_
timestamp 1701859473
transform -1 0 4510 0 -1 270
box -12 -8 32 272
use FILL  FILL_2__2001_
timestamp 1701859473
transform -1 0 5890 0 -1 2870
box -12 -8 32 272
use FILL  FILL_2__2002_
timestamp 1701859473
transform -1 0 1830 0 1 2870
box -12 -8 32 272
use FILL  FILL_2__2003_
timestamp 1701859473
transform 1 0 1330 0 -1 3390
box -12 -8 32 272
use FILL  FILL_2__2004_
timestamp 1701859473
transform 1 0 2750 0 -1 3390
box -12 -8 32 272
use FILL  FILL_2__2005_
timestamp 1701859473
transform -1 0 3030 0 1 2870
box -12 -8 32 272
use FILL  FILL_2__2006_
timestamp 1701859473
transform 1 0 2770 0 1 2870
box -12 -8 32 272
use FILL  FILL_2__2007_
timestamp 1701859473
transform 1 0 6790 0 -1 2870
box -12 -8 32 272
use FILL  FILL_2__2008_
timestamp 1701859473
transform 1 0 470 0 -1 1830
box -12 -8 32 272
use FILL  FILL_2__2009_
timestamp 1701859473
transform -1 0 3990 0 -1 3390
box -12 -8 32 272
use FILL  FILL_2__2010_
timestamp 1701859473
transform -1 0 4290 0 -1 2870
box -12 -8 32 272
use FILL  FILL_2__2011_
timestamp 1701859473
transform -1 0 2030 0 1 790
box -12 -8 32 272
use FILL  FILL_2__2012_
timestamp 1701859473
transform 1 0 1530 0 1 790
box -12 -8 32 272
use FILL  FILL_2__2013_
timestamp 1701859473
transform -1 0 1790 0 1 790
box -12 -8 32 272
use FILL  FILL_2__2014_
timestamp 1701859473
transform 1 0 4450 0 1 1310
box -12 -8 32 272
use FILL  FILL_2__2015_
timestamp 1701859473
transform 1 0 3170 0 1 1830
box -12 -8 32 272
use FILL  FILL_2__2016_
timestamp 1701859473
transform -1 0 3670 0 1 1830
box -12 -8 32 272
use FILL  FILL_2__2017_
timestamp 1701859473
transform -1 0 5190 0 -1 1830
box -12 -8 32 272
use FILL  FILL_2__2018_
timestamp 1701859473
transform 1 0 4950 0 -1 1830
box -12 -8 32 272
use FILL  FILL_2__2019_
timestamp 1701859473
transform -1 0 5470 0 -1 2870
box -12 -8 32 272
use FILL  FILL_2__2020_
timestamp 1701859473
transform -1 0 5230 0 -1 2870
box -12 -8 32 272
use FILL  FILL_2__2021_
timestamp 1701859473
transform -1 0 6870 0 -1 1310
box -12 -8 32 272
use FILL  FILL_2__2022_
timestamp 1701859473
transform -1 0 7110 0 1 790
box -12 -8 32 272
use FILL  FILL_2__2023_
timestamp 1701859473
transform 1 0 8150 0 1 1830
box -12 -8 32 272
use FILL  FILL_2__2024_
timestamp 1701859473
transform -1 0 8370 0 1 1830
box -12 -8 32 272
use FILL  FILL_2__2025_
timestamp 1701859473
transform 1 0 9530 0 -1 790
box -12 -8 32 272
use FILL  FILL_2__2026_
timestamp 1701859473
transform -1 0 8670 0 1 790
box -12 -8 32 272
use FILL  FILL_2__2027_
timestamp 1701859473
transform -1 0 6870 0 1 790
box -12 -8 32 272
use FILL  FILL_2__2028_
timestamp 1701859473
transform 1 0 6970 0 -1 790
box -12 -8 32 272
use FILL  FILL_2__2029_
timestamp 1701859473
transform 1 0 7410 0 1 270
box -12 -8 32 272
use FILL  FILL_2__2030_
timestamp 1701859473
transform -1 0 7090 0 -1 1310
box -12 -8 32 272
use FILL  FILL_2__2031_
timestamp 1701859473
transform 1 0 7410 0 -1 790
box -12 -8 32 272
use FILL  FILL_2__2032_
timestamp 1701859473
transform -1 0 8710 0 1 270
box -12 -8 32 272
use FILL  FILL_2__2033_
timestamp 1701859473
transform 1 0 8190 0 1 1310
box -12 -8 32 272
use FILL  FILL_2__2034_
timestamp 1701859473
transform -1 0 8870 0 -1 1310
box -12 -8 32 272
use FILL  FILL_2__2035_
timestamp 1701859473
transform -1 0 8450 0 1 790
box -12 -8 32 272
use FILL  FILL_2__2036_
timestamp 1701859473
transform -1 0 8610 0 -1 1830
box -12 -8 32 272
use FILL  FILL_2__2037_
timestamp 1701859473
transform -1 0 8670 0 -1 790
box -12 -8 32 272
use FILL  FILL_2__2038_
timestamp 1701859473
transform 1 0 7970 0 1 790
box -12 -8 32 272
use FILL  FILL_2__2039_
timestamp 1701859473
transform 1 0 7750 0 1 790
box -12 -8 32 272
use FILL  FILL_2__2040_
timestamp 1701859473
transform -1 0 7670 0 -1 790
box -12 -8 32 272
use FILL  FILL_2__2041_
timestamp 1701859473
transform -1 0 6890 0 -1 270
box -12 -8 32 272
use FILL  FILL_2__2042_
timestamp 1701859473
transform 1 0 8870 0 -1 790
box -12 -8 32 272
use FILL  FILL_2__2043_
timestamp 1701859473
transform 1 0 7190 0 1 270
box -12 -8 32 272
use FILL  FILL_2__2044_
timestamp 1701859473
transform 1 0 6930 0 1 270
box -12 -8 32 272
use FILL  FILL_2__2045_
timestamp 1701859473
transform -1 0 6250 0 1 270
box -12 -8 32 272
use FILL  FILL_2__2046_
timestamp 1701859473
transform 1 0 6430 0 -1 270
box -12 -8 32 272
use FILL  FILL_2__2047_
timestamp 1701859473
transform -1 0 6210 0 -1 270
box -12 -8 32 272
use FILL  FILL_2__2048_
timestamp 1701859473
transform -1 0 6010 0 -1 270
box -12 -8 32 272
use FILL  FILL_2__2049_
timestamp 1701859473
transform -1 0 7190 0 -1 790
box -12 -8 32 272
use FILL  FILL_2__2050_
timestamp 1701859473
transform 1 0 1430 0 -1 2870
box -12 -8 32 272
use FILL  FILL_2__2051_
timestamp 1701859473
transform 1 0 6230 0 -1 2350
box -12 -8 32 272
use FILL  FILL_2__2052_
timestamp 1701859473
transform -1 0 6130 0 1 790
box -12 -8 32 272
use FILL  FILL_2__2053_
timestamp 1701859473
transform -1 0 4350 0 1 1830
box -12 -8 32 272
use FILL  FILL_2__2054_
timestamp 1701859473
transform 1 0 2850 0 1 1310
box -12 -8 32 272
use FILL  FILL_2__2055_
timestamp 1701859473
transform -1 0 3110 0 1 1310
box -12 -8 32 272
use FILL  FILL_2__2056_
timestamp 1701859473
transform -1 0 1830 0 -1 1310
box -12 -8 32 272
use FILL  FILL_2__2057_
timestamp 1701859473
transform 1 0 2690 0 1 790
box -12 -8 32 272
use FILL  FILL_2__2058_
timestamp 1701859473
transform 1 0 3610 0 1 790
box -12 -8 32 272
use FILL  FILL_2__2059_
timestamp 1701859473
transform 1 0 3850 0 1 790
box -12 -8 32 272
use FILL  FILL_2__2060_
timestamp 1701859473
transform -1 0 4090 0 1 790
box -12 -8 32 272
use FILL  FILL_2__2061_
timestamp 1701859473
transform -1 0 2950 0 -1 270
box -12 -8 32 272
use FILL  FILL_2__2062_
timestamp 1701859473
transform 1 0 2730 0 1 270
box -12 -8 32 272
use FILL  FILL_2__2063_
timestamp 1701859473
transform 1 0 3110 0 -1 270
box -12 -8 32 272
use FILL  FILL_2__2064_
timestamp 1701859473
transform 1 0 3350 0 -1 270
box -12 -8 32 272
use FILL  FILL_2__2065_
timestamp 1701859473
transform -1 0 3590 0 -1 270
box -12 -8 32 272
use FILL  FILL_2__2066_
timestamp 1701859473
transform -1 0 5370 0 -1 270
box -12 -8 32 272
use FILL  FILL_2__2067_
timestamp 1701859473
transform 1 0 7310 0 1 790
box -12 -8 32 272
use FILL  FILL_2__2068_
timestamp 1701859473
transform 1 0 5870 0 1 790
box -12 -8 32 272
use FILL  FILL_2__2069_
timestamp 1701859473
transform 1 0 3350 0 -1 1830
box -12 -8 32 272
use FILL  FILL_2__2070_
timestamp 1701859473
transform -1 0 3830 0 -1 1830
box -12 -8 32 272
use FILL  FILL_2__2071_
timestamp 1701859473
transform -1 0 5670 0 1 790
box -12 -8 32 272
use FILL  FILL_2__2072_
timestamp 1701859473
transform -1 0 7730 0 1 1310
box -12 -8 32 272
use FILL  FILL_2__2073_
timestamp 1701859473
transform 1 0 6610 0 1 1310
box -12 -8 32 272
use FILL  FILL_2__2074_
timestamp 1701859473
transform 1 0 1750 0 1 1310
box -12 -8 32 272
use FILL  FILL_2__2075_
timestamp 1701859473
transform -1 0 2230 0 1 1310
box -12 -8 32 272
use FILL  FILL_2__2076_
timestamp 1701859473
transform -1 0 2270 0 -1 1310
box -12 -8 32 272
use FILL  FILL_2__2077_
timestamp 1701859473
transform 1 0 4130 0 -1 1310
box -12 -8 32 272
use FILL  FILL_2__2078_
timestamp 1701859473
transform -1 0 2270 0 1 1830
box -12 -8 32 272
use FILL  FILL_2__2079_
timestamp 1701859473
transform -1 0 910 0 -1 1830
box -12 -8 32 272
use FILL  FILL_2__2080_
timestamp 1701859473
transform 1 0 2230 0 -1 1830
box -12 -8 32 272
use FILL  FILL_2__2081_
timestamp 1701859473
transform 1 0 2470 0 -1 1830
box -12 -8 32 272
use FILL  FILL_2__2082_
timestamp 1701859473
transform -1 0 2690 0 -1 1830
box -12 -8 32 272
use FILL  FILL_2__2083_
timestamp 1701859473
transform 1 0 4370 0 -1 1310
box -12 -8 32 272
use FILL  FILL_2__2084_
timestamp 1701859473
transform -1 0 5210 0 1 790
box -12 -8 32 272
use FILL  FILL_2__2085_
timestamp 1701859473
transform -1 0 5050 0 -1 270
box -12 -8 32 272
use FILL  FILL_2__2086_
timestamp 1701859473
transform -1 0 4270 0 -1 270
box -12 -8 32 272
use FILL  FILL_2__2087_
timestamp 1701859473
transform -1 0 4750 0 1 790
box -12 -8 32 272
use FILL  FILL_2__2088_
timestamp 1701859473
transform -1 0 5590 0 1 270
box -12 -8 32 272
use FILL  FILL_2__2089_
timestamp 1701859473
transform 1 0 5350 0 1 270
box -12 -8 32 272
use FILL  FILL_2__2090_
timestamp 1701859473
transform -1 0 4930 0 -1 790
box -12 -8 32 272
use FILL  FILL_2__2091_
timestamp 1701859473
transform 1 0 3150 0 1 790
box -12 -8 32 272
use FILL  FILL_2__2092_
timestamp 1701859473
transform 1 0 2710 0 -1 270
box -12 -8 32 272
use FILL  FILL_2__2093_
timestamp 1701859473
transform -1 0 2870 0 -1 790
box -12 -8 32 272
use FILL  FILL_2__2094_
timestamp 1701859473
transform 1 0 2270 0 -1 270
box -12 -8 32 272
use FILL  FILL_2__2095_
timestamp 1701859473
transform 1 0 2470 0 -1 270
box -12 -8 32 272
use FILL  FILL_2__2096_
timestamp 1701859473
transform -1 0 4930 0 1 270
box -12 -8 32 272
use FILL  FILL_2__2097_
timestamp 1701859473
transform -1 0 5150 0 1 270
box -12 -8 32 272
use FILL  FILL_2__2098_
timestamp 1701859473
transform 1 0 4690 0 1 270
box -12 -8 32 272
use FILL  FILL_2__2099_
timestamp 1701859473
transform 1 0 4010 0 -1 270
box -12 -8 32 272
use FILL  FILL_2__2100_
timestamp 1701859473
transform -1 0 5870 0 -1 1830
box -12 -8 32 272
use FILL  FILL_2__2101_
timestamp 1701859473
transform -1 0 5790 0 1 1310
box -12 -8 32 272
use FILL  FILL_2__2102_
timestamp 1701859473
transform -1 0 6190 0 1 1310
box -12 -8 32 272
use FILL  FILL_2__2103_
timestamp 1701859473
transform 1 0 5750 0 -1 1310
box -12 -8 32 272
use FILL  FILL_2__2104_
timestamp 1701859473
transform -1 0 5990 0 1 1310
box -12 -8 32 272
use FILL  FILL_2__2105_
timestamp 1701859473
transform -1 0 4290 0 -1 1830
box -12 -8 32 272
use FILL  FILL_2__2106_
timestamp 1701859473
transform 1 0 3970 0 -1 790
box -12 -8 32 272
use FILL  FILL_2__2107_
timestamp 1701859473
transform -1 0 3550 0 -1 790
box -12 -8 32 272
use FILL  FILL_2__2108_
timestamp 1701859473
transform 1 0 2910 0 1 790
box -12 -8 32 272
use FILL  FILL_2__2109_
timestamp 1701859473
transform -1 0 3330 0 -1 790
box -12 -8 32 272
use FILL  FILL_2__2110_
timestamp 1701859473
transform 1 0 3090 0 -1 790
box -12 -8 32 272
use FILL  FILL_2__2111_
timestamp 1701859473
transform -1 0 3770 0 -1 790
box -12 -8 32 272
use FILL  FILL_2__2112_
timestamp 1701859473
transform -1 0 5130 0 -1 790
box -12 -8 32 272
use FILL  FILL_2__2113_
timestamp 1701859473
transform -1 0 5110 0 1 1310
box -12 -8 32 272
use FILL  FILL_2__2114_
timestamp 1701859473
transform -1 0 5550 0 1 1310
box -12 -8 32 272
use FILL  FILL_2__2115_
timestamp 1701859473
transform -1 0 5590 0 -1 790
box -12 -8 32 272
use FILL  FILL_2__2116_
timestamp 1701859473
transform 1 0 2410 0 1 1310
box -12 -8 32 272
use FILL  FILL_2__2117_
timestamp 1701859473
transform 1 0 2610 0 1 1310
box -12 -8 32 272
use FILL  FILL_2__2118_
timestamp 1701859473
transform 1 0 3790 0 1 1310
box -12 -8 32 272
use FILL  FILL_2__2119_
timestamp 1701859473
transform -1 0 4050 0 1 1310
box -12 -8 32 272
use FILL  FILL_2__2120_
timestamp 1701859473
transform 1 0 3910 0 -1 1310
box -12 -8 32 272
use FILL  FILL_2__2121_
timestamp 1701859473
transform -1 0 4490 0 1 270
box -12 -8 32 272
use FILL  FILL_2__2122_
timestamp 1701859473
transform -1 0 2830 0 1 2350
box -12 -8 32 272
use FILL  FILL_2__2123_
timestamp 1701859473
transform 1 0 2770 0 -1 2350
box -12 -8 32 272
use FILL  FILL_2__2124_
timestamp 1701859473
transform -1 0 3670 0 -1 2350
box -12 -8 32 272
use FILL  FILL_2__2125_
timestamp 1701859473
transform 1 0 5790 0 -1 3390
box -12 -8 32 272
use FILL  FILL_2__2126_
timestamp 1701859473
transform 1 0 5470 0 1 2870
box -12 -8 32 272
use FILL  FILL_2__2127_
timestamp 1701859473
transform -1 0 5950 0 1 2870
box -12 -8 32 272
use FILL  FILL_2__2128_
timestamp 1701859473
transform 1 0 4570 0 1 2870
box -12 -8 32 272
use FILL  FILL_2__2129_
timestamp 1701859473
transform 1 0 5250 0 1 2870
box -12 -8 32 272
use FILL  FILL_2__2130_
timestamp 1701859473
transform -1 0 4610 0 -1 2350
box -12 -8 32 272
use FILL  FILL_2__2131_
timestamp 1701859473
transform 1 0 4650 0 1 1310
box -12 -8 32 272
use FILL  FILL_2__2132_
timestamp 1701859473
transform -1 0 4530 0 1 790
box -12 -8 32 272
use FILL  FILL_2__2133_
timestamp 1701859473
transform 1 0 4450 0 -1 790
box -12 -8 32 272
use FILL  FILL_2__2134_
timestamp 1701859473
transform 1 0 3570 0 -1 2870
box -12 -8 32 272
use FILL  FILL_2__2135_
timestamp 1701859473
transform 1 0 4190 0 -1 3390
box -12 -8 32 272
use FILL  FILL_2__2136_
timestamp 1701859473
transform -1 0 2730 0 1 3390
box -12 -8 32 272
use FILL  FILL_2__2137_
timestamp 1701859473
transform 1 0 2290 0 1 3390
box -12 -8 32 272
use FILL  FILL_2__2138_
timestamp 1701859473
transform 1 0 3090 0 -1 4430
box -12 -8 32 272
use FILL  FILL_2__2139_
timestamp 1701859473
transform -1 0 2870 0 -1 4430
box -12 -8 32 272
use FILL  FILL_2__2140_
timestamp 1701859473
transform 1 0 2790 0 1 4430
box -12 -8 32 272
use FILL  FILL_2__2141_
timestamp 1701859473
transform -1 0 3030 0 1 4430
box -12 -8 32 272
use FILL  FILL_2__2142_
timestamp 1701859473
transform 1 0 2910 0 1 3390
box -12 -8 32 272
use FILL  FILL_2__2143_
timestamp 1701859473
transform -1 0 7410 0 -1 3390
box -12 -8 32 272
use FILL  FILL_2__2144_
timestamp 1701859473
transform 1 0 2050 0 1 2870
box -12 -8 32 272
use FILL  FILL_2__2145_
timestamp 1701859473
transform -1 0 10030 0 -1 2870
box -12 -8 32 272
use FILL  FILL_2__2146_
timestamp 1701859473
transform -1 0 7610 0 -1 3390
box -12 -8 32 272
use FILL  FILL_2__2147_
timestamp 1701859473
transform 1 0 7570 0 -1 3910
box -12 -8 32 272
use FILL  FILL_2__2148_
timestamp 1701859473
transform 1 0 7410 0 1 3390
box -12 -8 32 272
use FILL  FILL_2__2149_
timestamp 1701859473
transform 1 0 7610 0 1 3390
box -12 -8 32 272
use FILL  FILL_2__2150_
timestamp 1701859473
transform -1 0 7870 0 1 3390
box -12 -8 32 272
use FILL  FILL_2__2151_
timestamp 1701859473
transform 1 0 7150 0 -1 3390
box -12 -8 32 272
use FILL  FILL_2__2152_
timestamp 1701859473
transform 1 0 6910 0 -1 3390
box -12 -8 32 272
use FILL  FILL_2__2153_
timestamp 1701859473
transform -1 0 6050 0 -1 3390
box -12 -8 32 272
use FILL  FILL_2__2154_
timestamp 1701859473
transform 1 0 2810 0 -1 7030
box -12 -8 32 272
use FILL  FILL_2__2155_
timestamp 1701859473
transform 1 0 6370 0 1 5990
box -12 -8 32 272
use FILL  FILL_2__2156_
timestamp 1701859473
transform -1 0 4590 0 1 3910
box -12 -8 32 272
use FILL  FILL_2__2157_
timestamp 1701859473
transform -1 0 4730 0 -1 4430
box -12 -8 32 272
use FILL  FILL_2__2158_
timestamp 1701859473
transform -1 0 2590 0 1 2350
box -12 -8 32 272
use FILL  FILL_2__2159_
timestamp 1701859473
transform 1 0 3490 0 1 3910
box -12 -8 32 272
use FILL  FILL_2__2160_
timestamp 1701859473
transform -1 0 3810 0 -1 4430
box -12 -8 32 272
use FILL  FILL_2__2161_
timestamp 1701859473
transform -1 0 3950 0 1 3910
box -12 -8 32 272
use FILL  FILL_2__2162_
timestamp 1701859473
transform -1 0 4390 0 1 3910
box -12 -8 32 272
use FILL  FILL_2__2163_
timestamp 1701859473
transform 1 0 3710 0 -1 3910
box -12 -8 32 272
use FILL  FILL_2__2164_
timestamp 1701859473
transform -1 0 530 0 -1 4950
box -12 -8 32 272
use FILL  FILL_2__2165_
timestamp 1701859473
transform -1 0 3230 0 -1 3910
box -12 -8 32 272
use FILL  FILL_2__2166_
timestamp 1701859473
transform 1 0 3930 0 -1 3910
box -12 -8 32 272
use FILL  FILL_2__2167_
timestamp 1701859473
transform 1 0 4130 0 1 3910
box -12 -8 32 272
use FILL  FILL_2__2168_
timestamp 1701859473
transform 1 0 3050 0 1 3910
box -12 -8 32 272
use FILL  FILL_2__2169_
timestamp 1701859473
transform 1 0 2410 0 -1 4430
box -12 -8 32 272
use FILL  FILL_2__2170_
timestamp 1701859473
transform -1 0 2670 0 -1 4430
box -12 -8 32 272
use FILL  FILL_2__2171_
timestamp 1701859473
transform 1 0 4010 0 -1 4430
box -12 -8 32 272
use FILL  FILL_2__2172_
timestamp 1701859473
transform 1 0 4250 0 -1 4430
box -12 -8 32 272
use FILL  FILL_2__2173_
timestamp 1701859473
transform -1 0 4490 0 -1 4430
box -12 -8 32 272
use FILL  FILL_2__2174_
timestamp 1701859473
transform 1 0 5990 0 1 7030
box -12 -8 32 272
use FILL  FILL_2__2175_
timestamp 1701859473
transform -1 0 2490 0 1 8070
box -12 -8 32 272
use FILL  FILL_2__2176_
timestamp 1701859473
transform -1 0 6410 0 -1 8070
box -12 -8 32 272
use FILL  FILL_2__2177_
timestamp 1701859473
transform 1 0 4930 0 1 8070
box -12 -8 32 272
use FILL  FILL_2__2178_
timestamp 1701859473
transform -1 0 4110 0 -1 8590
box -12 -8 32 272
use FILL  FILL_2__2179_
timestamp 1701859473
transform -1 0 5930 0 -1 8070
box -12 -8 32 272
use FILL  FILL_2__2180_
timestamp 1701859473
transform -1 0 2950 0 -1 9630
box -12 -8 32 272
use FILL  FILL_2__2181_
timestamp 1701859473
transform 1 0 5010 0 1 7550
box -12 -8 32 272
use FILL  FILL_2__2182_
timestamp 1701859473
transform 1 0 5530 0 -1 10150
box -12 -8 32 272
use FILL  FILL_2__2183_
timestamp 1701859473
transform -1 0 3510 0 1 10150
box -12 -8 32 272
use FILL  FILL_2__2184_
timestamp 1701859473
transform 1 0 4330 0 1 8070
box -12 -8 32 272
use FILL  FILL_2__2185_
timestamp 1701859473
transform 1 0 5930 0 1 10150
box -12 -8 32 272
use FILL  FILL_2__2186_
timestamp 1701859473
transform 1 0 3490 0 1 10670
box -12 -8 32 272
use FILL  FILL_2__2187_
timestamp 1701859473
transform -1 0 5410 0 -1 10670
box -12 -8 32 272
use FILL  FILL_2__2188_
timestamp 1701859473
transform 1 0 2090 0 -1 10670
box -12 -8 32 272
use FILL  FILL_2__2189_
timestamp 1701859473
transform 1 0 5650 0 -1 10670
box -12 -8 32 272
use FILL  FILL_2__2190_
timestamp 1701859473
transform -1 0 2810 0 1 10150
box -12 -8 32 272
use FILL  FILL_2__2191_
timestamp 1701859473
transform -1 0 5290 0 -1 10150
box -12 -8 32 272
use FILL  FILL_2__2192_
timestamp 1701859473
transform -1 0 11090 0 1 3910
box -12 -8 32 272
use FILL  FILL_2__2193_
timestamp 1701859473
transform 1 0 1210 0 -1 3910
box -12 -8 32 272
use FILL  FILL_2__2194_
timestamp 1701859473
transform 1 0 1010 0 -1 3910
box -12 -8 32 272
use FILL  FILL_2__2195_
timestamp 1701859473
transform 1 0 2590 0 1 3910
box -12 -8 32 272
use FILL  FILL_2__2196_
timestamp 1701859473
transform 1 0 2830 0 1 3910
box -12 -8 32 272
use FILL  FILL_2__2197_
timestamp 1701859473
transform 1 0 5310 0 1 3910
box -12 -8 32 272
use FILL  FILL_2__2198_
timestamp 1701859473
transform 1 0 250 0 1 1830
box -12 -8 32 272
use FILL  FILL_2__2199_
timestamp 1701859473
transform -1 0 2810 0 -1 3910
box -12 -8 32 272
use FILL  FILL_2__2200_
timestamp 1701859473
transform 1 0 5330 0 -1 3910
box -12 -8 32 272
use FILL  FILL_2__2201_
timestamp 1701859473
transform -1 0 5570 0 1 3910
box -12 -8 32 272
use FILL  FILL_2__2202_
timestamp 1701859473
transform -1 0 8150 0 -1 4430
box -12 -8 32 272
use FILL  FILL_2__2203_
timestamp 1701859473
transform -1 0 4870 0 -1 3910
box -12 -8 32 272
use FILL  FILL_2__2204_
timestamp 1701859473
transform 1 0 5090 0 -1 3910
box -12 -8 32 272
use FILL  FILL_2__2205_
timestamp 1701859473
transform -1 0 8950 0 -1 3910
box -12 -8 32 272
use FILL  FILL_2__2206_
timestamp 1701859473
transform 1 0 9030 0 1 3910
box -12 -8 32 272
use FILL  FILL_2__2207_
timestamp 1701859473
transform 1 0 9490 0 -1 3910
box -12 -8 32 272
use FILL  FILL_2__2208_
timestamp 1701859473
transform -1 0 9750 0 -1 3910
box -12 -8 32 272
use FILL  FILL_2__2209_
timestamp 1701859473
transform -1 0 9550 0 1 4430
box -12 -8 32 272
use FILL  FILL_2__2210_
timestamp 1701859473
transform -1 0 10550 0 -1 4950
box -12 -8 32 272
use FILL  FILL_2__2211_
timestamp 1701859473
transform 1 0 9250 0 -1 3910
box -12 -8 32 272
use FILL  FILL_2__2212_
timestamp 1701859473
transform -1 0 8830 0 1 3910
box -12 -8 32 272
use FILL  FILL_2__2213_
timestamp 1701859473
transform -1 0 9270 0 1 3910
box -12 -8 32 272
use FILL  FILL_2__2214_
timestamp 1701859473
transform -1 0 9470 0 -1 4430
box -12 -8 32 272
use FILL  FILL_2__2215_
timestamp 1701859473
transform 1 0 9670 0 -1 4430
box -12 -8 32 272
use FILL  FILL_2__2216_
timestamp 1701859473
transform -1 0 9430 0 -1 7030
box -12 -8 32 272
use FILL  FILL_2__2217_
timestamp 1701859473
transform 1 0 9210 0 -1 4430
box -12 -8 32 272
use FILL  FILL_2__2218_
timestamp 1701859473
transform -1 0 9730 0 1 3910
box -12 -8 32 272
use FILL  FILL_2__2219_
timestamp 1701859473
transform 1 0 9910 0 1 3910
box -12 -8 32 272
use FILL  FILL_2__2220_
timestamp 1701859473
transform 1 0 10290 0 -1 4950
box -12 -8 32 272
use FILL  FILL_2__2221_
timestamp 1701859473
transform -1 0 9670 0 -1 7030
box -12 -8 32 272
use FILL  FILL_2__2222_
timestamp 1701859473
transform 1 0 10030 0 1 4430
box -12 -8 32 272
use FILL  FILL_2__2223_
timestamp 1701859473
transform -1 0 9930 0 -1 4430
box -12 -8 32 272
use FILL  FILL_2__2224_
timestamp 1701859473
transform -1 0 9790 0 1 4430
box -12 -8 32 272
use FILL  FILL_2__2225_
timestamp 1701859473
transform 1 0 10030 0 -1 4950
box -12 -8 32 272
use FILL  FILL_2__2226_
timestamp 1701859473
transform 1 0 8910 0 -1 7030
box -12 -8 32 272
use FILL  FILL_2__2227_
timestamp 1701859473
transform -1 0 9190 0 -1 7030
box -12 -8 32 272
use FILL  FILL_2__2228_
timestamp 1701859473
transform -1 0 5730 0 -1 7030
box -12 -8 32 272
use FILL  FILL_2__2229_
timestamp 1701859473
transform 1 0 4290 0 1 3390
box -12 -8 32 272
use FILL  FILL_2__2230_
timestamp 1701859473
transform -1 0 4390 0 -1 3910
box -12 -8 32 272
use FILL  FILL_2__2231_
timestamp 1701859473
transform -1 0 4170 0 -1 3910
box -12 -8 32 272
use FILL  FILL_2__2232_
timestamp 1701859473
transform 1 0 1570 0 1 2870
box -12 -8 32 272
use FILL  FILL_2__2233_
timestamp 1701859473
transform 1 0 2290 0 1 2870
box -12 -8 32 272
use FILL  FILL_2__2234_
timestamp 1701859473
transform -1 0 2550 0 1 2870
box -12 -8 32 272
use FILL  FILL_2__2235_
timestamp 1701859473
transform 1 0 6310 0 1 3390
box -12 -8 32 272
use FILL  FILL_2__2236_
timestamp 1701859473
transform -1 0 5590 0 -1 3910
box -12 -8 32 272
use FILL  FILL_2__2237_
timestamp 1701859473
transform -1 0 4630 0 -1 3910
box -12 -8 32 272
use FILL  FILL_2__2238_
timestamp 1701859473
transform 1 0 4690 0 -1 4950
box -12 -8 32 272
use FILL  FILL_2__2239_
timestamp 1701859473
transform 1 0 2810 0 1 4950
box -12 -8 32 272
use FILL  FILL_2__2240_
timestamp 1701859473
transform 1 0 2370 0 1 3910
box -12 -8 32 272
use FILL  FILL_2__2241_
timestamp 1701859473
transform -1 0 2390 0 1 4950
box -12 -8 32 272
use FILL  FILL_2__2242_
timestamp 1701859473
transform 1 0 2430 0 -1 4950
box -12 -8 32 272
use FILL  FILL_2__2243_
timestamp 1701859473
transform 1 0 2610 0 1 4950
box -12 -8 32 272
use FILL  FILL_2__2244_
timestamp 1701859473
transform 1 0 3030 0 1 4950
box -12 -8 32 272
use FILL  FILL_2__2245_
timestamp 1701859473
transform 1 0 2870 0 1 5990
box -12 -8 32 272
use FILL  FILL_2__2246_
timestamp 1701859473
transform 1 0 2890 0 -1 4950
box -12 -8 32 272
use FILL  FILL_2__2247_
timestamp 1701859473
transform -1 0 3010 0 -1 6510
box -12 -8 32 272
use FILL  FILL_2__2248_
timestamp 1701859473
transform 1 0 3470 0 -1 7030
box -12 -8 32 272
use FILL  FILL_2__2249_
timestamp 1701859473
transform 1 0 6250 0 1 7030
box -12 -8 32 272
use FILL  FILL_2__2250_
timestamp 1701859473
transform -1 0 10550 0 -1 7550
box -12 -8 32 272
use FILL  FILL_2__2251_
timestamp 1701859473
transform -1 0 10610 0 1 8070
box -12 -8 32 272
use FILL  FILL_2__2252_
timestamp 1701859473
transform -1 0 10910 0 -1 8070
box -12 -8 32 272
use FILL  FILL_2__2253_
timestamp 1701859473
transform -1 0 10670 0 -1 8070
box -12 -8 32 272
use FILL  FILL_2__2254_
timestamp 1701859473
transform 1 0 5370 0 1 8070
box -12 -8 32 272
use FILL  FILL_2__2255_
timestamp 1701859473
transform 1 0 2990 0 1 7030
box -12 -8 32 272
use FILL  FILL_2__2256_
timestamp 1701859473
transform -1 0 5110 0 1 7030
box -12 -8 32 272
use FILL  FILL_2__2257_
timestamp 1701859473
transform 1 0 5050 0 -1 7550
box -12 -8 32 272
use FILL  FILL_2__2258_
timestamp 1701859473
transform 1 0 5690 0 -1 8590
box -12 -8 32 272
use FILL  FILL_2__2259_
timestamp 1701859473
transform 1 0 10310 0 -1 7550
box -12 -8 32 272
use FILL  FILL_2__2260_
timestamp 1701859473
transform 1 0 9890 0 1 8070
box -12 -8 32 272
use FILL  FILL_2__2261_
timestamp 1701859473
transform -1 0 10190 0 1 7550
box -12 -8 32 272
use FILL  FILL_2__2262_
timestamp 1701859473
transform -1 0 9950 0 1 7550
box -12 -8 32 272
use FILL  FILL_2__2263_
timestamp 1701859473
transform 1 0 5450 0 1 7550
box -12 -8 32 272
use FILL  FILL_2__2264_
timestamp 1701859473
transform 1 0 1610 0 -1 6510
box -12 -8 32 272
use FILL  FILL_2__2265_
timestamp 1701859473
transform 1 0 1790 0 -1 6510
box -12 -8 32 272
use FILL  FILL_2__2266_
timestamp 1701859473
transform 1 0 3890 0 1 6510
box -12 -8 32 272
use FILL  FILL_2__2267_
timestamp 1701859473
transform -1 0 3650 0 -1 7550
box -12 -8 32 272
use FILL  FILL_2__2268_
timestamp 1701859473
transform 1 0 4330 0 -1 7550
box -12 -8 32 272
use FILL  FILL_2__2269_
timestamp 1701859473
transform 1 0 5650 0 1 7550
box -12 -8 32 272
use FILL  FILL_2__2270_
timestamp 1701859473
transform 1 0 8570 0 1 7550
box -12 -8 32 272
use FILL  FILL_2__2271_
timestamp 1701859473
transform -1 0 8850 0 -1 8070
box -12 -8 32 272
use FILL  FILL_2__2272_
timestamp 1701859473
transform -1 0 9110 0 -1 8070
box -12 -8 32 272
use FILL  FILL_2__2273_
timestamp 1701859473
transform -1 0 8610 0 -1 8070
box -12 -8 32 272
use FILL  FILL_2__2274_
timestamp 1701859473
transform -1 0 5970 0 -1 9630
box -12 -8 32 272
use FILL  FILL_2__2275_
timestamp 1701859473
transform -1 0 2270 0 1 8070
box -12 -8 32 272
use FILL  FILL_2__2276_
timestamp 1701859473
transform -1 0 3150 0 1 8070
box -12 -8 32 272
use FILL  FILL_2__2277_
timestamp 1701859473
transform -1 0 3630 0 -1 8590
box -12 -8 32 272
use FILL  FILL_2__2278_
timestamp 1701859473
transform 1 0 6530 0 1 9110
box -12 -8 32 272
use FILL  FILL_2__2279_
timestamp 1701859473
transform -1 0 10230 0 1 5990
box -12 -8 32 272
use FILL  FILL_2__2280_
timestamp 1701859473
transform 1 0 10410 0 1 5990
box -12 -8 32 272
use FILL  FILL_2__2281_
timestamp 1701859473
transform -1 0 10690 0 -1 5990
box -12 -8 32 272
use FILL  FILL_2__2282_
timestamp 1701859473
transform -1 0 10470 0 -1 6510
box -12 -8 32 272
use FILL  FILL_2__2283_
timestamp 1701859473
transform 1 0 5930 0 -1 8590
box -12 -8 32 272
use FILL  FILL_2__2284_
timestamp 1701859473
transform -1 0 2050 0 1 8070
box -12 -8 32 272
use FILL  FILL_2__2285_
timestamp 1701859473
transform -1 0 4110 0 1 8070
box -12 -8 32 272
use FILL  FILL_2__2286_
timestamp 1701859473
transform 1 0 5010 0 -1 8590
box -12 -8 32 272
use FILL  FILL_2__2287_
timestamp 1701859473
transform -1 0 6090 0 1 8590
box -12 -8 32 272
use FILL  FILL_2__2288_
timestamp 1701859473
transform -1 0 8810 0 1 7550
box -12 -8 32 272
use FILL  FILL_2__2289_
timestamp 1701859473
transform 1 0 8470 0 1 8070
box -12 -8 32 272
use FILL  FILL_2__2290_
timestamp 1701859473
transform -1 0 9970 0 -1 8070
box -12 -8 32 272
use FILL  FILL_2__2291_
timestamp 1701859473
transform -1 0 8750 0 1 8070
box -12 -8 32 272
use FILL  FILL_2__2292_
timestamp 1701859473
transform -1 0 6190 0 -1 9110
box -12 -8 32 272
use FILL  FILL_2__2293_
timestamp 1701859473
transform -1 0 2510 0 -1 8590
box -12 -8 32 272
use FILL  FILL_2__2294_
timestamp 1701859473
transform -1 0 3990 0 1 8590
box -12 -8 32 272
use FILL  FILL_2__2295_
timestamp 1701859473
transform 1 0 4910 0 1 8590
box -12 -8 32 272
use FILL  FILL_2__2296_
timestamp 1701859473
transform 1 0 6630 0 -1 9110
box -12 -8 32 272
use FILL  FILL_2__2297_
timestamp 1701859473
transform -1 0 9530 0 -1 5990
box -12 -8 32 272
use FILL  FILL_2__2298_
timestamp 1701859473
transform -1 0 9970 0 -1 5470
box -12 -8 32 272
use FILL  FILL_2__2299_
timestamp 1701859473
transform -1 0 9310 0 -1 6510
box -12 -8 32 272
use FILL  FILL_2__2300_
timestamp 1701859473
transform 1 0 9510 0 1 5990
box -12 -8 32 272
use FILL  FILL_2__2301_
timestamp 1701859473
transform 1 0 5550 0 1 9630
box -12 -8 32 272
use FILL  FILL_2__2302_
timestamp 1701859473
transform -1 0 3450 0 -1 9110
box -12 -8 32 272
use FILL  FILL_2__2303_
timestamp 1701859473
transform 1 0 2570 0 1 9110
box -12 -8 32 272
use FILL  FILL_2__2304_
timestamp 1701859473
transform 1 0 2770 0 -1 9110
box -12 -8 32 272
use FILL  FILL_2__2305_
timestamp 1701859473
transform -1 0 3750 0 1 8590
box -12 -8 32 272
use FILL  FILL_2__2306_
timestamp 1701859473
transform 1 0 4430 0 1 8590
box -12 -8 32 272
use FILL  FILL_2__2307_
timestamp 1701859473
transform 1 0 6290 0 1 9110
box -12 -8 32 272
use FILL  FILL_2__2308_
timestamp 1701859473
transform -1 0 8870 0 -1 6510
box -12 -8 32 272
use FILL  FILL_2__2309_
timestamp 1701859473
transform -1 0 8570 0 1 5990
box -12 -8 32 272
use FILL  FILL_2__2310_
timestamp 1701859473
transform -1 0 9070 0 -1 6510
box -12 -8 32 272
use FILL  FILL_2__2311_
timestamp 1701859473
transform -1 0 8630 0 -1 6510
box -12 -8 32 272
use FILL  FILL_2__2312_
timestamp 1701859473
transform -1 0 5530 0 -1 9630
box -12 -8 32 272
use FILL  FILL_2__2313_
timestamp 1701859473
transform -1 0 1810 0 1 8590
box -12 -8 32 272
use FILL  FILL_2__2314_
timestamp 1701859473
transform 1 0 1410 0 -1 8590
box -12 -8 32 272
use FILL  FILL_2__2315_
timestamp 1701859473
transform 1 0 1850 0 -1 8590
box -12 -8 32 272
use FILL  FILL_2__2316_
timestamp 1701859473
transform -1 0 4210 0 1 8590
box -12 -8 32 272
use FILL  FILL_2__2317_
timestamp 1701859473
transform 1 0 4670 0 1 8590
box -12 -8 32 272
use FILL  FILL_2__2318_
timestamp 1701859473
transform 1 0 6770 0 1 9110
box -12 -8 32 272
use FILL  FILL_2__2319_
timestamp 1701859473
transform -1 0 11090 0 1 4430
box -12 -8 32 272
use FILL  FILL_2__2320_
timestamp 1701859473
transform 1 0 5070 0 1 3910
box -12 -8 32 272
use FILL  FILL_2__2321_
timestamp 1701859473
transform 1 0 6490 0 1 3910
box -12 -8 32 272
use FILL  FILL_2__2322_
timestamp 1701859473
transform -1 0 7870 0 1 3910
box -12 -8 32 272
use FILL  FILL_2__2323_
timestamp 1701859473
transform 1 0 7910 0 -1 4430
box -12 -8 32 272
use FILL  FILL_2__2324_
timestamp 1701859473
transform -1 0 11130 0 -1 2870
box -12 -8 32 272
use FILL  FILL_2__2325_
timestamp 1701859473
transform -1 0 8110 0 1 3910
box -12 -8 32 272
use FILL  FILL_2__2326_
timestamp 1701859473
transform -1 0 3150 0 -1 4950
box -12 -8 32 272
use FILL  FILL_2__2327_
timestamp 1701859473
transform -1 0 3350 0 -1 4950
box -12 -8 32 272
use FILL  FILL_2__2328_
timestamp 1701859473
transform 1 0 3830 0 -1 5470
box -12 -8 32 272
use FILL  FILL_2__2329_
timestamp 1701859473
transform 1 0 3590 0 -1 5470
box -12 -8 32 272
use FILL  FILL_2__2330_
timestamp 1701859473
transform 1 0 3730 0 1 4950
box -12 -8 32 272
use FILL  FILL_2__2331_
timestamp 1701859473
transform 1 0 4810 0 1 3910
box -12 -8 32 272
use FILL  FILL_2__2332_
timestamp 1701859473
transform -1 0 4150 0 1 4950
box -12 -8 32 272
use FILL  FILL_2__2333_
timestamp 1701859473
transform -1 0 11110 0 -1 4430
box -12 -8 32 272
use FILL  FILL_2__2334_
timestamp 1701859473
transform 1 0 8990 0 -1 4430
box -12 -8 32 272
use FILL  FILL_2__2335_
timestamp 1701859473
transform 1 0 5170 0 -1 5470
box -12 -8 32 272
use FILL  FILL_2__2336_
timestamp 1701859473
transform -1 0 5030 0 1 5990
box -12 -8 32 272
use FILL  FILL_2__2337_
timestamp 1701859473
transform 1 0 4530 0 1 3390
box -12 -8 32 272
use FILL  FILL_2__2338_
timestamp 1701859473
transform 1 0 3130 0 1 3390
box -12 -8 32 272
use FILL  FILL_2__2339_
timestamp 1701859473
transform 1 0 4710 0 1 3390
box -12 -8 32 272
use FILL  FILL_2__2340_
timestamp 1701859473
transform 1 0 4950 0 1 3390
box -12 -8 32 272
use FILL  FILL_2__2341_
timestamp 1701859473
transform -1 0 530 0 1 5990
box -12 -8 32 272
use FILL  FILL_2__2342_
timestamp 1701859473
transform 1 0 2630 0 1 5470
box -12 -8 32 272
use FILL  FILL_2__2343_
timestamp 1701859473
transform -1 0 4570 0 1 6510
box -12 -8 32 272
use FILL  FILL_2__2344_
timestamp 1701859473
transform -1 0 4850 0 1 5470
box -12 -8 32 272
use FILL  FILL_2__2345_
timestamp 1701859473
transform -1 0 4650 0 1 5470
box -12 -8 32 272
use FILL  FILL_2__2346_
timestamp 1701859473
transform -1 0 4810 0 -1 5990
box -12 -8 32 272
use FILL  FILL_2__2347_
timestamp 1701859473
transform -1 0 5670 0 -1 5990
box -12 -8 32 272
use FILL  FILL_2__2348_
timestamp 1701859473
transform 1 0 5230 0 -1 6510
box -12 -8 32 272
use FILL  FILL_2__2349_
timestamp 1701859473
transform -1 0 5010 0 -1 6510
box -12 -8 32 272
use FILL  FILL_2__2350_
timestamp 1701859473
transform -1 0 4430 0 -1 6510
box -12 -8 32 272
use FILL  FILL_2__2351_
timestamp 1701859473
transform 1 0 5570 0 1 7030
box -12 -8 32 272
use FILL  FILL_2__2352_
timestamp 1701859473
transform -1 0 5790 0 1 7030
box -12 -8 32 272
use FILL  FILL_2__2353_
timestamp 1701859473
transform -1 0 730 0 1 7030
box -12 -8 32 272
use FILL  FILL_2__2354_
timestamp 1701859473
transform 1 0 5430 0 -1 5990
box -12 -8 32 272
use FILL  FILL_2__2355_
timestamp 1701859473
transform 1 0 5330 0 1 7030
box -12 -8 32 272
use FILL  FILL_2__2356_
timestamp 1701859473
transform -1 0 4830 0 -1 7550
box -12 -8 32 272
use FILL  FILL_2__2357_
timestamp 1701859473
transform 1 0 4690 0 1 8070
box -12 -8 32 272
use FILL  FILL_2__2358_
timestamp 1701859473
transform 1 0 5170 0 1 8070
box -12 -8 32 272
use FILL  FILL_2__2359_
timestamp 1701859473
transform -1 0 5490 0 -1 8590
box -12 -8 32 272
use FILL  FILL_2__2360_
timestamp 1701859473
transform -1 0 730 0 -1 6510
box -12 -8 32 272
use FILL  FILL_2__2361_
timestamp 1701859473
transform -1 0 5230 0 1 5990
box -12 -8 32 272
use FILL  FILL_2__2362_
timestamp 1701859473
transform 1 0 5230 0 1 6510
box -12 -8 32 272
use FILL  FILL_2__2363_
timestamp 1701859473
transform 1 0 5250 0 -1 7030
box -12 -8 32 272
use FILL  FILL_2__2364_
timestamp 1701859473
transform 1 0 5250 0 -1 8070
box -12 -8 32 272
use FILL  FILL_2__2365_
timestamp 1701859473
transform 1 0 5490 0 -1 8070
box -12 -8 32 272
use FILL  FILL_2__2366_
timestamp 1701859473
transform -1 0 5710 0 -1 8070
box -12 -8 32 272
use FILL  FILL_2__2367_
timestamp 1701859473
transform 1 0 2670 0 -1 7550
box -12 -8 32 272
use FILL  FILL_2__2368_
timestamp 1701859473
transform -1 0 5510 0 -1 7030
box -12 -8 32 272
use FILL  FILL_2__2369_
timestamp 1701859473
transform 1 0 5210 0 1 7550
box -12 -8 32 272
use FILL  FILL_2__2370_
timestamp 1701859473
transform -1 0 5250 0 -1 8590
box -12 -8 32 272
use FILL  FILL_2__2371_
timestamp 1701859473
transform 1 0 5930 0 -1 9110
box -12 -8 32 272
use FILL  FILL_2__2372_
timestamp 1701859473
transform 1 0 6090 0 1 9110
box -12 -8 32 272
use FILL  FILL_2__2373_
timestamp 1701859473
transform -1 0 6170 0 -1 9630
box -12 -8 32 272
use FILL  FILL_2__2374_
timestamp 1701859473
transform 1 0 50 0 -1 9110
box -12 -8 32 272
use FILL  FILL_2__2375_
timestamp 1701859473
transform -1 0 4190 0 1 5470
box -12 -8 32 272
use FILL  FILL_2__2376_
timestamp 1701859473
transform 1 0 4530 0 -1 5990
box -12 -8 32 272
use FILL  FILL_2__2377_
timestamp 1701859473
transform -1 0 3950 0 -1 6510
box -12 -8 32 272
use FILL  FILL_2__2378_
timestamp 1701859473
transform 1 0 3690 0 -1 6510
box -12 -8 32 272
use FILL  FILL_2__2379_
timestamp 1701859473
transform -1 0 5010 0 1 6510
box -12 -8 32 272
use FILL  FILL_2__2380_
timestamp 1701859473
transform -1 0 4790 0 -1 8590
box -12 -8 32 272
use FILL  FILL_2__2381_
timestamp 1701859473
transform 1 0 3850 0 -1 8590
box -12 -8 32 272
use FILL  FILL_2__2382_
timestamp 1701859473
transform -1 0 4550 0 -1 8590
box -12 -8 32 272
use FILL  FILL_2__2383_
timestamp 1701859473
transform -1 0 5630 0 1 8590
box -12 -8 32 272
use FILL  FILL_2__2384_
timestamp 1701859473
transform -1 0 5850 0 1 8590
box -12 -8 32 272
use FILL  FILL_2__2385_
timestamp 1701859473
transform 1 0 1230 0 -1 10150
box -12 -8 32 272
use FILL  FILL_2__2386_
timestamp 1701859473
transform 1 0 5490 0 -1 7550
box -12 -8 32 272
use FILL  FILL_2__2387_
timestamp 1701859473
transform 1 0 5470 0 -1 9110
box -12 -8 32 272
use FILL  FILL_2__2388_
timestamp 1701859473
transform -1 0 5270 0 -1 9110
box -12 -8 32 272
use FILL  FILL_2__2389_
timestamp 1701859473
transform -1 0 5050 0 -1 9630
box -12 -8 32 272
use FILL  FILL_2__2390_
timestamp 1701859473
transform 1 0 5110 0 1 9630
box -12 -8 32 272
use FILL  FILL_2__2391_
timestamp 1701859473
transform -1 0 5330 0 1 9630
box -12 -8 32 272
use FILL  FILL_2__2392_
timestamp 1701859473
transform 1 0 1430 0 -1 10150
box -12 -8 32 272
use FILL  FILL_2__2393_
timestamp 1701859473
transform -1 0 5290 0 -1 7550
box -12 -8 32 272
use FILL  FILL_2__2394_
timestamp 1701859473
transform 1 0 5370 0 1 8590
box -12 -8 32 272
use FILL  FILL_2__2395_
timestamp 1701859473
transform -1 0 5730 0 -1 9110
box -12 -8 32 272
use FILL  FILL_2__2396_
timestamp 1701859473
transform 1 0 5650 0 1 9110
box -12 -8 32 272
use FILL  FILL_2__2397_
timestamp 1701859473
transform 1 0 5890 0 1 9110
box -12 -8 32 272
use FILL  FILL_2__2398_
timestamp 1701859473
transform 1 0 5710 0 -1 9630
box -12 -8 32 272
use FILL  FILL_2__2399_
timestamp 1701859473
transform -1 0 3150 0 -1 5470
box -12 -8 32 272
use FILL  FILL_2__2400_
timestamp 1701859473
transform -1 0 3330 0 1 5990
box -12 -8 32 272
use FILL  FILL_2__2401_
timestamp 1701859473
transform 1 0 3250 0 -1 6510
box -12 -8 32 272
use FILL  FILL_2__2402_
timestamp 1701859473
transform -1 0 2190 0 -1 4430
box -12 -8 32 272
use FILL  FILL_2__2403_
timestamp 1701859473
transform -1 0 2590 0 1 4430
box -12 -8 32 272
use FILL  FILL_2__2404_
timestamp 1701859473
transform -1 0 2910 0 -1 5470
box -12 -8 32 272
use FILL  FILL_2__2405_
timestamp 1701859473
transform 1 0 2290 0 -1 2870
box -12 -8 32 272
use FILL  FILL_2__2406_
timestamp 1701859473
transform 1 0 2990 0 -1 3390
box -12 -8 32 272
use FILL  FILL_2__2407_
timestamp 1701859473
transform -1 0 3130 0 1 5470
box -12 -8 32 272
use FILL  FILL_2__2408_
timestamp 1701859473
transform 1 0 750 0 -1 2870
box -12 -8 32 272
use FILL  FILL_2__2409_
timestamp 1701859473
transform 1 0 770 0 -1 3910
box -12 -8 32 272
use FILL  FILL_2__2410_
timestamp 1701859473
transform 1 0 1170 0 1 4430
box -12 -8 32 272
use FILL  FILL_2__2411_
timestamp 1701859473
transform -1 0 730 0 -1 4950
box -12 -8 32 272
use FILL  FILL_2__2412_
timestamp 1701859473
transform 1 0 2410 0 -1 5990
box -12 -8 32 272
use FILL  FILL_2__2413_
timestamp 1701859473
transform 1 0 2870 0 1 5470
box -12 -8 32 272
use FILL  FILL_2__2414_
timestamp 1701859473
transform 1 0 4030 0 -1 5470
box -12 -8 32 272
use FILL  FILL_2__2415_
timestamp 1701859473
transform -1 0 3970 0 1 7030
box -12 -8 32 272
use FILL  FILL_2__2416_
timestamp 1701859473
transform 1 0 3930 0 1 4950
box -12 -8 32 272
use FILL  FILL_2__2417_
timestamp 1701859473
transform 1 0 4270 0 -1 5470
box -12 -8 32 272
use FILL  FILL_2__2418_
timestamp 1701859473
transform -1 0 1530 0 -1 4950
box -12 -8 32 272
use FILL  FILL_2__2419_
timestamp 1701859473
transform 1 0 2110 0 1 4430
box -12 -8 32 272
use FILL  FILL_2__2420_
timestamp 1701859473
transform 1 0 3770 0 1 5990
box -12 -8 32 272
use FILL  FILL_2__2421_
timestamp 1701859473
transform -1 0 3550 0 1 5990
box -12 -8 32 272
use FILL  FILL_2__2422_
timestamp 1701859473
transform -1 0 3430 0 -1 5990
box -12 -8 32 272
use FILL  FILL_2__2423_
timestamp 1701859473
transform -1 0 3650 0 -1 5990
box -12 -8 32 272
use FILL  FILL_2__2424_
timestamp 1701859473
transform 1 0 3190 0 -1 5990
box -12 -8 32 272
use FILL  FILL_2__2425_
timestamp 1701859473
transform 1 0 4330 0 1 5990
box -12 -8 32 272
use FILL  FILL_2__2426_
timestamp 1701859473
transform 1 0 3930 0 -1 7030
box -12 -8 32 272
use FILL  FILL_2__2427_
timestamp 1701859473
transform 1 0 4750 0 1 5990
box -12 -8 32 272
use FILL  FILL_2__2428_
timestamp 1701859473
transform 1 0 4510 0 1 5990
box -12 -8 32 272
use FILL  FILL_2__2429_
timestamp 1701859473
transform -1 0 4190 0 -1 6510
box -12 -8 32 272
use FILL  FILL_2__2430_
timestamp 1701859473
transform 1 0 4750 0 1 6510
box -12 -8 32 272
use FILL  FILL_2__2431_
timestamp 1701859473
transform -1 0 4850 0 -1 7030
box -12 -8 32 272
use FILL  FILL_2__2432_
timestamp 1701859473
transform 1 0 5070 0 -1 7030
box -12 -8 32 272
use FILL  FILL_2__2433_
timestamp 1701859473
transform -1 0 4330 0 -1 8070
box -12 -8 32 272
use FILL  FILL_2__2434_
timestamp 1701859473
transform 1 0 4810 0 1 7550
box -12 -8 32 272
use FILL  FILL_2__2435_
timestamp 1701859473
transform 1 0 4150 0 1 7030
box -12 -8 32 272
use FILL  FILL_2__2436_
timestamp 1701859473
transform -1 0 4590 0 -1 7550
box -12 -8 32 272
use FILL  FILL_2__2437_
timestamp 1701859473
transform -1 0 4570 0 -1 8070
box -12 -8 32 272
use FILL  FILL_2__2438_
timestamp 1701859473
transform -1 0 4810 0 -1 8070
box -12 -8 32 272
use FILL  FILL_2__2439_
timestamp 1701859473
transform -1 0 5050 0 -1 8070
box -12 -8 32 272
use FILL  FILL_2__2440_
timestamp 1701859473
transform 1 0 4590 0 1 10150
box -12 -8 32 272
use FILL  FILL_2__2441_
timestamp 1701859473
transform 1 0 3870 0 -1 7550
box -12 -8 32 272
use FILL  FILL_2__2442_
timestamp 1701859473
transform -1 0 4090 0 -1 8070
box -12 -8 32 272
use FILL  FILL_2__2443_
timestamp 1701859473
transform -1 0 3870 0 1 8070
box -12 -8 32 272
use FILL  FILL_2__2444_
timestamp 1701859473
transform 1 0 3610 0 1 8070
box -12 -8 32 272
use FILL  FILL_2__2445_
timestamp 1701859473
transform -1 0 4590 0 1 7550
box -12 -8 32 272
use FILL  FILL_2__2446_
timestamp 1701859473
transform 1 0 4510 0 1 8070
box -12 -8 32 272
use FILL  FILL_2__2447_
timestamp 1701859473
transform 1 0 4250 0 1 9110
box -12 -8 32 272
use FILL  FILL_2__2448_
timestamp 1701859473
transform 1 0 4910 0 1 9110
box -12 -8 32 272
use FILL  FILL_2__2449_
timestamp 1701859473
transform 1 0 5170 0 1 9110
box -12 -8 32 272
use FILL  FILL_2__2450_
timestamp 1701859473
transform 1 0 5410 0 1 9110
box -12 -8 32 272
use FILL  FILL_2__2451_
timestamp 1701859473
transform -1 0 5290 0 -1 9630
box -12 -8 32 272
use FILL  FILL_2__2452_
timestamp 1701859473
transform -1 0 5210 0 -1 10670
box -12 -8 32 272
use FILL  FILL_2__2453_
timestamp 1701859473
transform 1 0 3750 0 -1 10150
box -12 -8 32 272
use FILL  FILL_2__2454_
timestamp 1701859473
transform 1 0 3870 0 1 7550
box -12 -8 32 272
use FILL  FILL_2__2455_
timestamp 1701859473
transform 1 0 3830 0 -1 8070
box -12 -8 32 272
use FILL  FILL_2__2456_
timestamp 1701859473
transform -1 0 3610 0 -1 8070
box -12 -8 32 272
use FILL  FILL_2__2457_
timestamp 1701859473
transform 1 0 3370 0 1 8070
box -12 -8 32 272
use FILL  FILL_2__2458_
timestamp 1701859473
transform -1 0 4310 0 -1 8590
box -12 -8 32 272
use FILL  FILL_2__2459_
timestamp 1701859473
transform -1 0 4470 0 -1 11190
box -12 -8 32 272
use FILL  FILL_2__2460_
timestamp 1701859473
transform 1 0 4110 0 -1 10670
box -12 -8 32 272
use FILL  FILL_2__2461_
timestamp 1701859473
transform 1 0 4290 0 -1 9110
box -12 -8 32 272
use FILL  FILL_2__2462_
timestamp 1701859473
transform -1 0 4550 0 -1 9110
box -12 -8 32 272
use FILL  FILL_2__2463_
timestamp 1701859473
transform -1 0 4790 0 -1 9110
box -12 -8 32 272
use FILL  FILL_2__2464_
timestamp 1701859473
transform -1 0 5030 0 -1 9110
box -12 -8 32 272
use FILL  FILL_2__2465_
timestamp 1701859473
transform -1 0 4890 0 -1 11190
box -12 -8 32 272
use FILL  FILL_2__2466_
timestamp 1701859473
transform -1 0 3970 0 -1 10150
box -12 -8 32 272
use FILL  FILL_2__2467_
timestamp 1701859473
transform -1 0 4070 0 -1 9630
box -12 -8 32 272
use FILL  FILL_2__2468_
timestamp 1701859473
transform -1 0 4330 0 -1 9630
box -12 -8 32 272
use FILL  FILL_2__2469_
timestamp 1701859473
transform -1 0 4190 0 1 9630
box -12 -8 32 272
use FILL  FILL_2__2470_
timestamp 1701859473
transform -1 0 4430 0 1 9630
box -12 -8 32 272
use FILL  FILL_2__2471_
timestamp 1701859473
transform -1 0 5010 0 -1 10670
box -12 -8 32 272
use FILL  FILL_2__2472_
timestamp 1701859473
transform 1 0 3970 0 1 9630
box -12 -8 32 272
use FILL  FILL_2__2473_
timestamp 1701859473
transform 1 0 4530 0 -1 9630
box -12 -8 32 272
use FILL  FILL_2__2474_
timestamp 1701859473
transform -1 0 4810 0 -1 9630
box -12 -8 32 272
use FILL  FILL_2__2475_
timestamp 1701859473
transform 1 0 4650 0 1 9630
box -12 -8 32 272
use FILL  FILL_2__2476_
timestamp 1701859473
transform -1 0 4890 0 1 9630
box -12 -8 32 272
use FILL  FILL_2__2477_
timestamp 1701859473
transform 1 0 4830 0 1 10670
box -12 -8 32 272
use FILL  FILL_2__2478_
timestamp 1701859473
transform 1 0 3070 0 1 5990
box -12 -8 32 272
use FILL  FILL_2__2479_
timestamp 1701859473
transform -1 0 2630 0 1 5990
box -12 -8 32 272
use FILL  FILL_2__2480_
timestamp 1701859473
transform -1 0 2650 0 -1 5990
box -12 -8 32 272
use FILL  FILL_2__2481_
timestamp 1701859473
transform -1 0 2890 0 -1 5990
box -12 -8 32 272
use FILL  FILL_2__2482_
timestamp 1701859473
transform 1 0 1470 0 -1 5990
box -12 -8 32 272
use FILL  FILL_2__2483_
timestamp 1701859473
transform 1 0 2290 0 1 6510
box -12 -8 32 272
use FILL  FILL_2__2484_
timestamp 1701859473
transform -1 0 1910 0 1 6510
box -12 -8 32 272
use FILL  FILL_2__2485_
timestamp 1701859473
transform -1 0 2110 0 1 6510
box -12 -8 32 272
use FILL  FILL_2__2486_
timestamp 1701859473
transform 1 0 2310 0 -1 7030
box -12 -8 32 272
use FILL  FILL_2__2487_
timestamp 1701859473
transform 1 0 2070 0 -1 7030
box -12 -8 32 272
use FILL  FILL_2__2488_
timestamp 1701859473
transform -1 0 1870 0 -1 7030
box -12 -8 32 272
use FILL  FILL_2__2489_
timestamp 1701859473
transform 1 0 1370 0 -1 7030
box -12 -8 32 272
use FILL  FILL_2__2490_
timestamp 1701859473
transform -1 0 970 0 1 5470
box -12 -8 32 272
use FILL  FILL_2__2491_
timestamp 1701859473
transform 1 0 1170 0 1 5470
box -12 -8 32 272
use FILL  FILL_2__2492_
timestamp 1701859473
transform -1 0 2030 0 -1 6510
box -12 -8 32 272
use FILL  FILL_2__2493_
timestamp 1701859473
transform 1 0 1910 0 1 5990
box -12 -8 32 272
use FILL  FILL_2__2494_
timestamp 1701859473
transform -1 0 1470 0 1 5990
box -12 -8 32 272
use FILL  FILL_2__2495_
timestamp 1701859473
transform 1 0 1210 0 1 5990
box -12 -8 32 272
use FILL  FILL_2__2496_
timestamp 1701859473
transform 1 0 1610 0 -1 7030
box -12 -8 32 272
use FILL  FILL_2__2497_
timestamp 1701859473
transform -1 0 1810 0 -1 7550
box -12 -8 32 272
use FILL  FILL_2__2498_
timestamp 1701859473
transform 1 0 750 0 1 8070
box -12 -8 32 272
use FILL  FILL_2__2499_
timestamp 1701859473
transform 1 0 2430 0 1 7550
box -12 -8 32 272
use FILL  FILL_2__2500_
timestamp 1701859473
transform 1 0 1850 0 1 7550
box -12 -8 32 272
use FILL  FILL_2__2501_
timestamp 1701859473
transform 1 0 1630 0 1 7550
box -12 -8 32 272
use FILL  FILL_2__2502_
timestamp 1701859473
transform -1 0 1170 0 1 7550
box -12 -8 32 272
use FILL  FILL_2__2503_
timestamp 1701859473
transform -1 0 1410 0 1 8070
box -12 -8 32 272
use FILL  FILL_2__2504_
timestamp 1701859473
transform -1 0 1830 0 1 8070
box -12 -8 32 272
use FILL  FILL_2__2505_
timestamp 1701859473
transform 1 0 1170 0 1 8070
box -12 -8 32 272
use FILL  FILL_2__2506_
timestamp 1701859473
transform -1 0 1690 0 -1 8070
box -12 -8 32 272
use FILL  FILL_2__2507_
timestamp 1701859473
transform 1 0 1430 0 -1 8070
box -12 -8 32 272
use FILL  FILL_2__2508_
timestamp 1701859473
transform 1 0 950 0 1 8070
box -12 -8 32 272
use FILL  FILL_2__2509_
timestamp 1701859473
transform 1 0 510 0 -1 8590
box -12 -8 32 272
use FILL  FILL_2__2510_
timestamp 1701859473
transform -1 0 1450 0 1 9110
box -12 -8 32 272
use FILL  FILL_2__2511_
timestamp 1701859473
transform -1 0 1390 0 -1 9630
box -12 -8 32 272
use FILL  FILL_2__2512_
timestamp 1701859473
transform 1 0 950 0 -1 9630
box -12 -8 32 272
use FILL  FILL_2__2513_
timestamp 1701859473
transform -1 0 950 0 1 8590
box -12 -8 32 272
use FILL  FILL_2__2514_
timestamp 1701859473
transform 1 0 2030 0 -1 8590
box -12 -8 32 272
use FILL  FILL_2__2515_
timestamp 1701859473
transform 1 0 1150 0 -1 9110
box -12 -8 32 272
use FILL  FILL_2__2516_
timestamp 1701859473
transform -1 0 990 0 1 9110
box -12 -8 32 272
use FILL  FILL_2__2517_
timestamp 1701859473
transform -1 0 750 0 1 9110
box -12 -8 32 272
use FILL  FILL_2__2518_
timestamp 1701859473
transform 1 0 1610 0 -1 9630
box -12 -8 32 272
use FILL  FILL_2__2519_
timestamp 1701859473
transform 1 0 1710 0 1 9630
box -12 -8 32 272
use FILL  FILL_2__2520_
timestamp 1701859473
transform -1 0 2550 0 -1 9110
box -12 -8 32 272
use FILL  FILL_2__2521_
timestamp 1701859473
transform 1 0 2290 0 -1 9110
box -12 -8 32 272
use FILL  FILL_2__2522_
timestamp 1701859473
transform -1 0 1910 0 1 9630
box -12 -8 32 272
use FILL  FILL_2__2523_
timestamp 1701859473
transform -1 0 2130 0 1 9630
box -12 -8 32 272
use FILL  FILL_2__2524_
timestamp 1701859473
transform -1 0 1870 0 -1 9110
box -12 -8 32 272
use FILL  FILL_2__2525_
timestamp 1701859473
transform 1 0 750 0 -1 8590
box -12 -8 32 272
use FILL  FILL_2__2526_
timestamp 1701859473
transform -1 0 1650 0 -1 8590
box -12 -8 32 272
use FILL  FILL_2__2527_
timestamp 1701859473
transform -1 0 1190 0 -1 8590
box -12 -8 32 272
use FILL  FILL_2__2528_
timestamp 1701859473
transform -1 0 970 0 -1 8590
box -12 -8 32 272
use FILL  FILL_2__2529_
timestamp 1701859473
transform -1 0 1210 0 1 9110
box -12 -8 32 272
use FILL  FILL_2__2530_
timestamp 1701859473
transform -1 0 7470 0 -1 6510
box -12 -8 32 272
use FILL  FILL_2__2531_
timestamp 1701859473
transform 1 0 7890 0 1 7550
box -12 -8 32 272
use FILL  FILL_2__2532_
timestamp 1701859473
transform -1 0 9790 0 1 2870
box -12 -8 32 272
use FILL  FILL_2__2533_
timestamp 1701859473
transform -1 0 8870 0 1 4430
box -12 -8 32 272
use FILL  FILL_2__2534_
timestamp 1701859473
transform -1 0 9270 0 -1 5470
box -12 -8 32 272
use FILL  FILL_2__2535_
timestamp 1701859473
transform 1 0 50 0 -1 4950
box -12 -8 32 272
use FILL  FILL_2__2536_
timestamp 1701859473
transform 1 0 610 0 1 4950
box -12 -8 32 272
use FILL  FILL_2__2537_
timestamp 1701859473
transform 1 0 750 0 1 3390
box -12 -8 32 272
use FILL  FILL_2__2538_
timestamp 1701859473
transform -1 0 310 0 -1 3910
box -12 -8 32 272
use FILL  FILL_2__2539_
timestamp 1701859473
transform -1 0 70 0 1 4950
box -12 -8 32 272
use FILL  FILL_2__2540_
timestamp 1701859473
transform 1 0 3010 0 1 2350
box -12 -8 32 272
use FILL  FILL_2__2541_
timestamp 1701859473
transform -1 0 3270 0 1 2870
box -12 -8 32 272
use FILL  FILL_2__2542_
timestamp 1701859473
transform -1 0 2270 0 -1 6510
box -12 -8 32 272
use FILL  FILL_2__2543_
timestamp 1701859473
transform 1 0 830 0 1 4950
box -12 -8 32 272
use FILL  FILL_2__2544_
timestamp 1701859473
transform 1 0 1390 0 1 4430
box -12 -8 32 272
use FILL  FILL_2__2545_
timestamp 1701859473
transform 1 0 1250 0 -1 5470
box -12 -8 32 272
use FILL  FILL_2__2546_
timestamp 1701859473
transform -1 0 1990 0 -1 5470
box -12 -8 32 272
use FILL  FILL_2__2547_
timestamp 1701859473
transform 1 0 1930 0 -1 4430
box -12 -8 32 272
use FILL  FILL_2__2548_
timestamp 1701859473
transform 1 0 1050 0 1 4950
box -12 -8 32 272
use FILL  FILL_2__2549_
timestamp 1701859473
transform 1 0 1270 0 1 4950
box -12 -8 32 272
use FILL  FILL_2__2550_
timestamp 1701859473
transform -1 0 1750 0 -1 5470
box -12 -8 32 272
use FILL  FILL_2__2551_
timestamp 1701859473
transform 1 0 2530 0 -1 9630
box -12 -8 32 272
use FILL  FILL_2__2552_
timestamp 1701859473
transform 1 0 3370 0 -1 5470
box -12 -8 32 272
use FILL  FILL_2__2553_
timestamp 1701859473
transform -1 0 2750 0 -1 6510
box -12 -8 32 272
use FILL  FILL_2__2554_
timestamp 1701859473
transform -1 0 3210 0 1 6510
box -12 -8 32 272
use FILL  FILL_2__2555_
timestamp 1701859473
transform -1 0 3450 0 1 6510
box -12 -8 32 272
use FILL  FILL_2__2556_
timestamp 1701859473
transform -1 0 2770 0 1 6510
box -12 -8 32 272
use FILL  FILL_2__2557_
timestamp 1701859473
transform 1 0 2470 0 -1 6510
box -12 -8 32 272
use FILL  FILL_2__2558_
timestamp 1701859473
transform 1 0 3210 0 -1 7550
box -12 -8 32 272
use FILL  FILL_2__2559_
timestamp 1701859473
transform 1 0 3410 0 -1 7550
box -12 -8 32 272
use FILL  FILL_2__2560_
timestamp 1701859473
transform -1 0 3470 0 1 7030
box -12 -8 32 272
use FILL  FILL_2__2561_
timestamp 1701859473
transform -1 0 1490 0 1 4950
box -12 -8 32 272
use FILL  FILL_2__2562_
timestamp 1701859473
transform 1 0 3210 0 1 7030
box -12 -8 32 272
use FILL  FILL_2__2563_
timestamp 1701859473
transform 1 0 3770 0 1 5470
box -12 -8 32 272
use FILL  FILL_2__2564_
timestamp 1701859473
transform -1 0 3650 0 1 6510
box -12 -8 32 272
use FILL  FILL_2__2565_
timestamp 1701859473
transform 1 0 3710 0 1 7030
box -12 -8 32 272
use FILL  FILL_2__2566_
timestamp 1701859473
transform 1 0 3170 0 1 7550
box -12 -8 32 272
use FILL  FILL_2__2567_
timestamp 1701859473
transform 1 0 3130 0 -1 8070
box -12 -8 32 272
use FILL  FILL_2__2568_
timestamp 1701859473
transform -1 0 2950 0 -1 8590
box -12 -8 32 272
use FILL  FILL_2__2569_
timestamp 1701859473
transform 1 0 2710 0 -1 8590
box -12 -8 32 272
use FILL  FILL_2__2570_
timestamp 1701859473
transform 1 0 2890 0 -1 8070
box -12 -8 32 272
use FILL  FILL_2__2571_
timestamp 1701859473
transform -1 0 3850 0 -1 9630
box -12 -8 32 272
use FILL  FILL_2__2572_
timestamp 1701859473
transform -1 0 3870 0 -1 5990
box -12 -8 32 272
use FILL  FILL_2__2573_
timestamp 1701859473
transform -1 0 3730 0 -1 7030
box -12 -8 32 272
use FILL  FILL_2__2574_
timestamp 1701859473
transform 1 0 3450 0 -1 6510
box -12 -8 32 272
use FILL  FILL_2__2575_
timestamp 1701859473
transform 1 0 3350 0 -1 8070
box -12 -8 32 272
use FILL  FILL_2__2576_
timestamp 1701859473
transform -1 0 3390 0 -1 8590
box -12 -8 32 272
use FILL  FILL_2__2577_
timestamp 1701859473
transform 1 0 3270 0 1 9110
box -12 -8 32 272
use FILL  FILL_2__2578_
timestamp 1701859473
transform 1 0 3770 0 1 9110
box -12 -8 32 272
use FILL  FILL_2__2579_
timestamp 1701859473
transform -1 0 2750 0 -1 9630
box -12 -8 32 272
use FILL  FILL_2__2580_
timestamp 1701859473
transform -1 0 4110 0 -1 9110
box -12 -8 32 272
use FILL  FILL_2__2581_
timestamp 1701859473
transform -1 0 4030 0 1 9110
box -12 -8 32 272
use FILL  FILL_2__2582_
timestamp 1701859473
transform 1 0 3530 0 1 9110
box -12 -8 32 272
use FILL  FILL_2__2583_
timestamp 1701859473
transform 1 0 3030 0 1 9110
box -12 -8 32 272
use FILL  FILL_2__2584_
timestamp 1701859473
transform 1 0 2790 0 1 9110
box -12 -8 32 272
use FILL  FILL_2__2585_
timestamp 1701859473
transform 1 0 3890 0 -1 9110
box -12 -8 32 272
use FILL  FILL_2__2586_
timestamp 1701859473
transform 1 0 3050 0 1 9630
box -12 -8 32 272
use FILL  FILL_2__2587_
timestamp 1701859473
transform 1 0 3630 0 -1 9110
box -12 -8 32 272
use FILL  FILL_2__2588_
timestamp 1701859473
transform 1 0 3230 0 1 8590
box -12 -8 32 272
use FILL  FILL_2__2589_
timestamp 1701859473
transform 1 0 3070 0 -1 10150
box -12 -8 32 272
use FILL  FILL_2__2590_
timestamp 1701859473
transform 1 0 2810 0 -1 10150
box -12 -8 32 272
use FILL  FILL_2__2591_
timestamp 1701859473
transform -1 0 3570 0 -1 11190
box -12 -8 32 272
use FILL  FILL_2__2592_
timestamp 1701859473
transform -1 0 3630 0 -1 9630
box -12 -8 32 272
use FILL  FILL_2__2593_
timestamp 1701859473
transform -1 0 3150 0 -1 9630
box -12 -8 32 272
use FILL  FILL_2__2594_
timestamp 1701859473
transform -1 0 3310 0 -1 10150
box -12 -8 32 272
use FILL  FILL_2__2595_
timestamp 1701859473
transform 1 0 3030 0 -1 11190
box -12 -8 32 272
use FILL  FILL_2__2596_
timestamp 1701859473
transform 1 0 3310 0 -1 11190
box -12 -8 32 272
use FILL  FILL_2__2597_
timestamp 1701859473
transform 1 0 2770 0 -1 10670
box -12 -8 32 272
use FILL  FILL_2__2598_
timestamp 1701859473
transform -1 0 3510 0 1 9630
box -12 -8 32 272
use FILL  FILL_2__2599_
timestamp 1701859473
transform -1 0 3290 0 1 9630
box -12 -8 32 272
use FILL  FILL_2__2600_
timestamp 1701859473
transform -1 0 3010 0 1 10150
box -12 -8 32 272
use FILL  FILL_2__2601_
timestamp 1701859473
transform 1 0 2970 0 -1 10670
box -12 -8 32 272
use FILL  FILL_2__2602_
timestamp 1701859473
transform -1 0 3230 0 -1 10670
box -12 -8 32 272
use FILL  FILL_2__2603_
timestamp 1701859473
transform 1 0 3430 0 -1 10670
box -12 -8 32 272
use FILL  FILL_2__2604_
timestamp 1701859473
transform 1 0 3230 0 1 10150
box -12 -8 32 272
use FILL  FILL_2__2605_
timestamp 1701859473
transform 1 0 2350 0 1 10670
box -12 -8 32 272
use FILL  FILL_2__2606_
timestamp 1701859473
transform 1 0 2550 0 1 10670
box -12 -8 32 272
use FILL  FILL_2__2607_
timestamp 1701859473
transform -1 0 2790 0 1 10670
box -12 -8 32 272
use FILL  FILL_2__2608_
timestamp 1701859473
transform -1 0 3750 0 1 9630
box -12 -8 32 272
use FILL  FILL_2__2609_
timestamp 1701859473
transform -1 0 2370 0 1 9630
box -12 -8 32 272
use FILL  FILL_2__2610_
timestamp 1701859473
transform -1 0 2590 0 -1 10150
box -12 -8 32 272
use FILL  FILL_2__2611_
timestamp 1701859473
transform -1 0 2310 0 -1 10670
box -12 -8 32 272
use FILL  FILL_2__2612_
timestamp 1701859473
transform 1 0 2530 0 -1 10670
box -12 -8 32 272
use FILL  FILL_2__2613_
timestamp 1701859473
transform 1 0 1850 0 1 10670
box -12 -8 32 272
use FILL  FILL_2__2614_
timestamp 1701859473
transform 1 0 1850 0 -1 10670
box -12 -8 32 272
use FILL  FILL_2__2615_
timestamp 1701859473
transform -1 0 2370 0 -1 11190
box -12 -8 32 272
use FILL  FILL_2__2616_
timestamp 1701859473
transform -1 0 3390 0 -1 9630
box -12 -8 32 272
use FILL  FILL_2__2617_
timestamp 1701859473
transform 1 0 2290 0 -1 9630
box -12 -8 32 272
use FILL  FILL_2__2618_
timestamp 1701859473
transform -1 0 2570 0 1 10150
box -12 -8 32 272
use FILL  FILL_2__2619_
timestamp 1701859473
transform 1 0 2070 0 1 10670
box -12 -8 32 272
use FILL  FILL_2__2620_
timestamp 1701859473
transform 1 0 2110 0 -1 11190
box -12 -8 32 272
use FILL  FILL_2__2621_
timestamp 1701859473
transform -1 0 1390 0 1 5470
box -12 -8 32 272
use FILL  FILL_2__2622_
timestamp 1701859473
transform -1 0 1230 0 -1 5990
box -12 -8 32 272
use FILL  FILL_2__2623_
timestamp 1701859473
transform 1 0 2450 0 -1 5470
box -12 -8 32 272
use FILL  FILL_2__2624_
timestamp 1701859473
transform -1 0 2410 0 1 5470
box -12 -8 32 272
use FILL  FILL_2__2625_
timestamp 1701859473
transform 1 0 2210 0 -1 5470
box -12 -8 32 272
use FILL  FILL_2__2626_
timestamp 1701859473
transform -1 0 950 0 -1 5470
box -12 -8 32 272
use FILL  FILL_2__2627_
timestamp 1701859473
transform -1 0 1470 0 1 3910
box -12 -8 32 272
use FILL  FILL_2__2628_
timestamp 1701859473
transform 1 0 1150 0 1 3910
box -12 -8 32 272
use FILL  FILL_2__2629_
timestamp 1701859473
transform -1 0 750 0 -1 5470
box -12 -8 32 272
use FILL  FILL_2__2630_
timestamp 1701859473
transform 1 0 730 0 -1 5990
box -12 -8 32 272
use FILL  FILL_2__2631_
timestamp 1701859473
transform -1 0 730 0 1 5990
box -12 -8 32 272
use FILL  FILL_2__2632_
timestamp 1701859473
transform 1 0 2110 0 1 10150
box -12 -8 32 272
use FILL  FILL_2__2633_
timestamp 1701859473
transform -1 0 2350 0 1 10150
box -12 -8 32 272
use FILL  FILL_2__2634_
timestamp 1701859473
transform 1 0 2310 0 -1 10150
box -12 -8 32 272
use FILL  FILL_2__2635_
timestamp 1701859473
transform 1 0 2090 0 -1 10150
box -12 -8 32 272
use FILL  FILL_2__2636_
timestamp 1701859473
transform -1 0 730 0 -1 10150
box -12 -8 32 272
use FILL  FILL_2__2637_
timestamp 1701859473
transform -1 0 530 0 1 6510
box -12 -8 32 272
use FILL  FILL_2__2638_
timestamp 1701859473
transform -1 0 310 0 1 6510
box -12 -8 32 272
use FILL  FILL_2__2639_
timestamp 1701859473
transform -1 0 290 0 -1 6510
box -12 -8 32 272
use FILL  FILL_2__2640_
timestamp 1701859473
transform -1 0 290 0 1 5990
box -12 -8 32 272
use FILL  FILL_2__2641_
timestamp 1701859473
transform 1 0 50 0 -1 7550
box -12 -8 32 272
use FILL  FILL_2__2642_
timestamp 1701859473
transform -1 0 390 0 1 4950
box -12 -8 32 272
use FILL  FILL_2__2643_
timestamp 1701859473
transform -1 0 2530 0 1 6510
box -12 -8 32 272
use FILL  FILL_2__2644_
timestamp 1701859473
transform 1 0 2570 0 -1 7030
box -12 -8 32 272
use FILL  FILL_2__2645_
timestamp 1701859473
transform 1 0 2750 0 1 7030
box -12 -8 32 272
use FILL  FILL_2__2646_
timestamp 1701859473
transform 1 0 2050 0 1 7030
box -12 -8 32 272
use FILL  FILL_2__2647_
timestamp 1701859473
transform 1 0 730 0 1 7550
box -12 -8 32 272
use FILL  FILL_2__2648_
timestamp 1701859473
transform 1 0 270 0 1 7550
box -12 -8 32 272
use FILL  FILL_2__2649_
timestamp 1701859473
transform 1 0 250 0 -1 7550
box -12 -8 32 272
use FILL  FILL_2__2650_
timestamp 1701859473
transform -1 0 730 0 -1 7550
box -12 -8 32 272
use FILL  FILL_2__2651_
timestamp 1701859473
transform 1 0 470 0 -1 7550
box -12 -8 32 272
use FILL  FILL_2__2652_
timestamp 1701859473
transform 1 0 470 0 1 7030
box -12 -8 32 272
use FILL  FILL_2__2653_
timestamp 1701859473
transform 1 0 50 0 1 7550
box -12 -8 32 272
use FILL  FILL_2__2654_
timestamp 1701859473
transform -1 0 530 0 1 7550
box -12 -8 32 272
use FILL  FILL_2__2655_
timestamp 1701859473
transform 1 0 1850 0 1 7030
box -12 -8 32 272
use FILL  FILL_2__2656_
timestamp 1701859473
transform 1 0 1490 0 -1 5470
box -12 -8 32 272
use FILL  FILL_2__2657_
timestamp 1701859473
transform -1 0 1690 0 1 5990
box -12 -8 32 272
use FILL  FILL_2__2658_
timestamp 1701859473
transform -1 0 2170 0 1 5470
box -12 -8 32 272
use FILL  FILL_2__2659_
timestamp 1701859473
transform 1 0 1930 0 -1 5990
box -12 -8 32 272
use FILL  FILL_2__2660_
timestamp 1701859473
transform -1 0 1930 0 1 5470
box -12 -8 32 272
use FILL  FILL_2__2661_
timestamp 1701859473
transform -1 0 1610 0 1 5470
box -12 -8 32 272
use FILL  FILL_2__2662_
timestamp 1701859473
transform 1 0 710 0 1 5470
box -12 -8 32 272
use FILL  FILL_2__2663_
timestamp 1701859473
transform -1 0 990 0 -1 5990
box -12 -8 32 272
use FILL  FILL_2__2664_
timestamp 1701859473
transform 1 0 710 0 -1 7030
box -12 -8 32 272
use FILL  FILL_2__2665_
timestamp 1701859473
transform 1 0 1170 0 -1 7030
box -12 -8 32 272
use FILL  FILL_2__2666_
timestamp 1701859473
transform 1 0 1370 0 1 7030
box -12 -8 32 272
use FILL  FILL_2__2667_
timestamp 1701859473
transform 1 0 910 0 -1 7030
box -12 -8 32 272
use FILL  FILL_2__2668_
timestamp 1701859473
transform -1 0 2710 0 1 7550
box -12 -8 32 272
use FILL  FILL_2__2669_
timestamp 1701859473
transform 1 0 2650 0 -1 8070
box -12 -8 32 272
use FILL  FILL_2__2670_
timestamp 1701859473
transform 1 0 1910 0 -1 8070
box -12 -8 32 272
use FILL  FILL_2__2671_
timestamp 1701859473
transform -1 0 1410 0 1 7550
box -12 -8 32 272
use FILL  FILL_2__2672_
timestamp 1701859473
transform 1 0 1130 0 -1 7550
box -12 -8 32 272
use FILL  FILL_2__2673_
timestamp 1701859473
transform -1 0 1330 0 -1 7550
box -12 -8 32 272
use FILL  FILL_2__2674_
timestamp 1701859473
transform 1 0 1610 0 1 7030
box -12 -8 32 272
use FILL  FILL_2__2675_
timestamp 1701859473
transform 1 0 1550 0 -1 7550
box -12 -8 32 272
use FILL  FILL_2__2676_
timestamp 1701859473
transform -1 0 1990 0 -1 7550
box -12 -8 32 272
use FILL  FILL_2__2677_
timestamp 1701859473
transform 1 0 2390 0 -1 8070
box -12 -8 32 272
use FILL  FILL_2__2678_
timestamp 1701859473
transform -1 0 2170 0 -1 8070
box -12 -8 32 272
use FILL  FILL_2__2679_
timestamp 1701859473
transform -1 0 1610 0 1 8070
box -12 -8 32 272
use FILL  FILL_2__2680_
timestamp 1701859473
transform -1 0 290 0 -1 8590
box -12 -8 32 272
use FILL  FILL_2__2681_
timestamp 1701859473
transform 1 0 910 0 -1 7550
box -12 -8 32 272
use FILL  FILL_2__2682_
timestamp 1701859473
transform -1 0 290 0 -1 8070
box -12 -8 32 272
use FILL  FILL_2__2683_
timestamp 1701859473
transform -1 0 70 0 -1 9630
box -12 -8 32 272
use FILL  FILL_2__2684_
timestamp 1701859473
transform -1 0 70 0 1 10150
box -12 -8 32 272
use FILL  FILL_2__2685_
timestamp 1701859473
transform 1 0 950 0 1 5990
box -12 -8 32 272
use FILL  FILL_2__2686_
timestamp 1701859473
transform 1 0 930 0 1 7550
box -12 -8 32 272
use FILL  FILL_2__2687_
timestamp 1701859473
transform -1 0 930 0 -1 10150
box -12 -8 32 272
use FILL  FILL_2__2688_
timestamp 1701859473
transform 1 0 50 0 -1 10150
box -12 -8 32 272
use FILL  FILL_2__2689_
timestamp 1701859473
transform 1 0 270 0 -1 9630
box -12 -8 32 272
use FILL  FILL_2__2690_
timestamp 1701859473
transform 1 0 270 0 1 9110
box -12 -8 32 272
use FILL  FILL_2__2691_
timestamp 1701859473
transform 1 0 2730 0 1 8590
box -12 -8 32 272
use FILL  FILL_2__2692_
timestamp 1701859473
transform 1 0 2490 0 1 8590
box -12 -8 32 272
use FILL  FILL_2__2693_
timestamp 1701859473
transform -1 0 1150 0 -1 9630
box -12 -8 32 272
use FILL  FILL_2__2694_
timestamp 1701859473
transform 1 0 730 0 -1 9630
box -12 -8 32 272
use FILL  FILL_2__2695_
timestamp 1701859473
transform 1 0 50 0 1 9630
box -12 -8 32 272
use FILL  FILL_2__2696_
timestamp 1701859473
transform -1 0 530 0 -1 10150
box -12 -8 32 272
use FILL  FILL_2__2697_
timestamp 1701859473
transform 1 0 270 0 -1 10150
box -12 -8 32 272
use FILL  FILL_2__2698_
timestamp 1701859473
transform 1 0 290 0 1 9630
box -12 -8 32 272
use FILL  FILL_2__2699_
timestamp 1701859473
transform 1 0 510 0 -1 9630
box -12 -8 32 272
use FILL  FILL_2__2700_
timestamp 1701859473
transform 1 0 530 0 1 9630
box -12 -8 32 272
use FILL  FILL_2__2701_
timestamp 1701859473
transform -1 0 750 0 -1 10670
box -12 -8 32 272
use FILL  FILL_2__2702_
timestamp 1701859473
transform 1 0 3470 0 1 8590
box -12 -8 32 272
use FILL  FILL_2__2703_
timestamp 1701859473
transform -1 0 3010 0 1 8590
box -12 -8 32 272
use FILL  FILL_2__2704_
timestamp 1701859473
transform -1 0 1490 0 1 9630
box -12 -8 32 272
use FILL  FILL_2__2705_
timestamp 1701859473
transform 1 0 1230 0 1 9630
box -12 -8 32 272
use FILL  FILL_2__2706_
timestamp 1701859473
transform 1 0 250 0 1 10150
box -12 -8 32 272
use FILL  FILL_2__2707_
timestamp 1701859473
transform -1 0 490 0 1 10150
box -12 -8 32 272
use FILL  FILL_2__2708_
timestamp 1701859473
transform 1 0 690 0 1 10150
box -12 -8 32 272
use FILL  FILL_2__2709_
timestamp 1701859473
transform -1 0 510 0 -1 10670
box -12 -8 32 272
use FILL  FILL_2__2710_
timestamp 1701859473
transform 1 0 1690 0 1 10150
box -12 -8 32 272
use FILL  FILL_2__2711_
timestamp 1701859473
transform 1 0 2230 0 1 8590
box -12 -8 32 272
use FILL  FILL_2__2712_
timestamp 1701859473
transform -1 0 2010 0 1 8590
box -12 -8 32 272
use FILL  FILL_2__2713_
timestamp 1701859473
transform -1 0 1870 0 -1 9630
box -12 -8 32 272
use FILL  FILL_2__2714_
timestamp 1701859473
transform 1 0 1630 0 -1 10150
box -12 -8 32 272
use FILL  FILL_2__2715_
timestamp 1701859473
transform 1 0 950 0 1 10150
box -12 -8 32 272
use FILL  FILL_2__2716_
timestamp 1701859473
transform 1 0 1190 0 1 10150
box -12 -8 32 272
use FILL  FILL_2__2717_
timestamp 1701859473
transform 1 0 1450 0 1 10150
box -12 -8 32 272
use FILL  FILL_2__2718_
timestamp 1701859473
transform -1 0 10030 0 1 4950
box -12 -8 32 272
use FILL  FILL_2__2719_
timestamp 1701859473
transform -1 0 9790 0 1 4950
box -12 -8 32 272
use FILL  FILL_2__2720_
timestamp 1701859473
transform -1 0 4570 0 1 4950
box -12 -8 32 272
use FILL  FILL_2__2721_
timestamp 1701859473
transform -1 0 7330 0 -1 2350
box -12 -8 32 272
use FILL  FILL_2__2722_
timestamp 1701859473
transform 1 0 9970 0 -1 790
box -12 -8 32 272
use FILL  FILL_2__2723_
timestamp 1701859473
transform -1 0 7090 0 1 1830
box -12 -8 32 272
use FILL  FILL_2__2724_
timestamp 1701859473
transform -1 0 7090 0 -1 2350
box -12 -8 32 272
use FILL  FILL_2__2725_
timestamp 1701859473
transform 1 0 6950 0 1 3390
box -12 -8 32 272
use FILL  FILL_2__2726_
timestamp 1701859473
transform -1 0 7190 0 1 3390
box -12 -8 32 272
use FILL  FILL_2__2727_
timestamp 1701859473
transform -1 0 5410 0 1 3390
box -12 -8 32 272
use FILL  FILL_2__2728_
timestamp 1701859473
transform -1 0 5630 0 1 3390
box -12 -8 32 272
use FILL  FILL_2__2729_
timestamp 1701859473
transform -1 0 6730 0 -1 3910
box -12 -8 32 272
use FILL  FILL_2__2730_
timestamp 1701859473
transform 1 0 8230 0 -1 3910
box -12 -8 32 272
use FILL  FILL_2__2731_
timestamp 1701859473
transform 1 0 9250 0 1 1830
box -12 -8 32 272
use FILL  FILL_2__2732_
timestamp 1701859473
transform 1 0 7690 0 1 1830
box -12 -8 32 272
use FILL  FILL_2__2733_
timestamp 1701859473
transform 1 0 8570 0 1 2350
box -12 -8 32 272
use FILL  FILL_2__2734_
timestamp 1701859473
transform 1 0 7150 0 -1 5470
box -12 -8 32 272
use FILL  FILL_2__2735_
timestamp 1701859473
transform 1 0 7230 0 -1 2870
box -12 -8 32 272
use FILL  FILL_2__2736_
timestamp 1701859473
transform -1 0 7510 0 1 1310
box -12 -8 32 272
use FILL  FILL_2__2737_
timestamp 1701859473
transform 1 0 8570 0 1 1830
box -12 -8 32 272
use FILL  FILL_2__2738_
timestamp 1701859473
transform -1 0 7950 0 -1 2870
box -12 -8 32 272
use FILL  FILL_2__2739_
timestamp 1701859473
transform -1 0 7770 0 1 2870
box -12 -8 32 272
use FILL  FILL_2__2740_
timestamp 1701859473
transform -1 0 6550 0 -1 1830
box -12 -8 32 272
use FILL  FILL_2__2741_
timestamp 1701859473
transform 1 0 6750 0 -1 1830
box -12 -8 32 272
use FILL  FILL_2__2742_
timestamp 1701859473
transform -1 0 8190 0 -1 2870
box -12 -8 32 272
use FILL  FILL_2__2743_
timestamp 1701859473
transform -1 0 8210 0 1 2870
box -12 -8 32 272
use FILL  FILL_2__2744_
timestamp 1701859473
transform -1 0 7330 0 -1 270
box -12 -8 32 272
use FILL  FILL_2__2745_
timestamp 1701859473
transform -1 0 7290 0 1 1830
box -12 -8 32 272
use FILL  FILL_2__2746_
timestamp 1701859473
transform 1 0 7950 0 1 2870
box -12 -8 32 272
use FILL  FILL_2__2747_
timestamp 1701859473
transform -1 0 7750 0 -1 2350
box -12 -8 32 272
use FILL  FILL_2__2748_
timestamp 1701859473
transform 1 0 7930 0 -1 2350
box -12 -8 32 272
use FILL  FILL_2__2749_
timestamp 1701859473
transform 1 0 5890 0 1 1830
box -12 -8 32 272
use FILL  FILL_2__2750_
timestamp 1701859473
transform -1 0 6650 0 -1 1310
box -12 -8 32 272
use FILL  FILL_2__2751_
timestamp 1701859473
transform -1 0 6370 0 1 1830
box -12 -8 32 272
use FILL  FILL_2__2752_
timestamp 1701859473
transform -1 0 7730 0 1 2350
box -12 -8 32 272
use FILL  FILL_2__2753_
timestamp 1701859473
transform -1 0 7470 0 1 2350
box -12 -8 32 272
use FILL  FILL_2__2754_
timestamp 1701859473
transform 1 0 8810 0 -1 4950
box -12 -8 32 272
use FILL  FILL_2__2755_
timestamp 1701859473
transform 1 0 9710 0 1 790
box -12 -8 32 272
use FILL  FILL_2__2756_
timestamp 1701859473
transform -1 0 9950 0 1 790
box -12 -8 32 272
use FILL  FILL_2__2757_
timestamp 1701859473
transform 1 0 10650 0 -1 2870
box -12 -8 32 272
use FILL  FILL_2__2758_
timestamp 1701859473
transform -1 0 9150 0 -1 2870
box -12 -8 32 272
use FILL  FILL_2__2759_
timestamp 1701859473
transform 1 0 9070 0 1 4430
box -12 -8 32 272
use FILL  FILL_2__2760_
timestamp 1701859473
transform 1 0 10410 0 -1 790
box -12 -8 32 272
use FILL  FILL_2__2761_
timestamp 1701859473
transform 1 0 10170 0 -1 790
box -12 -8 32 272
use FILL  FILL_2__2762_
timestamp 1701859473
transform -1 0 10850 0 -1 1830
box -12 -8 32 272
use FILL  FILL_2__2763_
timestamp 1701859473
transform 1 0 6590 0 1 1830
box -12 -8 32 272
use FILL  FILL_2__2764_
timestamp 1701859473
transform -1 0 6850 0 1 1830
box -12 -8 32 272
use FILL  FILL_2__2765_
timestamp 1701859473
transform -1 0 10150 0 1 1830
box -12 -8 32 272
use FILL  FILL_2__2766_
timestamp 1701859473
transform -1 0 9970 0 -1 1830
box -12 -8 32 272
use FILL  FILL_2__2767_
timestamp 1701859473
transform -1 0 10390 0 -1 1830
box -12 -8 32 272
use FILL  FILL_2__2768_
timestamp 1701859473
transform -1 0 10370 0 1 1830
box -12 -8 32 272
use FILL  FILL_2__2769_
timestamp 1701859473
transform -1 0 10830 0 1 2350
box -12 -8 32 272
use FILL  FILL_2__2770_
timestamp 1701859473
transform -1 0 10610 0 -1 1830
box -12 -8 32 272
use FILL  FILL_2__2771_
timestamp 1701859473
transform 1 0 11030 0 1 2350
box -12 -8 32 272
use FILL  FILL_2__2772_
timestamp 1701859473
transform -1 0 10690 0 1 4950
box -12 -8 32 272
use FILL  FILL_2__2773_
timestamp 1701859473
transform 1 0 10430 0 -1 3910
box -12 -8 32 272
use FILL  FILL_2__2774_
timestamp 1701859473
transform -1 0 10730 0 -1 2350
box -12 -8 32 272
use FILL  FILL_2__2775_
timestamp 1701859473
transform -1 0 9090 0 -1 1310
box -12 -8 32 272
use FILL  FILL_2__2776_
timestamp 1701859473
transform 1 0 10630 0 -1 790
box -12 -8 32 272
use FILL  FILL_2__2777_
timestamp 1701859473
transform -1 0 8390 0 -1 270
box -12 -8 32 272
use FILL  FILL_2__2778_
timestamp 1701859473
transform 1 0 10930 0 1 270
box -12 -8 32 272
use FILL  FILL_2__2779_
timestamp 1701859473
transform 1 0 9010 0 -1 1830
box -12 -8 32 272
use FILL  FILL_2__2780_
timestamp 1701859473
transform -1 0 10030 0 1 1310
box -12 -8 32 272
use FILL  FILL_2__2781_
timestamp 1701859473
transform 1 0 10170 0 -1 1310
box -12 -8 32 272
use FILL  FILL_2__2782_
timestamp 1701859473
transform 1 0 8790 0 1 1830
box -12 -8 32 272
use FILL  FILL_2__2783_
timestamp 1701859473
transform 1 0 8350 0 -1 1310
box -12 -8 32 272
use FILL  FILL_2__2784_
timestamp 1701859473
transform 1 0 8590 0 -1 1310
box -12 -8 32 272
use FILL  FILL_2__2785_
timestamp 1701859473
transform 1 0 8810 0 -1 1830
box -12 -8 32 272
use FILL  FILL_2__2786_
timestamp 1701859473
transform -1 0 9290 0 -1 1310
box -12 -8 32 272
use FILL  FILL_2__2787_
timestamp 1701859473
transform -1 0 9490 0 -1 1830
box -12 -8 32 272
use FILL  FILL_2__2788_
timestamp 1701859473
transform 1 0 10170 0 -1 1830
box -12 -8 32 272
use FILL  FILL_2__2789_
timestamp 1701859473
transform 1 0 10250 0 1 1310
box -12 -8 32 272
use FILL  FILL_2__2790_
timestamp 1701859473
transform -1 0 10050 0 -1 2350
box -12 -8 32 272
use FILL  FILL_2__2791_
timestamp 1701859473
transform 1 0 9810 0 -1 2350
box -12 -8 32 272
use FILL  FILL_2__2792_
timestamp 1701859473
transform -1 0 10270 0 -1 2350
box -12 -8 32 272
use FILL  FILL_2__2793_
timestamp 1701859473
transform -1 0 10510 0 -1 2350
box -12 -8 32 272
use FILL  FILL_2__2794_
timestamp 1701859473
transform -1 0 10930 0 -1 2350
box -12 -8 32 272
use FILL  FILL_2__2795_
timestamp 1701859473
transform -1 0 10890 0 -1 2870
box -12 -8 32 272
use FILL  FILL_2__2796_
timestamp 1701859473
transform -1 0 10230 0 -1 2870
box -12 -8 32 272
use FILL  FILL_2__2797_
timestamp 1701859473
transform -1 0 9730 0 -1 1830
box -12 -8 32 272
use FILL  FILL_2__2798_
timestamp 1701859473
transform -1 0 10610 0 1 2350
box -12 -8 32 272
use FILL  FILL_2__2799_
timestamp 1701859473
transform 1 0 10390 0 -1 2870
box -12 -8 32 272
use FILL  FILL_2__2800_
timestamp 1701859473
transform -1 0 10410 0 -1 4430
box -12 -8 32 272
use FILL  FILL_2__2801_
timestamp 1701859473
transform -1 0 9370 0 -1 2870
box -12 -8 32 272
use FILL  FILL_2__2802_
timestamp 1701859473
transform -1 0 7230 0 -1 1830
box -12 -8 32 272
use FILL  FILL_2__2803_
timestamp 1701859473
transform 1 0 8430 0 -1 2870
box -12 -8 32 272
use FILL  FILL_2__2804_
timestamp 1701859473
transform -1 0 9490 0 -1 3390
box -12 -8 32 272
use FILL  FILL_2__2805_
timestamp 1701859473
transform -1 0 9790 0 -1 2870
box -12 -8 32 272
use FILL  FILL_2__2806_
timestamp 1701859473
transform 1 0 9550 0 -1 2870
box -12 -8 32 272
use FILL  FILL_2__2807_
timestamp 1701859473
transform 1 0 8890 0 -1 2350
box -12 -8 32 272
use FILL  FILL_2__2808_
timestamp 1701859473
transform 1 0 8650 0 -1 2350
box -12 -8 32 272
use FILL  FILL_2__2809_
timestamp 1701859473
transform 1 0 10370 0 1 2350
box -12 -8 32 272
use FILL  FILL_2__2810_
timestamp 1701859473
transform -1 0 10150 0 1 2350
box -12 -8 32 272
use FILL  FILL_2__2811_
timestamp 1701859473
transform 1 0 4930 0 -1 4430
box -12 -8 32 272
use FILL  FILL_2__2812_
timestamp 1701859473
transform -1 0 8890 0 1 4950
box -12 -8 32 272
use FILL  FILL_2__2813_
timestamp 1701859473
transform 1 0 8990 0 1 3390
box -12 -8 32 272
use FILL  FILL_2__2814_
timestamp 1701859473
transform -1 0 8810 0 -1 4430
box -12 -8 32 272
use FILL  FILL_2__2815_
timestamp 1701859473
transform -1 0 8590 0 1 3910
box -12 -8 32 272
use FILL  FILL_2__2816_
timestamp 1701859473
transform -1 0 8210 0 1 4950
box -12 -8 32 272
use FILL  FILL_2__2817_
timestamp 1701859473
transform 1 0 8650 0 1 4950
box -12 -8 32 272
use FILL  FILL_2__2818_
timestamp 1701859473
transform 1 0 8350 0 -1 4430
box -12 -8 32 272
use FILL  FILL_2__2819_
timestamp 1701859473
transform 1 0 8550 0 -1 4430
box -12 -8 32 272
use FILL  FILL_2__2820_
timestamp 1701859473
transform -1 0 9510 0 1 2350
box -12 -8 32 272
use FILL  FILL_2__2821_
timestamp 1701859473
transform 1 0 9030 0 1 2350
box -12 -8 32 272
use FILL  FILL_2__2822_
timestamp 1701859473
transform -1 0 9030 0 1 1830
box -12 -8 32 272
use FILL  FILL_2__2823_
timestamp 1701859473
transform -1 0 8810 0 1 2350
box -12 -8 32 272
use FILL  FILL_2__2824_
timestamp 1701859473
transform 1 0 9930 0 -1 3390
box -12 -8 32 272
use FILL  FILL_2__2825_
timestamp 1701859473
transform -1 0 10650 0 -1 3390
box -12 -8 32 272
use FILL  FILL_2__2826_
timestamp 1701859473
transform 1 0 9510 0 1 790
box -12 -8 32 272
use FILL  FILL_2__2827_
timestamp 1701859473
transform -1 0 9250 0 -1 1830
box -12 -8 32 272
use FILL  FILL_2__2828_
timestamp 1701859473
transform 1 0 6970 0 -1 1830
box -12 -8 32 272
use FILL  FILL_2__2829_
timestamp 1701859473
transform -1 0 9990 0 1 2870
box -12 -8 32 272
use FILL  FILL_2__2830_
timestamp 1701859473
transform 1 0 8290 0 -1 3390
box -12 -8 32 272
use FILL  FILL_2__2831_
timestamp 1701859473
transform 1 0 8330 0 1 3910
box -12 -8 32 272
use FILL  FILL_2__2832_
timestamp 1701859473
transform -1 0 9310 0 1 2350
box -12 -8 32 272
use FILL  FILL_2__2833_
timestamp 1701859473
transform -1 0 9250 0 -1 3390
box -12 -8 32 272
use FILL  FILL_2__2834_
timestamp 1701859473
transform -1 0 9010 0 -1 3390
box -12 -8 32 272
use FILL  FILL_2__2835_
timestamp 1701859473
transform -1 0 9310 0 1 790
box -12 -8 32 272
use FILL  FILL_2__2836_
timestamp 1701859473
transform 1 0 8890 0 1 1310
box -12 -8 32 272
use FILL  FILL_2__2837_
timestamp 1701859473
transform -1 0 9570 0 1 1310
box -12 -8 32 272
use FILL  FILL_2__2838_
timestamp 1701859473
transform -1 0 9690 0 1 3390
box -12 -8 32 272
use FILL  FILL_2__2839_
timestamp 1701859473
transform -1 0 9730 0 -1 3390
box -12 -8 32 272
use FILL  FILL_2__2840_
timestamp 1701859473
transform 1 0 9050 0 -1 270
box -12 -8 32 272
use FILL  FILL_2__2841_
timestamp 1701859473
transform -1 0 8850 0 -1 270
box -12 -8 32 272
use FILL  FILL_2__2842_
timestamp 1701859473
transform 1 0 9270 0 -1 270
box -12 -8 32 272
use FILL  FILL_2__2843_
timestamp 1701859473
transform 1 0 9510 0 -1 270
box -12 -8 32 272
use FILL  FILL_2__2844_
timestamp 1701859473
transform 1 0 9310 0 1 270
box -12 -8 32 272
use FILL  FILL_2__2845_
timestamp 1701859473
transform -1 0 9990 0 1 270
box -12 -8 32 272
use FILL  FILL_2__2846_
timestamp 1701859473
transform 1 0 9730 0 1 270
box -12 -8 32 272
use FILL  FILL_2__2847_
timestamp 1701859473
transform -1 0 11130 0 -1 10670
box -12 -8 32 272
use FILL  FILL_2__2848_
timestamp 1701859473
transform -1 0 10610 0 -1 1310
box -12 -8 32 272
use FILL  FILL_2__2849_
timestamp 1701859473
transform -1 0 10950 0 1 1310
box -12 -8 32 272
use FILL  FILL_2__2850_
timestamp 1701859473
transform -1 0 11090 0 -1 1830
box -12 -8 32 272
use FILL  FILL_2__2851_
timestamp 1701859473
transform 1 0 10690 0 -1 3910
box -12 -8 32 272
use FILL  FILL_2__2852_
timestamp 1701859473
transform -1 0 8890 0 1 270
box -12 -8 32 272
use FILL  FILL_2__2853_
timestamp 1701859473
transform -1 0 9110 0 1 270
box -12 -8 32 272
use FILL  FILL_2__2854_
timestamp 1701859473
transform 1 0 10610 0 1 790
box -12 -8 32 272
use FILL  FILL_2__2855_
timestamp 1701859473
transform -1 0 9810 0 1 1310
box -12 -8 32 272
use FILL  FILL_2__2856_
timestamp 1701859473
transform -1 0 10470 0 1 1310
box -12 -8 32 272
use FILL  FILL_2__2857_
timestamp 1701859473
transform -1 0 10710 0 1 1310
box -12 -8 32 272
use FILL  FILL_2__2858_
timestamp 1701859473
transform -1 0 11070 0 1 1830
box -12 -8 32 272
use FILL  FILL_2__2859_
timestamp 1701859473
transform 1 0 10930 0 -1 3910
box -12 -8 32 272
use FILL  FILL_2__2860_
timestamp 1701859473
transform 1 0 10850 0 -1 3390
box -12 -8 32 272
use FILL  FILL_2__2861_
timestamp 1701859473
transform 1 0 9730 0 -1 270
box -12 -8 32 272
use FILL  FILL_2__2862_
timestamp 1701859473
transform 1 0 8590 0 -1 270
box -12 -8 32 272
use FILL  FILL_2__2863_
timestamp 1701859473
transform -1 0 10230 0 1 270
box -12 -8 32 272
use FILL  FILL_2__2864_
timestamp 1701859473
transform 1 0 10470 0 1 270
box -12 -8 32 272
use FILL  FILL_2__2865_
timestamp 1701859473
transform -1 0 10710 0 1 270
box -12 -8 32 272
use FILL  FILL_2__2866_
timestamp 1701859473
transform -1 0 11090 0 -1 790
box -12 -8 32 272
use FILL  FILL_2__2867_
timestamp 1701859473
transform 1 0 11050 0 -1 3390
box -12 -8 32 272
use FILL  FILL_2__2868_
timestamp 1701859473
transform 1 0 11030 0 1 790
box -12 -8 32 272
use FILL  FILL_2__2869_
timestamp 1701859473
transform 1 0 10150 0 1 790
box -12 -8 32 272
use FILL  FILL_2__2870_
timestamp 1701859473
transform -1 0 10370 0 1 790
box -12 -8 32 272
use FILL  FILL_2__2871_
timestamp 1701859473
transform -1 0 10810 0 1 790
box -12 -8 32 272
use FILL  FILL_2__2872_
timestamp 1701859473
transform -1 0 11150 0 1 1310
box -12 -8 32 272
use FILL  FILL_2__2873_
timestamp 1701859473
transform -1 0 9930 0 1 3390
box -12 -8 32 272
use FILL  FILL_2__2874_
timestamp 1701859473
transform -1 0 10170 0 1 3390
box -12 -8 32 272
use FILL  FILL_2__2875_
timestamp 1701859473
transform -1 0 10750 0 -1 4950
box -12 -8 32 272
use FILL  FILL_2__2876_
timestamp 1701859473
transform -1 0 9710 0 1 1830
box -12 -8 32 272
use FILL  FILL_2__2877_
timestamp 1701859473
transform 1 0 9890 0 1 1830
box -12 -8 32 272
use FILL  FILL_2__2878_
timestamp 1701859473
transform 1 0 9710 0 -1 1310
box -12 -8 32 272
use FILL  FILL_2__2879_
timestamp 1701859473
transform -1 0 9950 0 -1 1310
box -12 -8 32 272
use FILL  FILL_2__2880_
timestamp 1701859473
transform 1 0 9450 0 1 1830
box -12 -8 32 272
use FILL  FILL_2__2881_
timestamp 1701859473
transform 1 0 10830 0 -1 790
box -12 -8 32 272
use FILL  FILL_2__2882_
timestamp 1701859473
transform -1 0 9510 0 -1 1310
box -12 -8 32 272
use FILL  FILL_2__2883_
timestamp 1701859473
transform -1 0 10410 0 -1 1310
box -12 -8 32 272
use FILL  FILL_2__2884_
timestamp 1701859473
transform 1 0 11050 0 -1 1310
box -12 -8 32 272
use FILL  FILL_2__2885_
timestamp 1701859473
transform -1 0 10830 0 -1 1310
box -12 -8 32 272
use FILL  FILL_2__2886_
timestamp 1701859473
transform 1 0 10590 0 1 1830
box -12 -8 32 272
use FILL  FILL_2__2887_
timestamp 1701859473
transform 1 0 10150 0 -1 4430
box -12 -8 32 272
use FILL  FILL_2__2888_
timestamp 1701859473
transform -1 0 3970 0 1 5470
box -12 -8 32 272
use FILL  FILL_2__2889_
timestamp 1701859473
transform 1 0 6090 0 1 2350
box -12 -8 32 272
use FILL  FILL_2__2890_
timestamp 1701859473
transform -1 0 8370 0 1 5990
box -12 -8 32 272
use FILL  FILL_2__2891_
timestamp 1701859473
transform -1 0 8170 0 1 5990
box -12 -8 32 272
use FILL  FILL_2__2892_
timestamp 1701859473
transform 1 0 7390 0 -1 5470
box -12 -8 32 272
use FILL  FILL_2__2893_
timestamp 1701859473
transform 1 0 7210 0 1 5470
box -12 -8 32 272
use FILL  FILL_2__2894_
timestamp 1701859473
transform 1 0 6490 0 -1 6510
box -12 -8 32 272
use FILL  FILL_2__2895_
timestamp 1701859473
transform 1 0 6630 0 1 6510
box -12 -8 32 272
use FILL  FILL_2__2896_
timestamp 1701859473
transform -1 0 7890 0 -1 5470
box -12 -8 32 272
use FILL  FILL_2__2897_
timestamp 1701859473
transform 1 0 7690 0 1 5470
box -12 -8 32 272
use FILL  FILL_2__2898_
timestamp 1701859473
transform 1 0 7210 0 -1 6510
box -12 -8 32 272
use FILL  FILL_2__2899_
timestamp 1701859473
transform 1 0 6730 0 -1 6510
box -12 -8 32 272
use FILL  FILL_2__2900_
timestamp 1701859473
transform -1 0 6270 0 -1 6510
box -12 -8 32 272
use FILL  FILL_2__2901_
timestamp 1701859473
transform 1 0 6010 0 -1 6510
box -12 -8 32 272
use FILL  FILL_2__2902_
timestamp 1701859473
transform -1 0 7930 0 1 5990
box -12 -8 32 272
use FILL  FILL_2__2903_
timestamp 1701859473
transform 1 0 7210 0 1 5990
box -12 -8 32 272
use FILL  FILL_2__2904_
timestamp 1701859473
transform 1 0 8330 0 -1 5470
box -12 -8 32 272
use FILL  FILL_2__2905_
timestamp 1701859473
transform 1 0 8350 0 1 5470
box -12 -8 32 272
use FILL  FILL_2__2906_
timestamp 1701859473
transform 1 0 8090 0 -1 5990
box -12 -8 32 272
use FILL  FILL_2__2907_
timestamp 1701859473
transform -1 0 7870 0 -1 5990
box -12 -8 32 272
use FILL  FILL_2__2908_
timestamp 1701859473
transform -1 0 8190 0 -1 4950
box -12 -8 32 272
use FILL  FILL_2__2909_
timestamp 1701859473
transform 1 0 3330 0 -1 4430
box -12 -8 32 272
use FILL  FILL_2__2910_
timestamp 1701859473
transform -1 0 6490 0 -1 4430
box -12 -8 32 272
use FILL  FILL_2__2911_
timestamp 1701859473
transform -1 0 6830 0 1 4430
box -12 -8 32 272
use FILL  FILL_2__2912_
timestamp 1701859473
transform 1 0 8610 0 -1 4950
box -12 -8 32 272
use FILL  FILL_2__2913_
timestamp 1701859473
transform -1 0 6790 0 -1 4950
box -12 -8 32 272
use FILL  FILL_2__2914_
timestamp 1701859473
transform 1 0 7050 0 -1 8070
box -12 -8 32 272
use FILL  FILL_2__2915_
timestamp 1701859473
transform 1 0 7170 0 -1 5990
box -12 -8 32 272
use FILL  FILL_2__2916_
timestamp 1701859473
transform 1 0 6930 0 -1 5990
box -12 -8 32 272
use FILL  FILL_2__2917_
timestamp 1701859473
transform -1 0 6310 0 -1 5990
box -12 -8 32 272
use FILL  FILL_2__2918_
timestamp 1701859473
transform 1 0 6230 0 1 5470
box -12 -8 32 272
use FILL  FILL_2__2919_
timestamp 1701859473
transform 1 0 6150 0 1 4950
box -12 -8 32 272
use FILL  FILL_2__2920_
timestamp 1701859473
transform 1 0 5910 0 1 4950
box -12 -8 32 272
use FILL  FILL_2__2921_
timestamp 1701859473
transform -1 0 7370 0 -1 3910
box -12 -8 32 272
use FILL  FILL_2__2922_
timestamp 1701859473
transform -1 0 7410 0 1 3910
box -12 -8 32 272
use FILL  FILL_2__2923_
timestamp 1701859473
transform -1 0 6730 0 -1 4430
box -12 -8 32 272
use FILL  FILL_2__2924_
timestamp 1701859473
transform 1 0 6350 0 1 4950
box -12 -8 32 272
use FILL  FILL_2__2925_
timestamp 1701859473
transform 1 0 7250 0 1 7550
box -12 -8 32 272
use FILL  FILL_2__2926_
timestamp 1701859473
transform -1 0 7490 0 1 4430
box -12 -8 32 272
use FILL  FILL_2__2927_
timestamp 1701859473
transform 1 0 7270 0 -1 4950
box -12 -8 32 272
use FILL  FILL_2__2928_
timestamp 1701859473
transform 1 0 7010 0 -1 4950
box -12 -8 32 272
use FILL  FILL_2__2929_
timestamp 1701859473
transform -1 0 6590 0 1 4950
box -12 -8 32 272
use FILL  FILL_2__2930_
timestamp 1701859473
transform 1 0 6130 0 1 1830
box -12 -8 32 272
use FILL  FILL_2__2931_
timestamp 1701859473
transform 1 0 7010 0 -1 2870
box -12 -8 32 272
use FILL  FILL_2__2932_
timestamp 1701859473
transform 1 0 5170 0 -1 4430
box -12 -8 32 272
use FILL  FILL_2__2933_
timestamp 1701859473
transform 1 0 5370 0 -1 4430
box -12 -8 32 272
use FILL  FILL_2__2934_
timestamp 1701859473
transform 1 0 5610 0 -1 4430
box -12 -8 32 272
use FILL  FILL_2__2935_
timestamp 1701859473
transform 1 0 6430 0 1 6510
box -12 -8 32 272
use FILL  FILL_2__2936_
timestamp 1701859473
transform 1 0 6310 0 -1 4950
box -12 -8 32 272
use FILL  FILL_2__2937_
timestamp 1701859473
transform 1 0 6530 0 -1 4950
box -12 -8 32 272
use FILL  FILL_2__2938_
timestamp 1701859473
transform 1 0 5010 0 1 4950
box -12 -8 32 272
use FILL  FILL_2__2939_
timestamp 1701859473
transform 1 0 4790 0 1 4950
box -12 -8 32 272
use FILL  FILL_2__2940_
timestamp 1701859473
transform -1 0 5850 0 -1 5470
box -12 -8 32 272
use FILL  FILL_2__2941_
timestamp 1701859473
transform 1 0 5610 0 -1 5470
box -12 -8 32 272
use FILL  FILL_2__2942_
timestamp 1701859473
transform -1 0 9310 0 1 4430
box -12 -8 32 272
use FILL  FILL_2__2943_
timestamp 1701859473
transform 1 0 6270 0 -1 4430
box -12 -8 32 272
use FILL  FILL_2__2944_
timestamp 1701859473
transform -1 0 6290 0 1 3910
box -12 -8 32 272
use FILL  FILL_2__2945_
timestamp 1701859473
transform -1 0 6370 0 1 4430
box -12 -8 32 272
use FILL  FILL_2__2946_
timestamp 1701859473
transform 1 0 6130 0 1 4430
box -12 -8 32 272
use FILL  FILL_2__2947_
timestamp 1701859473
transform -1 0 6530 0 -1 5990
box -12 -8 32 272
use FILL  FILL_2__2948_
timestamp 1701859473
transform 1 0 6070 0 -1 5990
box -12 -8 32 272
use FILL  FILL_2__2949_
timestamp 1701859473
transform -1 0 5890 0 -1 5990
box -12 -8 32 272
use FILL  FILL_2__2950_
timestamp 1701859473
transform 1 0 5750 0 1 5470
box -12 -8 32 272
use FILL  FILL_2__2951_
timestamp 1701859473
transform -1 0 6010 0 1 5470
box -12 -8 32 272
use FILL  FILL_2__2952_
timestamp 1701859473
transform -1 0 6090 0 -1 4950
box -12 -8 32 272
use FILL  FILL_2__2953_
timestamp 1701859473
transform -1 0 4370 0 1 4950
box -12 -8 32 272
use FILL  FILL_2__2954_
timestamp 1701859473
transform -1 0 6630 0 1 4430
box -12 -8 32 272
use FILL  FILL_2__2955_
timestamp 1701859473
transform -1 0 5910 0 1 4430
box -12 -8 32 272
use FILL  FILL_2__2956_
timestamp 1701859473
transform 1 0 5190 0 1 4430
box -12 -8 32 272
use FILL  FILL_2__2957_
timestamp 1701859473
transform 1 0 5130 0 -1 4950
box -12 -8 32 272
use FILL  FILL_2__2958_
timestamp 1701859473
transform -1 0 5450 0 1 4430
box -12 -8 32 272
use FILL  FILL_2__2959_
timestamp 1701859473
transform 1 0 6950 0 -1 5470
box -12 -8 32 272
use FILL  FILL_2__2960_
timestamp 1701859473
transform -1 0 6490 0 1 5470
box -12 -8 32 272
use FILL  FILL_2__2961_
timestamp 1701859473
transform 1 0 6250 0 -1 5470
box -12 -8 32 272
use FILL  FILL_2__2962_
timestamp 1701859473
transform -1 0 6510 0 -1 5470
box -12 -8 32 272
use FILL  FILL_2__2963_
timestamp 1701859473
transform -1 0 6750 0 -1 5470
box -12 -8 32 272
use FILL  FILL_2__2964_
timestamp 1701859473
transform -1 0 5390 0 -1 4950
box -12 -8 32 272
use FILL  FILL_2__2965_
timestamp 1701859473
transform 1 0 4890 0 -1 4950
box -12 -8 32 272
use FILL  FILL_2__2966_
timestamp 1701859473
transform -1 0 6350 0 1 2350
box -12 -8 32 272
use FILL  FILL_2__2967_
timestamp 1701859473
transform 1 0 7610 0 1 3910
box -12 -8 32 272
use FILL  FILL_2__2968_
timestamp 1701859473
transform -1 0 6930 0 -1 3910
box -12 -8 32 272
use FILL  FILL_2__2969_
timestamp 1701859473
transform -1 0 7150 0 -1 3910
box -12 -8 32 272
use FILL  FILL_2__2970_
timestamp 1701859473
transform -1 0 7190 0 1 3910
box -12 -8 32 272
use FILL  FILL_2__2971_
timestamp 1701859473
transform -1 0 6710 0 1 3910
box -12 -8 32 272
use FILL  FILL_2__2972_
timestamp 1701859473
transform 1 0 6930 0 1 3910
box -12 -8 32 272
use FILL  FILL_2__2973_
timestamp 1701859473
transform -1 0 7050 0 1 4430
box -12 -8 32 272
use FILL  FILL_2__2974_
timestamp 1701859473
transform 1 0 6950 0 -1 4430
box -12 -8 32 272
use FILL  FILL_2__2975_
timestamp 1701859473
transform -1 0 7710 0 -1 4430
box -12 -8 32 272
use FILL  FILL_2__2976_
timestamp 1701859473
transform -1 0 7470 0 -1 4430
box -12 -8 32 272
use FILL  FILL_2__2977_
timestamp 1701859473
transform 1 0 7190 0 -1 4430
box -12 -8 32 272
use FILL  FILL_2__2978_
timestamp 1701859473
transform 1 0 7250 0 1 4430
box -12 -8 32 272
use FILL  FILL_2__2979_
timestamp 1701859473
transform -1 0 3590 0 -1 4950
box -12 -8 32 272
use FILL  FILL_2__2980_
timestamp 1701859473
transform -1 0 2970 0 1 7550
box -12 -8 32 272
use FILL  FILL_2__2981_
timestamp 1701859473
transform 1 0 3490 0 1 4950
box -12 -8 32 272
use FILL  FILL_2__2982_
timestamp 1701859473
transform 1 0 9550 0 1 6510
box -12 -8 32 272
use FILL  FILL_2__2983_
timestamp 1701859473
transform 1 0 1870 0 1 4430
box -12 -8 32 272
use FILL  FILL_2__2984_
timestamp 1701859473
transform -1 0 3490 0 -1 3910
box -12 -8 32 272
use FILL  FILL_2__2985_
timestamp 1701859473
transform 1 0 3650 0 1 4430
box -12 -8 32 272
use FILL  FILL_2__2986_
timestamp 1701859473
transform -1 0 5850 0 -1 4430
box -12 -8 32 272
use FILL  FILL_2__2987_
timestamp 1701859473
transform -1 0 5670 0 1 4430
box -12 -8 32 272
use FILL  FILL_2__2988_
timestamp 1701859473
transform 1 0 9330 0 1 6510
box -12 -8 32 272
use FILL  FILL_2__2989_
timestamp 1701859473
transform 1 0 5950 0 1 6510
box -12 -8 32 272
use FILL  FILL_2__2990_
timestamp 1701859473
transform -1 0 6210 0 1 6510
box -12 -8 32 272
use FILL  FILL_2__2991_
timestamp 1701859473
transform 1 0 7110 0 1 6510
box -12 -8 32 272
use FILL  FILL_2__2992_
timestamp 1701859473
transform 1 0 9630 0 1 7030
box -12 -8 32 272
use FILL  FILL_2__2993_
timestamp 1701859473
transform 1 0 9830 0 1 7030
box -12 -8 32 272
use FILL  FILL_2__2994_
timestamp 1701859473
transform -1 0 10750 0 -1 7550
box -12 -8 32 272
use FILL  FILL_2__2995_
timestamp 1701859473
transform -1 0 7550 0 -1 7550
box -12 -8 32 272
use FILL  FILL_2__2996_
timestamp 1701859473
transform 1 0 7450 0 1 7550
box -12 -8 32 272
use FILL  FILL_2__2997_
timestamp 1701859473
transform -1 0 7330 0 -1 7550
box -12 -8 32 272
use FILL  FILL_2__2998_
timestamp 1701859473
transform -1 0 6390 0 -1 7550
box -12 -8 32 272
use FILL  FILL_2__2999_
timestamp 1701859473
transform 1 0 6110 0 1 7550
box -12 -8 32 272
use FILL  FILL_2__3000_
timestamp 1701859473
transform -1 0 5950 0 -1 7550
box -12 -8 32 272
use FILL  FILL_2__3001_
timestamp 1701859473
transform -1 0 5730 0 -1 7550
box -12 -8 32 272
use FILL  FILL_2__3002_
timestamp 1701859473
transform -1 0 6150 0 -1 7550
box -12 -8 32 272
use FILL  FILL_2__3003_
timestamp 1701859473
transform -1 0 6330 0 1 7550
box -12 -8 32 272
use FILL  FILL_2__3004_
timestamp 1701859473
transform 1 0 8130 0 1 7550
box -12 -8 32 272
use FILL  FILL_2__3005_
timestamp 1701859473
transform 1 0 10950 0 -1 7550
box -12 -8 32 272
use FILL  FILL_2__3006_
timestamp 1701859473
transform -1 0 10430 0 1 7550
box -12 -8 32 272
use FILL  FILL_2__3007_
timestamp 1701859473
transform 1 0 6950 0 1 7030
box -12 -8 32 272
use FILL  FILL_2__3008_
timestamp 1701859473
transform -1 0 6510 0 1 7030
box -12 -8 32 272
use FILL  FILL_2__3009_
timestamp 1701859473
transform -1 0 5910 0 -1 7030
box -12 -8 32 272
use FILL  FILL_2__3010_
timestamp 1701859473
transform 1 0 6130 0 -1 7030
box -12 -8 32 272
use FILL  FILL_2__3011_
timestamp 1701859473
transform 1 0 6710 0 1 7030
box -12 -8 32 272
use FILL  FILL_2__3012_
timestamp 1701859473
transform -1 0 7830 0 -1 7030
box -12 -8 32 272
use FILL  FILL_2__3013_
timestamp 1701859473
transform 1 0 8270 0 -1 7030
box -12 -8 32 272
use FILL  FILL_2__3014_
timestamp 1701859473
transform 1 0 10630 0 1 7550
box -12 -8 32 272
use FILL  FILL_2__3015_
timestamp 1701859473
transform -1 0 6350 0 -1 7030
box -12 -8 32 272
use FILL  FILL_2__3016_
timestamp 1701859473
transform -1 0 7230 0 1 7030
box -12 -8 32 272
use FILL  FILL_2__3017_
timestamp 1701859473
transform 1 0 6570 0 -1 7030
box -12 -8 32 272
use FILL  FILL_2__3018_
timestamp 1701859473
transform -1 0 6870 0 -1 7030
box -12 -8 32 272
use FILL  FILL_2__3019_
timestamp 1701859473
transform -1 0 7110 0 -1 7030
box -12 -8 32 272
use FILL  FILL_2__3020_
timestamp 1701859473
transform 1 0 8270 0 1 7030
box -12 -8 32 272
use FILL  FILL_2__3021_
timestamp 1701859473
transform -1 0 9330 0 -1 8070
box -12 -8 32 272
use FILL  FILL_2__3022_
timestamp 1701859473
transform 1 0 9510 0 -1 8070
box -12 -8 32 272
use FILL  FILL_2__3023_
timestamp 1701859473
transform -1 0 5730 0 1 6510
box -12 -8 32 272
use FILL  FILL_2__3024_
timestamp 1701859473
transform 1 0 5470 0 1 6510
box -12 -8 32 272
use FILL  FILL_2__3025_
timestamp 1701859473
transform -1 0 5490 0 -1 6510
box -12 -8 32 272
use FILL  FILL_2__3026_
timestamp 1701859473
transform 1 0 10910 0 -1 5990
box -12 -8 32 272
use FILL  FILL_2__3027_
timestamp 1701859473
transform -1 0 11150 0 -1 5990
box -12 -8 32 272
use FILL  FILL_2__3028_
timestamp 1701859473
transform -1 0 9770 0 -1 8070
box -12 -8 32 272
use FILL  FILL_2__3029_
timestamp 1701859473
transform -1 0 7090 0 -1 7550
box -12 -8 32 272
use FILL  FILL_2__3030_
timestamp 1701859473
transform -1 0 8070 0 -1 7030
box -12 -8 32 272
use FILL  FILL_2__3031_
timestamp 1701859473
transform 1 0 8050 0 1 7030
box -12 -8 32 272
use FILL  FILL_2__3032_
timestamp 1701859473
transform 1 0 7670 0 1 7550
box -12 -8 32 272
use FILL  FILL_2__3033_
timestamp 1701859473
transform -1 0 6750 0 1 8070
box -12 -8 32 272
use FILL  FILL_2__3034_
timestamp 1701859473
transform -1 0 7730 0 -1 8070
box -12 -8 32 272
use FILL  FILL_2__3035_
timestamp 1701859473
transform 1 0 7470 0 -1 8070
box -12 -8 32 272
use FILL  FILL_2__3036_
timestamp 1701859473
transform -1 0 6950 0 1 8070
box -12 -8 32 272
use FILL  FILL_2__3037_
timestamp 1701859473
transform -1 0 6510 0 1 8070
box -12 -8 32 272
use FILL  FILL_2__3038_
timestamp 1701859473
transform -1 0 7130 0 1 8070
box -12 -8 32 272
use FILL  FILL_2__3039_
timestamp 1701859473
transform 1 0 7350 0 1 8070
box -12 -8 32 272
use FILL  FILL_2__3040_
timestamp 1701859473
transform 1 0 9690 0 1 7550
box -12 -8 32 272
use FILL  FILL_2__3041_
timestamp 1701859473
transform -1 0 9550 0 -1 6510
box -12 -8 32 272
use FILL  FILL_2__3042_
timestamp 1701859473
transform 1 0 7250 0 -1 8070
box -12 -8 32 272
use FILL  FILL_2__3043_
timestamp 1701859473
transform -1 0 6570 0 1 7550
box -12 -8 32 272
use FILL  FILL_2__3044_
timestamp 1701859473
transform -1 0 6610 0 -1 7550
box -12 -8 32 272
use FILL  FILL_2__3045_
timestamp 1701859473
transform 1 0 6830 0 -1 7550
box -12 -8 32 272
use FILL  FILL_2__3046_
timestamp 1701859473
transform -1 0 7790 0 1 6510
box -12 -8 32 272
use FILL  FILL_2__3047_
timestamp 1701859473
transform 1 0 9130 0 1 6510
box -12 -8 32 272
use FILL  FILL_2__3048_
timestamp 1701859473
transform 1 0 9750 0 -1 6510
box -12 -8 32 272
use FILL  FILL_2__3049_
timestamp 1701859473
transform -1 0 6830 0 1 7550
box -12 -8 32 272
use FILL  FILL_2__3050_
timestamp 1701859473
transform -1 0 7050 0 1 7550
box -12 -8 32 272
use FILL  FILL_2__3051_
timestamp 1701859473
transform -1 0 7790 0 1 7030
box -12 -8 32 272
use FILL  FILL_2__3052_
timestamp 1701859473
transform 1 0 7490 0 1 7030
box -12 -8 32 272
use FILL  FILL_2__3053_
timestamp 1701859473
transform 1 0 7330 0 -1 7030
box -12 -8 32 272
use FILL  FILL_2__3054_
timestamp 1701859473
transform -1 0 7590 0 -1 7030
box -12 -8 32 272
use FILL  FILL_2__3055_
timestamp 1701859473
transform 1 0 8010 0 1 6510
box -12 -8 32 272
use FILL  FILL_2__3056_
timestamp 1701859473
transform -1 0 9530 0 1 5470
box -12 -8 32 272
use FILL  FILL_2__3057_
timestamp 1701859473
transform -1 0 9290 0 1 5470
box -12 -8 32 272
use FILL  FILL_2__3058_
timestamp 1701859473
transform 1 0 8710 0 -1 7550
box -12 -8 32 272
use FILL  FILL_2__3059_
timestamp 1701859473
transform -1 0 8590 0 -1 5990
box -12 -8 32 272
use FILL  FILL_2__3060_
timestamp 1701859473
transform 1 0 9770 0 1 6510
box -12 -8 32 272
use FILL  FILL_2__3061_
timestamp 1701859473
transform 1 0 10010 0 1 6510
box -12 -8 32 272
use FILL  FILL_2__3062_
timestamp 1701859473
transform -1 0 9630 0 -1 7550
box -12 -8 32 272
use FILL  FILL_2__3063_
timestamp 1701859473
transform 1 0 9370 0 -1 7550
box -12 -8 32 272
use FILL  FILL_2__3064_
timestamp 1701859473
transform -1 0 10330 0 -1 7030
box -12 -8 32 272
use FILL  FILL_2__3065_
timestamp 1701859473
transform -1 0 10570 0 -1 7030
box -12 -8 32 272
use FILL  FILL_2__3066_
timestamp 1701859473
transform -1 0 8490 0 -1 7550
box -12 -8 32 272
use FILL  FILL_2__3067_
timestamp 1701859473
transform 1 0 8230 0 -1 7550
box -12 -8 32 272
use FILL  FILL_2__3068_
timestamp 1701859473
transform 1 0 10190 0 -1 5990
box -12 -8 32 272
use FILL  FILL_2__3069_
timestamp 1701859473
transform 1 0 10430 0 -1 5990
box -12 -8 32 272
use FILL  FILL_2__3070_
timestamp 1701859473
transform 1 0 8890 0 -1 7550
box -12 -8 32 272
use FILL  FILL_2__3071_
timestamp 1701859473
transform -1 0 9150 0 -1 7550
box -12 -8 32 272
use FILL  FILL_2__3072_
timestamp 1701859473
transform -1 0 9770 0 1 5990
box -12 -8 32 272
use FILL  FILL_2__3073_
timestamp 1701859473
transform -1 0 9990 0 1 5990
box -12 -8 32 272
use FILL  FILL_2__3074_
timestamp 1701859473
transform 1 0 8810 0 1 5990
box -12 -8 32 272
use FILL  FILL_2__3075_
timestamp 1701859473
transform 1 0 8810 0 -1 5990
box -12 -8 32 272
use FILL  FILL_2__3076_
timestamp 1701859473
transform 1 0 10710 0 1 6510
box -12 -8 32 272
use FILL  FILL_2__3077_
timestamp 1701859473
transform 1 0 10910 0 1 6510
box -12 -8 32 272
use FILL  FILL_2__3078_
timestamp 1701859473
transform -1 0 8710 0 -1 7030
box -12 -8 32 272
use FILL  FILL_2__3079_
timestamp 1701859473
transform -1 0 8490 0 -1 7030
box -12 -8 32 272
use FILL  FILL_2__3080_
timestamp 1701859473
transform 1 0 10970 0 -1 8590
box -12 -8 32 272
use FILL  FILL_2__3081_
timestamp 1701859473
transform -1 0 10970 0 -1 270
box -12 -8 32 272
use FILL  FILL_2__3082_
timestamp 1701859473
transform 1 0 10070 0 -1 8590
box -12 -8 32 272
use FILL  FILL_2__3083_
timestamp 1701859473
transform -1 0 9850 0 -1 8590
box -12 -8 32 272
use FILL  FILL_2__3084_
timestamp 1701859473
transform -1 0 9030 0 1 7550
box -12 -8 32 272
use FILL  FILL_2__3085_
timestamp 1701859473
transform 1 0 8930 0 1 7030
box -12 -8 32 272
use FILL  FILL_2__3086_
timestamp 1701859473
transform -1 0 10690 0 1 5990
box -12 -8 32 272
use FILL  FILL_2__3087_
timestamp 1701859473
transform 1 0 10890 0 1 5990
box -12 -8 32 272
use FILL  FILL_2__3088_
timestamp 1701859473
transform 1 0 8250 0 1 8070
box -12 -8 32 272
use FILL  FILL_2__3089_
timestamp 1701859473
transform -1 0 8030 0 1 8070
box -12 -8 32 272
use FILL  FILL_2__3090_
timestamp 1701859473
transform -1 0 11130 0 1 4950
box -12 -8 32 272
use FILL  FILL_2__3091_
timestamp 1701859473
transform 1 0 10870 0 1 4950
box -12 -8 32 272
use FILL  FILL_2__3092_
timestamp 1701859473
transform 1 0 8790 0 -1 5470
box -12 -8 32 272
use FILL  FILL_2__3093_
timestamp 1701859473
transform -1 0 9030 0 -1 5470
box -12 -8 32 272
use FILL  FILL_2__3094_
timestamp 1701859473
transform -1 0 10230 0 -1 5470
box -12 -8 32 272
use FILL  FILL_2__3095_
timestamp 1701859473
transform 1 0 10170 0 1 5470
box -12 -8 32 272
use FILL  FILL_2__3096_
timestamp 1701859473
transform 1 0 8910 0 1 6510
box -12 -8 32 272
use FILL  FILL_2__3097_
timestamp 1701859473
transform -1 0 8690 0 1 6510
box -12 -8 32 272
use FILL  FILL_2__3098_
timestamp 1701859473
transform -1 0 10390 0 1 8070
box -12 -8 32 272
use FILL  FILL_2__3099_
timestamp 1701859473
transform -1 0 11150 0 -1 8070
box -12 -8 32 272
use FILL  FILL_2__3100_
timestamp 1701859473
transform 1 0 10150 0 1 8070
box -12 -8 32 272
use FILL  FILL_2__3101_
timestamp 1701859473
transform 1 0 10290 0 -1 8590
box -12 -8 32 272
use FILL  FILL_2__3102_
timestamp 1701859473
transform 1 0 8370 0 -1 8070
box -12 -8 32 272
use FILL  FILL_2__3103_
timestamp 1701859473
transform -1 0 8350 0 1 7550
box -12 -8 32 272
use FILL  FILL_2__3104_
timestamp 1701859473
transform -1 0 11150 0 1 6510
box -12 -8 32 272
use FILL  FILL_2__3105_
timestamp 1701859473
transform -1 0 10950 0 -1 4950
box -12 -8 32 272
use FILL  FILL_2__3106_
timestamp 1701859473
transform 1 0 9370 0 -1 8590
box -12 -8 32 272
use FILL  FILL_2__3107_
timestamp 1701859473
transform -1 0 9610 0 -1 8590
box -12 -8 32 272
use FILL  FILL_2__3108_
timestamp 1701859473
transform 1 0 9970 0 1 5470
box -12 -8 32 272
use FILL  FILL_2__3109_
timestamp 1701859473
transform -1 0 9750 0 1 5470
box -12 -8 32 272
use FILL  FILL_2__3110_
timestamp 1701859473
transform 1 0 8390 0 -1 6510
box -12 -8 32 272
use FILL  FILL_2__3111_
timestamp 1701859473
transform -1 0 8170 0 -1 6510
box -12 -8 32 272
use FILL  FILL_2__3112_
timestamp 1701859473
transform 1 0 510 0 -1 2870
box -12 -8 32 272
use FILL  FILL_2__3113_
timestamp 1701859473
transform 1 0 50 0 -1 2870
box -12 -8 32 272
use FILL  FILL_2__3114_
timestamp 1701859473
transform -1 0 310 0 -1 2870
box -12 -8 32 272
use FILL  FILL_2__3115_
timestamp 1701859473
transform -1 0 1190 0 1 2350
box -12 -8 32 272
use FILL  FILL_2__3116_
timestamp 1701859473
transform 1 0 950 0 -1 2350
box -12 -8 32 272
use FILL  FILL_2__3117_
timestamp 1701859473
transform 1 0 2030 0 -1 1310
box -12 -8 32 272
use FILL  FILL_2__3118_
timestamp 1701859473
transform -1 0 1410 0 -1 2350
box -12 -8 32 272
use FILL  FILL_2__3119_
timestamp 1701859473
transform -1 0 1170 0 -1 2350
box -12 -8 32 272
use FILL  FILL_2__3120_
timestamp 1701859473
transform -1 0 470 0 1 2350
box -12 -8 32 272
use FILL  FILL_2__3121_
timestamp 1701859473
transform 1 0 250 0 1 2870
box -12 -8 32 272
use FILL  FILL_2__3122_
timestamp 1701859473
transform 1 0 2510 0 -1 3390
box -12 -8 32 272
use FILL  FILL_2__3123_
timestamp 1701859473
transform 1 0 530 0 1 3390
box -12 -8 32 272
use FILL  FILL_2__3124_
timestamp 1701859473
transform -1 0 310 0 1 3390
box -12 -8 32 272
use FILL  FILL_2__3125_
timestamp 1701859473
transform -1 0 730 0 -1 2350
box -12 -8 32 272
use FILL  FILL_2__3126_
timestamp 1701859473
transform -1 0 1430 0 1 2350
box -12 -8 32 272
use FILL  FILL_2__3127_
timestamp 1701859473
transform -1 0 950 0 1 2350
box -12 -8 32 272
use FILL  FILL_2__3128_
timestamp 1701859473
transform -1 0 1890 0 1 2350
box -12 -8 32 272
use FILL  FILL_2__3129_
timestamp 1701859473
transform -1 0 1650 0 -1 2350
box -12 -8 32 272
use FILL  FILL_2__3130_
timestamp 1701859473
transform -1 0 1670 0 1 2350
box -12 -8 32 272
use FILL  FILL_2__3131_
timestamp 1701859473
transform -1 0 710 0 1 2350
box -12 -8 32 272
use FILL  FILL_2__3132_
timestamp 1701859473
transform 1 0 470 0 1 2870
box -12 -8 32 272
use FILL  FILL_2__3133_
timestamp 1701859473
transform 1 0 530 0 -1 3910
box -12 -8 32 272
use FILL  FILL_2__3134_
timestamp 1701859473
transform -1 0 1210 0 1 3390
box -12 -8 32 272
use FILL  FILL_2__3135_
timestamp 1701859473
transform 1 0 970 0 1 3390
box -12 -8 32 272
use FILL  FILL_2__3136_
timestamp 1701859473
transform -1 0 550 0 -1 3390
box -12 -8 32 272
use FILL  FILL_2__3137_
timestamp 1701859473
transform 1 0 270 0 -1 3390
box -12 -8 32 272
use FILL  FILL_2__3138_
timestamp 1701859473
transform -1 0 1670 0 1 4430
box -12 -8 32 272
use FILL  FILL_2__3139_
timestamp 1701859473
transform -1 0 1870 0 -1 3390
box -12 -8 32 272
use FILL  FILL_2__3140_
timestamp 1701859473
transform -1 0 290 0 1 3910
box -12 -8 32 272
use FILL  FILL_2__3141_
timestamp 1701859473
transform 1 0 730 0 1 4430
box -12 -8 32 272
use FILL  FILL_2__3142_
timestamp 1701859473
transform 1 0 970 0 1 4430
box -12 -8 32 272
use FILL  FILL_2__3143_
timestamp 1701859473
transform 1 0 990 0 -1 4430
box -12 -8 32 272
use FILL  FILL_2__3144_
timestamp 1701859473
transform -1 0 1230 0 -1 4430
box -12 -8 32 272
use FILL  FILL_2__3145_
timestamp 1701859473
transform -1 0 510 0 1 3910
box -12 -8 32 272
use FILL  FILL_2__3146_
timestamp 1701859473
transform -1 0 730 0 1 3910
box -12 -8 32 272
use FILL  FILL_2__3147_
timestamp 1701859473
transform 1 0 510 0 -1 4430
box -12 -8 32 272
use FILL  FILL_2__3148_
timestamp 1701859473
transform -1 0 770 0 -1 4430
box -12 -8 32 272
use FILL  FILL_2__3149_
timestamp 1701859473
transform -1 0 70 0 -1 3910
box -12 -8 32 272
use FILL  FILL_2__3150_
timestamp 1701859473
transform -1 0 930 0 1 3910
box -12 -8 32 272
use FILL  FILL_2__3151_
timestamp 1701859473
transform 1 0 50 0 1 3910
box -12 -8 32 272
use FILL  FILL_2__3152_
timestamp 1701859473
transform 1 0 50 0 -1 4430
box -12 -8 32 272
use FILL  FILL_2__3153_
timestamp 1701859473
transform -1 0 290 0 -1 4430
box -12 -8 32 272
use FILL  FILL_2__3154_
timestamp 1701859473
transform -1 0 790 0 -1 3390
box -12 -8 32 272
use FILL  FILL_2__3155_
timestamp 1701859473
transform -1 0 70 0 1 2870
box -12 -8 32 272
use FILL  FILL_2__3156_
timestamp 1701859473
transform 1 0 50 0 -1 3390
box -12 -8 32 272
use FILL  FILL_2__3157_
timestamp 1701859473
transform -1 0 70 0 1 3390
box -12 -8 32 272
use FILL  FILL_2__3158_
timestamp 1701859473
transform 1 0 50 0 1 4430
box -12 -8 32 272
use FILL  FILL_2__3159_
timestamp 1701859473
transform 1 0 270 0 1 4430
box -12 -8 32 272
use FILL  FILL_2__3160_
timestamp 1701859473
transform -1 0 510 0 1 4430
box -12 -8 32 272
use FILL  FILL_2__3161_
timestamp 1701859473
transform 1 0 4150 0 -1 7030
box -12 -8 32 272
use FILL  FILL_2__3162_
timestamp 1701859473
transform -1 0 4390 0 -1 7030
box -12 -8 32 272
use FILL  FILL_2__3163_
timestamp 1701859473
transform 1 0 4610 0 -1 7030
box -12 -8 32 272
use FILL  FILL_2__3164_
timestamp 1701859473
transform 1 0 4850 0 1 7030
box -12 -8 32 272
use FILL  FILL_2__3165_
timestamp 1701859473
transform 1 0 4110 0 1 7550
box -12 -8 32 272
use FILL  FILL_2__3166_
timestamp 1701859473
transform -1 0 4350 0 1 7550
box -12 -8 32 272
use FILL  FILL_2__3167_
timestamp 1701859473
transform 1 0 4830 0 -1 10150
box -12 -8 32 272
use FILL  FILL_2__3168_
timestamp 1701859473
transform 1 0 5030 0 -1 10150
box -12 -8 32 272
use FILL  FILL_2__3169_
timestamp 1701859473
transform -1 0 3670 0 -1 10670
box -12 -8 32 272
use FILL  FILL_2__3170_
timestamp 1701859473
transform -1 0 3890 0 -1 10670
box -12 -8 32 272
use FILL  FILL_2__3171_
timestamp 1701859473
transform 1 0 4310 0 -1 10670
box -12 -8 32 272
use FILL  FILL_2__3172_
timestamp 1701859473
transform -1 0 4550 0 -1 10670
box -12 -8 32 272
use FILL  FILL_2__3173_
timestamp 1701859473
transform 1 0 4150 0 1 10150
box -12 -8 32 272
use FILL  FILL_2__3174_
timestamp 1701859473
transform -1 0 4390 0 1 10150
box -12 -8 32 272
use FILL  FILL_2__3175_
timestamp 1701859473
transform 1 0 5490 0 1 10150
box -12 -8 32 272
use FILL  FILL_2__3176_
timestamp 1701859473
transform 1 0 5250 0 1 10150
box -12 -8 32 272
use FILL  FILL_2__3177_
timestamp 1701859473
transform -1 0 1730 0 -1 5990
box -12 -8 32 272
use FILL  FILL_2__3178_
timestamp 1701859473
transform 1 0 2170 0 -1 5990
box -12 -8 32 272
use FILL  FILL_2__3179_
timestamp 1701859473
transform -1 0 1450 0 1 6510
box -12 -8 32 272
use FILL  FILL_2__3180_
timestamp 1701859473
transform -1 0 1670 0 1 6510
box -12 -8 32 272
use FILL  FILL_2__3181_
timestamp 1701859473
transform -1 0 530 0 -1 6510
box -12 -8 32 272
use FILL  FILL_2__3182_
timestamp 1701859473
transform -1 0 930 0 -1 6510
box -12 -8 32 272
use FILL  FILL_2__3183_
timestamp 1701859473
transform 1 0 290 0 1 8070
box -12 -8 32 272
use FILL  FILL_2__3184_
timestamp 1701859473
transform -1 0 530 0 1 8070
box -12 -8 32 272
use FILL  FILL_2__3185_
timestamp 1701859473
transform -1 0 70 0 -1 8590
box -12 -8 32 272
use FILL  FILL_2__3186_
timestamp 1701859473
transform -1 0 70 0 1 8070
box -12 -8 32 272
use FILL  FILL_2__3187_
timestamp 1701859473
transform 1 0 690 0 -1 9110
box -12 -8 32 272
use FILL  FILL_2__3188_
timestamp 1701859473
transform 1 0 910 0 -1 9110
box -12 -8 32 272
use FILL  FILL_2__3189_
timestamp 1701859473
transform 1 0 2090 0 -1 9630
box -12 -8 32 272
use FILL  FILL_2__3190_
timestamp 1701859473
transform 1 0 2330 0 1 9110
box -12 -8 32 272
use FILL  FILL_2__3191_
timestamp 1701859473
transform 1 0 1390 0 -1 9110
box -12 -8 32 272
use FILL  FILL_2__3192_
timestamp 1701859473
transform -1 0 1630 0 -1 9110
box -12 -8 32 272
use FILL  FILL_2__3324_
timestamp 1701859473
transform 1 0 5570 0 1 8070
box -12 -8 32 272
use FILL  FILL_2__3325_
timestamp 1701859473
transform -1 0 6290 0 1 8070
box -12 -8 32 272
use FILL  FILL_2__3326_
timestamp 1701859473
transform -1 0 6190 0 -1 8070
box -12 -8 32 272
use FILL  FILL_2__3327_
timestamp 1701859473
transform -1 0 6150 0 -1 8590
box -12 -8 32 272
use FILL  FILL_2__3328_
timestamp 1701859473
transform -1 0 6050 0 1 8070
box -12 -8 32 272
use FILL  FILL_2__3329_
timestamp 1701859473
transform 1 0 5810 0 1 8070
box -12 -8 32 272
use FILL  FILL_2__3330_
timestamp 1701859473
transform -1 0 6990 0 1 8590
box -12 -8 32 272
use FILL  FILL_2__3331_
timestamp 1701859473
transform 1 0 7270 0 -1 8590
box -12 -8 32 272
use FILL  FILL_2__3332_
timestamp 1701859473
transform 1 0 6990 0 -1 8590
box -12 -8 32 272
use FILL  FILL_2__3333_
timestamp 1701859473
transform 1 0 10190 0 1 8590
box -12 -8 32 272
use FILL  FILL_2__3334_
timestamp 1701859473
transform 1 0 9310 0 1 8590
box -12 -8 32 272
use FILL  FILL_2__3335_
timestamp 1701859473
transform 1 0 7850 0 -1 10150
box -12 -8 32 272
use FILL  FILL_2__3336_
timestamp 1701859473
transform -1 0 6690 0 1 9630
box -12 -8 32 272
use FILL  FILL_2__3337_
timestamp 1701859473
transform -1 0 6210 0 1 9630
box -12 -8 32 272
use FILL  FILL_2__3338_
timestamp 1701859473
transform 1 0 7170 0 -1 10150
box -12 -8 32 272
use FILL  FILL_2__3339_
timestamp 1701859473
transform -1 0 8050 0 1 10150
box -12 -8 32 272
use FILL  FILL_2__3340_
timestamp 1701859473
transform 1 0 7810 0 1 10150
box -12 -8 32 272
use FILL  FILL_2__3341_
timestamp 1701859473
transform 1 0 7570 0 1 10150
box -12 -8 32 272
use FILL  FILL_2__3342_
timestamp 1701859473
transform 1 0 6790 0 -1 11190
box -12 -8 32 272
use FILL  FILL_2__3343_
timestamp 1701859473
transform -1 0 7390 0 -1 10150
box -12 -8 32 272
use FILL  FILL_2__3344_
timestamp 1701859473
transform 1 0 7610 0 -1 10150
box -12 -8 32 272
use FILL  FILL_2__3345_
timestamp 1701859473
transform -1 0 8990 0 1 9630
box -12 -8 32 272
use FILL  FILL_2__3346_
timestamp 1701859473
transform 1 0 8510 0 1 10150
box -12 -8 32 272
use FILL  FILL_2__3347_
timestamp 1701859473
transform -1 0 8290 0 1 10150
box -12 -8 32 272
use FILL  FILL_2__3348_
timestamp 1701859473
transform 1 0 9110 0 -1 10670
box -12 -8 32 272
use FILL  FILL_2__3349_
timestamp 1701859473
transform 1 0 7850 0 1 9630
box -12 -8 32 272
use FILL  FILL_2__3350_
timestamp 1701859473
transform 1 0 7550 0 -1 8590
box -12 -8 32 272
use FILL  FILL_2__3351_
timestamp 1701859473
transform -1 0 7730 0 1 8590
box -12 -8 32 272
use FILL  FILL_2__3352_
timestamp 1701859473
transform -1 0 8190 0 -1 9110
box -12 -8 32 272
use FILL  FILL_2__3353_
timestamp 1701859473
transform 1 0 8070 0 -1 10150
box -12 -8 32 272
use FILL  FILL_2__3354_
timestamp 1701859473
transform 1 0 7750 0 -1 10670
box -12 -8 32 272
use FILL  FILL_2__3355_
timestamp 1701859473
transform -1 0 7530 0 -1 10670
box -12 -8 32 272
use FILL  FILL_2__3356_
timestamp 1701859473
transform 1 0 7310 0 -1 10670
box -12 -8 32 272
use FILL  FILL_2__3357_
timestamp 1701859473
transform 1 0 7130 0 1 10670
box -12 -8 32 272
use FILL  FILL_2__3358_
timestamp 1701859473
transform 1 0 7390 0 1 10670
box -12 -8 32 272
use FILL  FILL_2__3359_
timestamp 1701859473
transform 1 0 7630 0 1 10670
box -12 -8 32 272
use FILL  FILL_2__3360_
timestamp 1701859473
transform -1 0 7890 0 1 10670
box -12 -8 32 272
use FILL  FILL_2__3361_
timestamp 1701859473
transform 1 0 8910 0 -1 10670
box -12 -8 32 272
use FILL  FILL_2__3362_
timestamp 1701859473
transform 1 0 7970 0 -1 10670
box -12 -8 32 272
use FILL  FILL_2__3363_
timestamp 1701859473
transform 1 0 8090 0 1 10670
box -12 -8 32 272
use FILL  FILL_2__3364_
timestamp 1701859473
transform 1 0 7930 0 -1 11190
box -12 -8 32 272
use FILL  FILL_2__3365_
timestamp 1701859473
transform -1 0 7470 0 -1 11190
box -12 -8 32 272
use FILL  FILL_2__3366_
timestamp 1701859473
transform 1 0 6990 0 -1 11190
box -12 -8 32 272
use FILL  FILL_2__3367_
timestamp 1701859473
transform 1 0 6870 0 1 10670
box -12 -8 32 272
use FILL  FILL_2__3368_
timestamp 1701859473
transform 1 0 7210 0 -1 11190
box -12 -8 32 272
use FILL  FILL_2__3369_
timestamp 1701859473
transform 1 0 7690 0 -1 11190
box -12 -8 32 272
use FILL  FILL_2__3370_
timestamp 1701859473
transform 1 0 8210 0 -1 10670
box -12 -8 32 272
use FILL  FILL_2__3371_
timestamp 1701859473
transform 1 0 8310 0 1 10670
box -12 -8 32 272
use FILL  FILL_2__3372_
timestamp 1701859473
transform 1 0 9490 0 1 10670
box -12 -8 32 272
use FILL  FILL_2__3373_
timestamp 1701859473
transform -1 0 6590 0 -1 11190
box -12 -8 32 272
use FILL  FILL_2__3374_
timestamp 1701859473
transform 1 0 5690 0 1 10670
box -12 -8 32 272
use FILL  FILL_2__3375_
timestamp 1701859473
transform -1 0 5950 0 1 10670
box -12 -8 32 272
use FILL  FILL_2__3376_
timestamp 1701859473
transform -1 0 6170 0 1 10670
box -12 -8 32 272
use FILL  FILL_2__3377_
timestamp 1701859473
transform 1 0 6410 0 1 10670
box -12 -8 32 272
use FILL  FILL_2__3378_
timestamp 1701859473
transform 1 0 6350 0 -1 11190
box -12 -8 32 272
use FILL  FILL_2__3379_
timestamp 1701859473
transform 1 0 8670 0 -1 10670
box -12 -8 32 272
use FILL  FILL_2__3380_
timestamp 1701859473
transform 1 0 8790 0 1 10670
box -12 -8 32 272
use FILL  FILL_2__3381_
timestamp 1701859473
transform -1 0 6670 0 1 10670
box -12 -8 32 272
use FILL  FILL_2__3382_
timestamp 1701859473
transform 1 0 6130 0 -1 10670
box -12 -8 32 272
use FILL  FILL_2__3383_
timestamp 1701859473
transform -1 0 6390 0 -1 10670
box -12 -8 32 272
use FILL  FILL_2__3384_
timestamp 1701859473
transform -1 0 6830 0 -1 10670
box -12 -8 32 272
use FILL  FILL_2__3385_
timestamp 1701859473
transform 1 0 6590 0 -1 10670
box -12 -8 32 272
use FILL  FILL_2__3386_
timestamp 1701859473
transform 1 0 7070 0 -1 10670
box -12 -8 32 272
use FILL  FILL_2__3387_
timestamp 1701859473
transform 1 0 8430 0 -1 10670
box -12 -8 32 272
use FILL  FILL_2__3388_
timestamp 1701859473
transform 1 0 8550 0 1 10670
box -12 -8 32 272
use FILL  FILL_2__3389_
timestamp 1701859473
transform 1 0 10210 0 -1 10670
box -12 -8 32 272
use FILL  FILL_2__3390_
timestamp 1701859473
transform 1 0 9770 0 -1 10670
box -12 -8 32 272
use FILL  FILL_2__3391_
timestamp 1701859473
transform 1 0 9970 0 -1 10670
box -12 -8 32 272
use FILL  FILL_2__3392_
timestamp 1701859473
transform 1 0 10430 0 -1 10670
box -12 -8 32 272
use FILL  FILL_2__3393_
timestamp 1701859473
transform -1 0 11170 0 -1 10150
box -12 -8 32 272
use FILL  FILL_2__3394_
timestamp 1701859473
transform 1 0 7350 0 1 10150
box -12 -8 32 272
use FILL  FILL_2__3395_
timestamp 1701859473
transform 1 0 6410 0 1 10150
box -12 -8 32 272
use FILL  FILL_2__3396_
timestamp 1701859473
transform -1 0 6670 0 1 10150
box -12 -8 32 272
use FILL  FILL_2__3397_
timestamp 1701859473
transform -1 0 6990 0 -1 10150
box -12 -8 32 272
use FILL  FILL_2__3398_
timestamp 1701859473
transform 1 0 6270 0 -1 10150
box -12 -8 32 272
use FILL  FILL_2__3399_
timestamp 1701859473
transform -1 0 6750 0 -1 10150
box -12 -8 32 272
use FILL  FILL_2__3400_
timestamp 1701859473
transform -1 0 6930 0 1 10150
box -12 -8 32 272
use FILL  FILL_2__3401_
timestamp 1701859473
transform 1 0 7110 0 1 10150
box -12 -8 32 272
use FILL  FILL_2__3402_
timestamp 1701859473
transform -1 0 9050 0 1 10150
box -12 -8 32 272
use FILL  FILL_2__3403_
timestamp 1701859473
transform 1 0 9490 0 1 10150
box -12 -8 32 272
use FILL  FILL_2__3404_
timestamp 1701859473
transform -1 0 5750 0 1 9630
box -12 -8 32 272
use FILL  FILL_2__3405_
timestamp 1701859473
transform -1 0 6030 0 -1 10150
box -12 -8 32 272
use FILL  FILL_2__3406_
timestamp 1701859473
transform 1 0 6390 0 -1 9630
box -12 -8 32 272
use FILL  FILL_2__3407_
timestamp 1701859473
transform -1 0 6610 0 -1 9630
box -12 -8 32 272
use FILL  FILL_2__3408_
timestamp 1701859473
transform 1 0 6870 0 1 9630
box -12 -8 32 272
use FILL  FILL_2__3409_
timestamp 1701859473
transform -1 0 6490 0 -1 10150
box -12 -8 32 272
use FILL  FILL_2__3410_
timestamp 1701859473
transform 1 0 9230 0 -1 10150
box -12 -8 32 272
use FILL  FILL_2__3411_
timestamp 1701859473
transform 1 0 9250 0 1 10150
box -12 -8 32 272
use FILL  FILL_2__3412_
timestamp 1701859473
transform 1 0 9970 0 1 10150
box -12 -8 32 272
use FILL  FILL_2__3413_
timestamp 1701859473
transform -1 0 5990 0 1 9630
box -12 -8 32 272
use FILL  FILL_2__3414_
timestamp 1701859473
transform 1 0 8130 0 1 9110
box -12 -8 32 272
use FILL  FILL_2__3415_
timestamp 1701859473
transform 1 0 6410 0 1 9630
box -12 -8 32 272
use FILL  FILL_2__3416_
timestamp 1701859473
transform 1 0 7250 0 1 8590
box -12 -8 32 272
use FILL  FILL_2__3417_
timestamp 1701859473
transform 1 0 7330 0 -1 9110
box -12 -8 32 272
use FILL  FILL_2__3418_
timestamp 1701859473
transform -1 0 7470 0 -1 9630
box -12 -8 32 272
use FILL  FILL_2__3419_
timestamp 1701859473
transform 1 0 7230 0 -1 9630
box -12 -8 32 272
use FILL  FILL_2__3420_
timestamp 1701859473
transform -1 0 6810 0 -1 9630
box -12 -8 32 272
use FILL  FILL_2__3421_
timestamp 1701859473
transform -1 0 7030 0 -1 9630
box -12 -8 32 272
use FILL  FILL_2__3422_
timestamp 1701859473
transform -1 0 7130 0 1 9630
box -12 -8 32 272
use FILL  FILL_2__3423_
timestamp 1701859473
transform -1 0 8190 0 -1 9630
box -12 -8 32 272
use FILL  FILL_2__3424_
timestamp 1701859473
transform -1 0 7710 0 -1 9630
box -12 -8 32 272
use FILL  FILL_2__3425_
timestamp 1701859473
transform -1 0 7370 0 1 9630
box -12 -8 32 272
use FILL  FILL_2__3426_
timestamp 1701859473
transform -1 0 9010 0 -1 10150
box -12 -8 32 272
use FILL  FILL_2__3427_
timestamp 1701859473
transform 1 0 8770 0 -1 10150
box -12 -8 32 272
use FILL  FILL_2__3428_
timestamp 1701859473
transform 1 0 7450 0 1 8590
box -12 -8 32 272
use FILL  FILL_2__3429_
timestamp 1701859473
transform 1 0 7530 0 -1 9110
box -12 -8 32 272
use FILL  FILL_2__3430_
timestamp 1701859473
transform -1 0 7750 0 -1 9110
box -12 -8 32 272
use FILL  FILL_2__3431_
timestamp 1701859473
transform 1 0 7670 0 1 9110
box -12 -8 32 272
use FILL  FILL_2__3432_
timestamp 1701859473
transform 1 0 7910 0 1 9110
box -12 -8 32 272
use FILL  FILL_2__3433_
timestamp 1701859473
transform -1 0 7950 0 -1 9630
box -12 -8 32 272
use FILL  FILL_2__3434_
timestamp 1701859473
transform 1 0 7590 0 1 9630
box -12 -8 32 272
use FILL  FILL_2__3435_
timestamp 1701859473
transform 1 0 10210 0 1 10150
box -12 -8 32 272
use FILL  FILL_2__3436_
timestamp 1701859473
transform -1 0 10210 0 -1 10150
box -12 -8 32 272
use FILL  FILL_2__3437_
timestamp 1701859473
transform 1 0 10650 0 1 10150
box -12 -8 32 272
use FILL  FILL_2__3438_
timestamp 1701859473
transform 1 0 10430 0 1 10150
box -12 -8 32 272
use FILL  FILL_2__3439_
timestamp 1701859473
transform 1 0 10870 0 1 10150
box -12 -8 32 272
use FILL  FILL_2__3440_
timestamp 1701859473
transform -1 0 10690 0 -1 10150
box -12 -8 32 272
use FILL  FILL_2__3441_
timestamp 1701859473
transform -1 0 10550 0 1 9630
box -12 -8 32 272
use FILL  FILL_2__3442_
timestamp 1701859473
transform -1 0 10430 0 -1 10150
box -12 -8 32 272
use FILL  FILL_2__3443_
timestamp 1701859473
transform -1 0 10990 0 1 9630
box -12 -8 32 272
use FILL  FILL_2__3444_
timestamp 1701859473
transform -1 0 8390 0 -1 9630
box -12 -8 32 272
use FILL  FILL_2__3445_
timestamp 1701859473
transform -1 0 8090 0 1 9630
box -12 -8 32 272
use FILL  FILL_2__3446_
timestamp 1701859473
transform 1 0 8530 0 1 9630
box -12 -8 32 272
use FILL  FILL_2__3447_
timestamp 1701859473
transform 1 0 8310 0 1 9630
box -12 -8 32 272
use FILL  FILL_2__3448_
timestamp 1701859473
transform -1 0 8750 0 1 9630
box -12 -8 32 272
use FILL  FILL_2__3449_
timestamp 1701859473
transform -1 0 9790 0 1 10150
box -12 -8 32 272
use FILL  FILL_2__3450_
timestamp 1701859473
transform -1 0 9750 0 -1 10150
box -12 -8 32 272
use FILL  FILL_2__3451_
timestamp 1701859473
transform 1 0 9470 0 -1 10150
box -12 -8 32 272
use FILL  FILL_2__3452_
timestamp 1701859473
transform -1 0 9210 0 1 9630
box -12 -8 32 272
use FILL  FILL_2__3453_
timestamp 1701859473
transform -1 0 9970 0 -1 10150
box -12 -8 32 272
use FILL  FILL_2__3454_
timestamp 1701859473
transform 1 0 9410 0 1 9630
box -12 -8 32 272
use FILL  FILL_2__3455_
timestamp 1701859473
transform 1 0 9630 0 1 9630
box -12 -8 32 272
use FILL  FILL_2__3456_
timestamp 1701859473
transform -1 0 10330 0 1 9630
box -12 -8 32 272
use FILL  FILL_2__3457_
timestamp 1701859473
transform -1 0 9870 0 1 9630
box -12 -8 32 272
use FILL  FILL_2__3458_
timestamp 1701859473
transform -1 0 10110 0 1 9630
box -12 -8 32 272
use FILL  FILL_2__3459_
timestamp 1701859473
transform -1 0 10250 0 -1 9630
box -12 -8 32 272
use FILL  FILL_2__3460_
timestamp 1701859473
transform 1 0 10910 0 -1 10150
box -12 -8 32 272
use FILL  FILL_2__3461_
timestamp 1701859473
transform -1 0 11150 0 -1 9630
box -12 -8 32 272
use FILL  FILL_2__3462_
timestamp 1701859473
transform -1 0 10690 0 -1 9630
box -12 -8 32 272
use FILL  FILL_2__3463_
timestamp 1701859473
transform 1 0 10370 0 -1 11190
box -12 -8 32 272
use FILL  FILL_2__3464_
timestamp 1701859473
transform 1 0 9710 0 -1 11190
box -12 -8 32 272
use FILL  FILL_2__3465_
timestamp 1701859473
transform 1 0 9950 0 -1 11190
box -12 -8 32 272
use FILL  FILL_2__3466_
timestamp 1701859473
transform 1 0 10130 0 -1 11190
box -12 -8 32 272
use FILL  FILL_2__3467_
timestamp 1701859473
transform -1 0 11110 0 1 10670
box -12 -8 32 272
use FILL  FILL_2__3468_
timestamp 1701859473
transform 1 0 10610 0 1 10670
box -12 -8 32 272
use FILL  FILL_2__3469_
timestamp 1701859473
transform 1 0 9330 0 -1 10670
box -12 -8 32 272
use FILL  FILL_2__3470_
timestamp 1701859473
transform 1 0 9570 0 -1 10670
box -12 -8 32 272
use FILL  FILL_2__3471_
timestamp 1701859473
transform 1 0 9710 0 1 10670
box -12 -8 32 272
use FILL  FILL_2__3472_
timestamp 1701859473
transform -1 0 9970 0 1 10670
box -12 -8 32 272
use FILL  FILL_2__3473_
timestamp 1701859473
transform 1 0 8590 0 -1 11190
box -12 -8 32 272
use FILL  FILL_2__3474_
timestamp 1701859473
transform 1 0 8150 0 -1 11190
box -12 -8 32 272
use FILL  FILL_2__3475_
timestamp 1701859473
transform 1 0 8390 0 -1 11190
box -12 -8 32 272
use FILL  FILL_2__3476_
timestamp 1701859473
transform -1 0 8830 0 -1 11190
box -12 -8 32 272
use FILL  FILL_2__3477_
timestamp 1701859473
transform 1 0 9050 0 -1 11190
box -12 -8 32 272
use FILL  FILL_2__3478_
timestamp 1701859473
transform 1 0 9030 0 1 10670
box -12 -8 32 272
use FILL  FILL_2__3479_
timestamp 1701859473
transform 1 0 8310 0 -1 10150
box -12 -8 32 272
use FILL  FILL_2__3480_
timestamp 1701859473
transform -1 0 8570 0 -1 10150
box -12 -8 32 272
use FILL  FILL_2__3481_
timestamp 1701859473
transform -1 0 8350 0 1 9110
box -12 -8 32 272
use FILL  FILL_2__3482_
timestamp 1701859473
transform -1 0 8570 0 1 9110
box -12 -8 32 272
use FILL  FILL_2__3483_
timestamp 1701859473
transform 1 0 8750 0 1 10150
box -12 -8 32 272
use FILL  FILL_2__3484_
timestamp 1701859473
transform -1 0 10050 0 -1 9630
box -12 -8 32 272
use FILL  FILL_2__3485_
timestamp 1701859473
transform 1 0 11070 0 1 10150
box -12 -8 32 272
use FILL  FILL_2__3486_
timestamp 1701859473
transform 1 0 10410 0 1 9110
box -12 -8 32 272
use FILL  FILL_2__3487_
timestamp 1701859473
transform 1 0 10450 0 -1 9630
box -12 -8 32 272
use FILL  FILL_2__3488_
timestamp 1701859473
transform -1 0 10750 0 1 9630
box -12 -8 32 272
use FILL  FILL_2__3489_
timestamp 1701859473
transform 1 0 10590 0 -1 11190
box -12 -8 32 272
use FILL  FILL_2__3490_
timestamp 1701859473
transform 1 0 11050 0 -1 11190
box -12 -8 32 272
use FILL  FILL_2__3491_
timestamp 1701859473
transform -1 0 10850 0 -1 11190
box -12 -8 32 272
use FILL  FILL_2__3492_
timestamp 1701859473
transform -1 0 10410 0 1 10670
box -12 -8 32 272
use FILL  FILL_2__3493_
timestamp 1701859473
transform -1 0 10190 0 1 10670
box -12 -8 32 272
use FILL  FILL_2__3494_
timestamp 1701859473
transform 1 0 9290 0 1 10670
box -12 -8 32 272
use FILL  FILL_2__3495_
timestamp 1701859473
transform -1 0 9490 0 -1 11190
box -12 -8 32 272
use FILL  FILL_2__3496_
timestamp 1701859473
transform 1 0 9250 0 -1 11190
box -12 -8 32 272
use FILL  FILL_2__3497_
timestamp 1701859473
transform -1 0 9350 0 -1 9630
box -12 -8 32 272
use FILL  FILL_2__3498_
timestamp 1701859473
transform -1 0 8850 0 1 9110
box -12 -8 32 272
use FILL  FILL_2__3499_
timestamp 1701859473
transform 1 0 8370 0 -1 9110
box -12 -8 32 272
use FILL  FILL_2__3500_
timestamp 1701859473
transform 1 0 9750 0 1 9110
box -12 -8 32 272
use FILL  FILL_2__3501_
timestamp 1701859473
transform -1 0 9990 0 1 9110
box -12 -8 32 272
use FILL  FILL_2__3502_
timestamp 1701859473
transform -1 0 8250 0 -1 8590
box -12 -8 32 272
use FILL  FILL_2__3503_
timestamp 1701859473
transform -1 0 8630 0 -1 9630
box -12 -8 32 272
use FILL  FILL_2__3504_
timestamp 1701859473
transform 1 0 8850 0 -1 9630
box -12 -8 32 272
use FILL  FILL_2__3505_
timestamp 1701859473
transform -1 0 9110 0 -1 9630
box -12 -8 32 272
use FILL  FILL_2__3506_
timestamp 1701859473
transform -1 0 8630 0 1 8590
box -12 -8 32 272
use FILL  FILL_2__3507_
timestamp 1701859473
transform 1 0 10710 0 -1 9110
box -12 -8 32 272
use FILL  FILL_2__3508_
timestamp 1701859473
transform 1 0 10470 0 -1 9110
box -12 -8 32 272
use FILL  FILL_2__3509_
timestamp 1701859473
transform 1 0 8410 0 1 8590
box -12 -8 32 272
use FILL  FILL_2__3510_
timestamp 1701859473
transform -1 0 8870 0 1 8590
box -12 -8 32 272
use FILL  FILL_2__3511_
timestamp 1701859473
transform 1 0 9930 0 -1 270
box -12 -8 32 272
use FILL  FILL_2__3512_
timestamp 1701859473
transform 1 0 10930 0 -1 9110
box -12 -8 32 272
use FILL  FILL_2__3513_
timestamp 1701859473
transform 1 0 10910 0 -1 9630
box -12 -8 32 272
use FILL  FILL_2__3514_
timestamp 1701859473
transform 1 0 10870 0 1 10670
box -12 -8 32 272
use FILL  FILL_2__3515_
timestamp 1701859473
transform -1 0 10670 0 -1 10670
box -12 -8 32 272
use FILL  FILL_2__3516_
timestamp 1701859473
transform 1 0 10890 0 -1 10670
box -12 -8 32 272
use FILL  FILL_2__3517_
timestamp 1701859473
transform 1 0 9570 0 -1 9630
box -12 -8 32 272
use FILL  FILL_2__3518_
timestamp 1701859473
transform 1 0 9790 0 -1 9630
box -12 -8 32 272
use FILL  FILL_2__3519_
timestamp 1701859473
transform 1 0 9070 0 1 9110
box -12 -8 32 272
use FILL  FILL_2__3520_
timestamp 1701859473
transform -1 0 9310 0 1 9110
box -12 -8 32 272
use FILL  FILL_2__3521_
timestamp 1701859473
transform 1 0 6550 0 1 8590
box -12 -8 32 272
use FILL  FILL_2__3522_
timestamp 1701859473
transform 1 0 7950 0 -1 9110
box -12 -8 32 272
use FILL  FILL_2__3523_
timestamp 1701859473
transform 1 0 6750 0 1 8590
box -12 -8 32 272
use FILL  FILL_2__3524_
timestamp 1701859473
transform 1 0 7470 0 1 9110
box -12 -8 32 272
use FILL  FILL_2__3525_
timestamp 1701859473
transform 1 0 7010 0 1 9110
box -12 -8 32 272
use FILL  FILL_2__3526_
timestamp 1701859473
transform -1 0 7250 0 1 9110
box -12 -8 32 272
use FILL  FILL_2__3539_
timestamp 1701859473
transform 1 0 11110 0 -1 7030
box -12 -8 32 272
use FILL  FILL_2__3540_
timestamp 1701859473
transform 1 0 4610 0 1 10670
box -12 -8 32 272
use FILL  FILL_2__3541_
timestamp 1701859473
transform -1 0 70 0 1 5990
box -12 -8 32 272
use FILL  FILL_2__3542_
timestamp 1701859473
transform -1 0 70 0 -1 8070
box -12 -8 32 272
use FILL  FILL_2__3543_
timestamp 1701859473
transform -1 0 70 0 1 8590
box -12 -8 32 272
use FILL  FILL_2__3544_
timestamp 1701859473
transform -1 0 70 0 1 9110
box -12 -8 32 272
use FILL  FILL_2__3545_
timestamp 1701859473
transform -1 0 1910 0 -1 11190
box -12 -8 32 272
use FILL  FILL_2__3546_
timestamp 1701859473
transform -1 0 530 0 1 9110
box -12 -8 32 272
use FILL  FILL_2__3547_
timestamp 1701859473
transform 1 0 4650 0 -1 11190
box -12 -8 32 272
use FILL  FILL_2__3548_
timestamp 1701859473
transform 1 0 5250 0 1 10670
box -12 -8 32 272
use FILL  FILL_2__3549_
timestamp 1701859473
transform -1 0 4250 0 -1 11190
box -12 -8 32 272
use FILL  FILL_2__3550_
timestamp 1701859473
transform -1 0 5090 0 -1 11190
box -12 -8 32 272
use FILL  FILL_2__3551_
timestamp 1701859473
transform 1 0 5490 0 -1 11190
box -12 -8 32 272
use FILL  FILL_2__3552_
timestamp 1701859473
transform 1 0 5270 0 -1 11190
box -12 -8 32 272
use FILL  FILL_2__3553_
timestamp 1701859473
transform -1 0 70 0 -1 5990
box -12 -8 32 272
use FILL  FILL_2__3554_
timestamp 1701859473
transform -1 0 270 0 1 7030
box -12 -8 32 272
use FILL  FILL_2__3555_
timestamp 1701859473
transform -1 0 5050 0 1 10670
box -12 -8 32 272
use FILL  FILL_2__3556_
timestamp 1701859473
transform 1 0 6190 0 1 10150
box -12 -8 32 272
use FILL  FILL_2__3557_
timestamp 1701859473
transform -1 0 5730 0 -1 11190
box -12 -8 32 272
use FILL  FILL_2__3558_
timestamp 1701859473
transform 1 0 6130 0 -1 11190
box -12 -8 32 272
use FILL  FILL_2__3559_
timestamp 1701859473
transform -1 0 4790 0 -1 10670
box -12 -8 32 272
use FILL  FILL_2__3560_
timestamp 1701859473
transform 1 0 5470 0 1 10670
box -12 -8 32 272
use FILL  FILL_2__3561_
timestamp 1701859473
transform 1 0 5910 0 -1 11190
box -12 -8 32 272
use FILL  FILL_2__3562_
timestamp 1701859473
transform 1 0 5710 0 1 10150
box -12 -8 32 272
use FILL  FILL_2__3563_
timestamp 1701859473
transform 1 0 5170 0 1 3390
box -12 -8 32 272
use FILL  FILL_2_BUFX2_insert0
timestamp 1701859473
transform 1 0 5790 0 -1 10150
box -12 -8 32 272
use FILL  FILL_2_BUFX2_insert1
timestamp 1701859473
transform 1 0 6550 0 1 2350
box -12 -8 32 272
use FILL  FILL_2_BUFX2_insert2
timestamp 1701859473
transform 1 0 5390 0 -1 1830
box -12 -8 32 272
use FILL  FILL_2_BUFX2_insert3
timestamp 1701859473
transform -1 0 530 0 -1 5470
box -12 -8 32 272
use FILL  FILL_2_BUFX2_insert4
timestamp 1701859473
transform 1 0 3270 0 1 4950
box -12 -8 32 272
use FILL  FILL_2_BUFX2_insert5
timestamp 1701859473
transform 1 0 1330 0 -1 1830
box -12 -8 32 272
use FILL  FILL_2_BUFX2_insert6
timestamp 1701859473
transform -1 0 70 0 -1 11190
box -12 -8 32 272
use FILL  FILL_2_BUFX2_insert7
timestamp 1701859473
transform 1 0 1630 0 1 10670
box -12 -8 32 272
use FILL  FILL_2_BUFX2_insert8
timestamp 1701859473
transform 1 0 1590 0 1 1830
box -12 -8 32 272
use FILL  FILL_2_BUFX2_insert9
timestamp 1701859473
transform 1 0 1890 0 -1 3910
box -12 -8 32 272
use FILL  FILL_2_BUFX2_insert10
timestamp 1701859473
transform 1 0 1710 0 -1 4430
box -12 -8 32 272
use FILL  FILL_2_BUFX2_insert11
timestamp 1701859473
transform -1 0 1690 0 -1 3910
box -12 -8 32 272
use FILL  FILL_2_BUFX2_insert12
timestamp 1701859473
transform -1 0 1470 0 -1 3910
box -12 -8 32 272
use FILL  FILL_2_BUFX2_insert13
timestamp 1701859473
transform -1 0 1370 0 -1 1310
box -12 -8 32 272
use FILL  FILL_2_BUFX2_insert14
timestamp 1701859473
transform -1 0 3610 0 1 3390
box -12 -8 32 272
use FILL  FILL_2_BUFX2_insert15
timestamp 1701859473
transform 1 0 4490 0 -1 5470
box -12 -8 32 272
use FILL  FILL_2_BUFX2_insert16
timestamp 1701859473
transform 1 0 1290 0 -1 4950
box -12 -8 32 272
use FILL  FILL_2_BUFX2_insert17
timestamp 1701859473
transform 1 0 3570 0 1 1310
box -12 -8 32 272
use FILL  FILL_2_BUFX2_insert18
timestamp 1701859473
transform -1 0 9710 0 1 2350
box -12 -8 32 272
use FILL  FILL_2_BUFX2_insert19
timestamp 1701859473
transform -1 0 8450 0 -1 790
box -12 -8 32 272
use FILL  FILL_2_BUFX2_insert20
timestamp 1701859473
transform 1 0 9910 0 1 2350
box -12 -8 32 272
use FILL  FILL_2_BUFX2_insert21
timestamp 1701859473
transform -1 0 7750 0 -1 1310
box -12 -8 32 272
use FILL  FILL_2_BUFX2_insert22
timestamp 1701859473
transform -1 0 3150 0 -1 2870
box -12 -8 32 272
use FILL  FILL_2_BUFX2_insert23
timestamp 1701859473
transform -1 0 2690 0 -1 4950
box -12 -8 32 272
use FILL  FILL_2_BUFX2_insert24
timestamp 1701859473
transform -1 0 3590 0 -1 4430
box -12 -8 32 272
use FILL  FILL_2_BUFX2_insert25
timestamp 1701859473
transform 1 0 4330 0 1 4430
box -12 -8 32 272
use FILL  FILL_2_BUFX2_insert26
timestamp 1701859473
transform 1 0 4150 0 1 2870
box -12 -8 32 272
use FILL  FILL_2_BUFX2_insert27
timestamp 1701859473
transform 1 0 9550 0 1 4950
box -12 -8 32 272
use FILL  FILL_2_BUFX2_insert28
timestamp 1701859473
transform -1 0 7430 0 -1 5990
box -12 -8 32 272
use FILL  FILL_2_BUFX2_insert29
timestamp 1701859473
transform -1 0 1230 0 1 6510
box -12 -8 32 272
use FILL  FILL_2_BUFX2_insert30
timestamp 1701859473
transform -1 0 8730 0 -1 3910
box -12 -8 32 272
use FILL  FILL_2_BUFX2_insert31
timestamp 1701859473
transform -1 0 9510 0 1 3910
box -12 -8 32 272
use FILL  FILL_2_BUFX2_insert32
timestamp 1701859473
transform 1 0 5810 0 -1 3910
box -12 -8 32 272
use FILL  FILL_2_BUFX2_insert33
timestamp 1701859473
transform -1 0 9490 0 -1 4950
box -12 -8 32 272
use FILL  FILL_2_BUFX2_insert34
timestamp 1701859473
transform 1 0 5150 0 1 8590
box -12 -8 32 272
use FILL  FILL_2_BUFX2_insert35
timestamp 1701859473
transform -1 0 5910 0 1 7550
box -12 -8 32 272
use FILL  FILL_2_BUFX2_insert36
timestamp 1701859473
transform -1 0 1150 0 1 8590
box -12 -8 32 272
use FILL  FILL_2_BUFX2_insert37
timestamp 1701859473
transform -1 0 9530 0 1 8590
box -12 -8 32 272
use FILL  FILL_2_BUFX2_insert49
timestamp 1701859473
transform -1 0 2990 0 1 6510
box -12 -8 32 272
use FILL  FILL_2_BUFX2_insert50
timestamp 1701859473
transform 1 0 2290 0 -1 8590
box -12 -8 32 272
use FILL  FILL_2_BUFX2_insert51
timestamp 1701859473
transform 1 0 3150 0 -1 8590
box -12 -8 32 272
use FILL  FILL_2_BUFX2_insert52
timestamp 1701859473
transform 1 0 3330 0 1 5470
box -12 -8 32 272
use FILL  FILL_2_BUFX2_insert53
timestamp 1701859473
transform -1 0 11170 0 1 9110
box -12 -8 32 272
use FILL  FILL_2_BUFX2_insert54
timestamp 1701859473
transform -1 0 9110 0 1 8590
box -12 -8 32 272
use FILL  FILL_2_BUFX2_insert55
timestamp 1701859473
transform -1 0 9550 0 1 9110
box -12 -8 32 272
use FILL  FILL_2_BUFX2_insert56
timestamp 1701859473
transform -1 0 10210 0 1 9110
box -12 -8 32 272
use FILL  FILL_2_BUFX2_insert57
timestamp 1701859473
transform -1 0 11170 0 -1 2350
box -12 -8 32 272
use FILL  FILL_2_BUFX2_insert58
timestamp 1701859473
transform -1 0 8910 0 1 2870
box -12 -8 32 272
use FILL  FILL_2_BUFX2_insert59
timestamp 1701859473
transform -1 0 7490 0 1 1830
box -12 -8 32 272
use FILL  FILL_2_BUFX2_insert60
timestamp 1701859473
transform 1 0 10830 0 1 1830
box -12 -8 32 272
use FILL  FILL_2_BUFX2_insert61
timestamp 1701859473
transform -1 0 11110 0 1 2870
box -12 -8 32 272
use FILL  FILL_2_BUFX2_insert62
timestamp 1701859473
transform 1 0 2150 0 1 3910
box -12 -8 32 272
use FILL  FILL_2_BUFX2_insert63
timestamp 1701859473
transform 1 0 2070 0 1 3390
box -12 -8 32 272
use FILL  FILL_2_BUFX2_insert64
timestamp 1701859473
transform -1 0 1730 0 1 3910
box -12 -8 32 272
use FILL  FILL_2_BUFX2_insert65
timestamp 1701859473
transform -1 0 1670 0 1 3390
box -12 -8 32 272
use FILL  FILL_2_BUFX2_insert66
timestamp 1701859473
transform -1 0 4250 0 1 1310
box -12 -8 32 272
use FILL  FILL_2_BUFX2_insert67
timestamp 1701859473
transform -1 0 3550 0 -1 10150
box -12 -8 32 272
use FILL  FILL_2_BUFX2_insert68
timestamp 1701859473
transform -1 0 7110 0 1 2870
box -12 -8 32 272
use FILL  FILL_2_BUFX2_insert69
timestamp 1701859473
transform -1 0 5590 0 -1 3390
box -12 -8 32 272
use FILL  FILL_2_BUFX2_insert70
timestamp 1701859473
transform -1 0 3610 0 -1 1830
box -12 -8 32 272
use FILL  FILL_2_BUFX2_insert71
timestamp 1701859473
transform -1 0 7250 0 1 2350
box -12 -8 32 272
use FILL  FILL_2_BUFX2_insert72
timestamp 1701859473
transform -1 0 6430 0 1 1310
box -12 -8 32 272
use FILL  FILL_2_BUFX2_insert73
timestamp 1701859473
transform 1 0 3550 0 1 5470
box -12 -8 32 272
use FILL  FILL_2_BUFX2_insert74
timestamp 1701859473
transform 1 0 7510 0 -1 2350
box -12 -8 32 272
use FILL  FILL_2_BUFX2_insert75
timestamp 1701859473
transform 1 0 7530 0 1 2870
box -12 -8 32 272
use FILL  FILL_2_BUFX2_insert76
timestamp 1701859473
transform 1 0 7310 0 1 2870
box -12 -8 32 272
use FILL  FILL_2_BUFX2_insert77
timestamp 1701859473
transform -1 0 3370 0 -1 2870
box -12 -8 32 272
use FILL  FILL_2_BUFX2_insert78
timestamp 1701859473
transform 1 0 1870 0 -1 2870
box -12 -8 32 272
use FILL  FILL_2_BUFX2_insert79
timestamp 1701859473
transform -1 0 2110 0 -1 2870
box -12 -8 32 272
use FILL  FILL_2_BUFX2_insert80
timestamp 1701859473
transform 1 0 2350 0 1 4430
box -12 -8 32 272
use FILL  FILL_2_BUFX2_insert81
timestamp 1701859473
transform -1 0 1950 0 1 3910
box -12 -8 32 272
use FILL  FILL_2_BUFX2_insert82
timestamp 1701859473
transform -1 0 270 0 1 8590
box -12 -8 32 272
use FILL  FILL_2_BUFX2_insert83
timestamp 1701859473
transform 1 0 4150 0 -1 10150
box -12 -8 32 272
use FILL  FILL_2_BUFX2_insert84
timestamp 1701859473
transform 1 0 4110 0 -1 7550
box -12 -8 32 272
use FILL  FILL_2_BUFX2_insert85
timestamp 1701859473
transform -1 0 70 0 -1 6510
box -12 -8 32 272
use FILL  FILL_2_BUFX2_insert86
timestamp 1701859473
transform 1 0 1870 0 -1 10150
box -12 -8 32 272
use FILL  FILL_2_CLKBUF1_insert38
timestamp 1701859473
transform 1 0 2870 0 -1 7550
box -12 -8 32 272
use FILL  FILL_2_CLKBUF1_insert39
timestamp 1701859473
transform -1 0 4670 0 -1 6510
box -12 -8 32 272
use FILL  FILL_2_CLKBUF1_insert40
timestamp 1701859473
transform -1 0 970 0 -1 4950
box -12 -8 32 272
use FILL  FILL_2_CLKBUF1_insert41
timestamp 1701859473
transform -1 0 10630 0 -1 270
box -12 -8 32 272
use FILL  FILL_2_CLKBUF1_insert42
timestamp 1701859473
transform 1 0 9690 0 -1 4950
box -12 -8 32 272
use FILL  FILL_2_CLKBUF1_insert43
timestamp 1701859473
transform -1 0 11010 0 1 7030
box -12 -8 32 272
use FILL  FILL_2_CLKBUF1_insert44
timestamp 1701859473
transform -1 0 10750 0 1 4430
box -12 -8 32 272
use FILL  FILL_2_CLKBUF1_insert45
timestamp 1701859473
transform 1 0 5670 0 -1 6510
box -12 -8 32 272
use FILL  FILL_2_CLKBUF1_insert46
timestamp 1701859473
transform 1 0 3990 0 1 5990
box -12 -8 32 272
use FILL  FILL_2_CLKBUF1_insert47
timestamp 1701859473
transform -1 0 2110 0 1 7550
box -12 -8 32 272
use FILL  FILL_2_CLKBUF1_insert48
timestamp 1701859473
transform -1 0 10790 0 -1 7030
box -12 -8 32 272
use FILL  FILL_3__1668_
timestamp 1701859473
transform 1 0 6750 0 -1 3390
box -12 -8 32 272
use FILL  FILL_3__1669_
timestamp 1701859473
transform -1 0 6790 0 -1 790
box -12 -8 32 272
use FILL  FILL_3__1670_
timestamp 1701859473
transform 1 0 6570 0 -1 2870
box -12 -8 32 272
use FILL  FILL_3__1671_
timestamp 1701859473
transform -1 0 6370 0 -1 8590
box -12 -8 32 272
use FILL  FILL_3__1672_
timestamp 1701859473
transform 1 0 5930 0 -1 10670
box -12 -8 32 272
use FILL  FILL_3__1673_
timestamp 1701859473
transform 1 0 6330 0 1 8590
box -12 -8 32 272
use FILL  FILL_3__1674_
timestamp 1701859473
transform -1 0 6410 0 -1 9110
box -12 -8 32 272
use FILL  FILL_3__1675_
timestamp 1701859473
transform 1 0 70 0 -1 5470
box -12 -8 32 272
use FILL  FILL_3__1676_
timestamp 1701859473
transform -1 0 310 0 -1 5470
box -12 -8 32 272
use FILL  FILL_3__1677_
timestamp 1701859473
transform -1 0 550 0 1 5470
box -12 -8 32 272
use FILL  FILL_3__1678_
timestamp 1701859473
transform 1 0 70 0 -1 10670
box -12 -8 32 272
use FILL  FILL_3__1679_
timestamp 1701859473
transform -1 0 290 0 -1 11190
box -12 -8 32 272
use FILL  FILL_3__1680_
timestamp 1701859473
transform 1 0 270 0 -1 10670
box -12 -8 32 272
use FILL  FILL_3__1681_
timestamp 1701859473
transform -1 0 90 0 -1 7030
box -12 -8 32 272
use FILL  FILL_3__1682_
timestamp 1701859473
transform -1 0 90 0 1 7030
box -12 -8 32 272
use FILL  FILL_3__1683_
timestamp 1701859473
transform 1 0 70 0 1 6510
box -12 -8 32 272
use FILL  FILL_3__1684_
timestamp 1701859473
transform 1 0 950 0 -1 11190
box -12 -8 32 272
use FILL  FILL_3__1685_
timestamp 1701859473
transform -1 0 1210 0 -1 11190
box -12 -8 32 272
use FILL  FILL_3__1686_
timestamp 1701859473
transform -1 0 1010 0 1 10670
box -12 -8 32 272
use FILL  FILL_3__1687_
timestamp 1701859473
transform 1 0 1430 0 -1 11190
box -12 -8 32 272
use FILL  FILL_3__1688_
timestamp 1701859473
transform -1 0 1690 0 -1 11190
box -12 -8 32 272
use FILL  FILL_3__1689_
timestamp 1701859473
transform -1 0 1950 0 1 10150
box -12 -8 32 272
use FILL  FILL_3__1690_
timestamp 1701859473
transform 1 0 2110 0 1 9110
box -12 -8 32 272
use FILL  FILL_3__1691_
timestamp 1701859473
transform -1 0 2130 0 -1 9110
box -12 -8 32 272
use FILL  FILL_3__1692_
timestamp 1701859473
transform 1 0 70 0 1 790
box -12 -8 32 272
use FILL  FILL_3__1693_
timestamp 1701859473
transform 1 0 70 0 -1 1310
box -12 -8 32 272
use FILL  FILL_3__1694_
timestamp 1701859473
transform 1 0 490 0 -1 270
box -12 -8 32 272
use FILL  FILL_3__1695_
timestamp 1701859473
transform -1 0 710 0 -1 270
box -12 -8 32 272
use FILL  FILL_3__1696_
timestamp 1701859473
transform 1 0 1130 0 1 2870
box -12 -8 32 272
use FILL  FILL_3__1697_
timestamp 1701859473
transform -1 0 2790 0 -1 2870
box -12 -8 32 272
use FILL  FILL_3__1698_
timestamp 1701859473
transform -1 0 1890 0 1 3390
box -12 -8 32 272
use FILL  FILL_3__1699_
timestamp 1701859473
transform 1 0 3810 0 1 3390
box -12 -8 32 272
use FILL  FILL_3__1700_
timestamp 1701859473
transform -1 0 2610 0 -1 3910
box -12 -8 32 272
use FILL  FILL_3__1701_
timestamp 1701859473
transform -1 0 1150 0 1 270
box -12 -8 32 272
use FILL  FILL_3__1702_
timestamp 1701859473
transform 1 0 910 0 1 270
box -12 -8 32 272
use FILL  FILL_3__1703_
timestamp 1701859473
transform -1 0 1390 0 1 1830
box -12 -8 32 272
use FILL  FILL_3__1704_
timestamp 1701859473
transform -1 0 9150 0 1 2870
box -12 -8 32 272
use FILL  FILL_3__1705_
timestamp 1701859473
transform 1 0 9770 0 -1 790
box -12 -8 32 272
use FILL  FILL_3__1706_
timestamp 1701859473
transform -1 0 7990 0 -1 4950
box -12 -8 32 272
use FILL  FILL_3__1707_
timestamp 1701859473
transform 1 0 8430 0 -1 4950
box -12 -8 32 272
use FILL  FILL_3__1708_
timestamp 1701859473
transform 1 0 5050 0 -1 5990
box -12 -8 32 272
use FILL  FILL_3__1709_
timestamp 1701859473
transform -1 0 11150 0 1 5990
box -12 -8 32 272
use FILL  FILL_3__1710_
timestamp 1701859473
transform 1 0 5430 0 -1 5470
box -12 -8 32 272
use FILL  FILL_3__1711_
timestamp 1701859473
transform -1 0 5270 0 -1 5990
box -12 -8 32 272
use FILL  FILL_3__1712_
timestamp 1701859473
transform -1 0 5090 0 1 5470
box -12 -8 32 272
use FILL  FILL_3__1713_
timestamp 1701859473
transform 1 0 7950 0 1 4430
box -12 -8 32 272
use FILL  FILL_3__1714_
timestamp 1701859473
transform 1 0 7750 0 1 4950
box -12 -8 32 272
use FILL  FILL_3__1715_
timestamp 1701859473
transform -1 0 7990 0 1 4950
box -12 -8 32 272
use FILL  FILL_3__1716_
timestamp 1701859473
transform -1 0 8210 0 1 4430
box -12 -8 32 272
use FILL  FILL_3__1717_
timestamp 1701859473
transform -1 0 7990 0 1 1310
box -12 -8 32 272
use FILL  FILL_3__1718_
timestamp 1701859473
transform -1 0 5930 0 1 5990
box -12 -8 32 272
use FILL  FILL_3__1719_
timestamp 1701859473
transform -1 0 6790 0 -1 5990
box -12 -8 32 272
use FILL  FILL_3__1720_
timestamp 1701859473
transform -1 0 6770 0 1 5470
box -12 -8 32 272
use FILL  FILL_3__1721_
timestamp 1701859473
transform -1 0 7010 0 1 5470
box -12 -8 32 272
use FILL  FILL_3__1722_
timestamp 1701859473
transform -1 0 7710 0 1 4430
box -12 -8 32 272
use FILL  FILL_3__1723_
timestamp 1701859473
transform 1 0 7930 0 1 1830
box -12 -8 32 272
use FILL  FILL_3__1724_
timestamp 1701859473
transform -1 0 7970 0 -1 1310
box -12 -8 32 272
use FILL  FILL_3__1725_
timestamp 1701859473
transform 1 0 6570 0 1 5990
box -12 -8 32 272
use FILL  FILL_3__1726_
timestamp 1701859473
transform 1 0 6770 0 1 5990
box -12 -8 32 272
use FILL  FILL_3__1727_
timestamp 1701859473
transform -1 0 7010 0 1 5990
box -12 -8 32 272
use FILL  FILL_3__1728_
timestamp 1701859473
transform 1 0 7710 0 1 5990
box -12 -8 32 272
use FILL  FILL_3__1729_
timestamp 1701859473
transform -1 0 7650 0 -1 5990
box -12 -8 32 272
use FILL  FILL_3__1730_
timestamp 1701859473
transform -1 0 8130 0 1 3390
box -12 -8 32 272
use FILL  FILL_3__1731_
timestamp 1701859473
transform -1 0 7990 0 -1 270
box -12 -8 32 272
use FILL  FILL_3__1732_
timestamp 1701859473
transform -1 0 7950 0 1 5470
box -12 -8 32 272
use FILL  FILL_3__1733_
timestamp 1701859473
transform -1 0 8170 0 1 5470
box -12 -8 32 272
use FILL  FILL_3__1734_
timestamp 1701859473
transform 1 0 8130 0 -1 5470
box -12 -8 32 272
use FILL  FILL_3__1735_
timestamp 1701859473
transform 1 0 8590 0 -1 5470
box -12 -8 32 272
use FILL  FILL_3__1736_
timestamp 1701859473
transform 1 0 8430 0 1 4950
box -12 -8 32 272
use FILL  FILL_3__1737_
timestamp 1701859473
transform -1 0 8510 0 -1 3910
box -12 -8 32 272
use FILL  FILL_3__1738_
timestamp 1701859473
transform 1 0 8910 0 1 790
box -12 -8 32 272
use FILL  FILL_3__1739_
timestamp 1701859473
transform -1 0 9130 0 -1 790
box -12 -8 32 272
use FILL  FILL_3__1740_
timestamp 1701859473
transform 1 0 6490 0 1 270
box -12 -8 32 272
use FILL  FILL_3__1741_
timestamp 1701859473
transform 1 0 6390 0 1 790
box -12 -8 32 272
use FILL  FILL_3__1742_
timestamp 1701859473
transform -1 0 6330 0 -1 790
box -12 -8 32 272
use FILL  FILL_3__1743_
timestamp 1701859473
transform -1 0 2330 0 -1 3390
box -12 -8 32 272
use FILL  FILL_3__1744_
timestamp 1701859473
transform 1 0 310 0 -1 4950
box -12 -8 32 272
use FILL  FILL_3__1745_
timestamp 1701859473
transform 1 0 2130 0 -1 3910
box -12 -8 32 272
use FILL  FILL_3__1746_
timestamp 1701859473
transform -1 0 5150 0 -1 3390
box -12 -8 32 272
use FILL  FILL_3__1747_
timestamp 1701859473
transform -1 0 310 0 -1 270
box -12 -8 32 272
use FILL  FILL_3__1748_
timestamp 1701859473
transform -1 0 510 0 1 270
box -12 -8 32 272
use FILL  FILL_3__1749_
timestamp 1701859473
transform -1 0 950 0 1 1310
box -12 -8 32 272
use FILL  FILL_3__1750_
timestamp 1701859473
transform -1 0 1170 0 1 1310
box -12 -8 32 272
use FILL  FILL_3__1751_
timestamp 1701859473
transform -1 0 4530 0 -1 2870
box -12 -8 32 272
use FILL  FILL_3__1752_
timestamp 1701859473
transform 1 0 4730 0 -1 2870
box -12 -8 32 272
use FILL  FILL_3__1753_
timestamp 1701859473
transform -1 0 4350 0 1 790
box -12 -8 32 272
use FILL  FILL_3__1754_
timestamp 1701859473
transform 1 0 290 0 -1 790
box -12 -8 32 272
use FILL  FILL_3__1755_
timestamp 1701859473
transform -1 0 510 0 -1 790
box -12 -8 32 272
use FILL  FILL_3__1756_
timestamp 1701859473
transform -1 0 90 0 -1 270
box -12 -8 32 272
use FILL  FILL_3__1757_
timestamp 1701859473
transform 1 0 690 0 -1 790
box -12 -8 32 272
use FILL  FILL_3__1758_
timestamp 1701859473
transform 1 0 70 0 1 2350
box -12 -8 32 272
use FILL  FILL_3__1759_
timestamp 1701859473
transform -1 0 2570 0 -1 2870
box -12 -8 32 272
use FILL  FILL_3__1760_
timestamp 1701859473
transform 1 0 2950 0 -1 2870
box -12 -8 32 272
use FILL  FILL_3__1761_
timestamp 1701859473
transform -1 0 3270 0 -1 3390
box -12 -8 32 272
use FILL  FILL_3__1762_
timestamp 1701859473
transform -1 0 90 0 1 270
box -12 -8 32 272
use FILL  FILL_3__1763_
timestamp 1701859473
transform 1 0 70 0 -1 790
box -12 -8 32 272
use FILL  FILL_3__1764_
timestamp 1701859473
transform 1 0 510 0 1 1310
box -12 -8 32 272
use FILL  FILL_3__1765_
timestamp 1701859473
transform 1 0 1370 0 1 1310
box -12 -8 32 272
use FILL  FILL_3__1766_
timestamp 1701859473
transform -1 0 3170 0 -1 1830
box -12 -8 32 272
use FILL  FILL_3__1767_
timestamp 1701859473
transform 1 0 1470 0 -1 4430
box -12 -8 32 272
use FILL  FILL_3__1768_
timestamp 1701859473
transform 1 0 290 0 -1 1310
box -12 -8 32 272
use FILL  FILL_3__1769_
timestamp 1701859473
transform -1 0 510 0 1 1830
box -12 -8 32 272
use FILL  FILL_3__1770_
timestamp 1701859473
transform 1 0 2110 0 -1 3390
box -12 -8 32 272
use FILL  FILL_3__1771_
timestamp 1701859473
transform -1 0 2370 0 -1 3910
box -12 -8 32 272
use FILL  FILL_3__1772_
timestamp 1701859473
transform -1 0 3030 0 -1 3910
box -12 -8 32 272
use FILL  FILL_3__1773_
timestamp 1701859473
transform 1 0 3930 0 1 2870
box -12 -8 32 272
use FILL  FILL_3__1774_
timestamp 1701859473
transform -1 0 5310 0 -1 2350
box -12 -8 32 272
use FILL  FILL_3__1775_
timestamp 1701859473
transform 1 0 270 0 1 790
box -12 -8 32 272
use FILL  FILL_3__1776_
timestamp 1701859473
transform -1 0 310 0 1 1310
box -12 -8 32 272
use FILL  FILL_3__1777_
timestamp 1701859473
transform 1 0 730 0 -1 1830
box -12 -8 32 272
use FILL  FILL_3__1778_
timestamp 1701859473
transform -1 0 4450 0 1 5470
box -12 -8 32 272
use FILL  FILL_3__1779_
timestamp 1701859473
transform -1 0 6090 0 -1 5470
box -12 -8 32 272
use FILL  FILL_3__1780_
timestamp 1701859473
transform 1 0 4810 0 1 2870
box -12 -8 32 272
use FILL  FILL_3__1781_
timestamp 1701859473
transform 1 0 4390 0 1 2870
box -12 -8 32 272
use FILL  FILL_3__1782_
timestamp 1701859473
transform -1 0 90 0 1 1310
box -12 -8 32 272
use FILL  FILL_3__1783_
timestamp 1701859473
transform -1 0 1370 0 1 2870
box -12 -8 32 272
use FILL  FILL_3__1784_
timestamp 1701859473
transform -1 0 5070 0 1 2870
box -12 -8 32 272
use FILL  FILL_3__1785_
timestamp 1701859473
transform 1 0 4990 0 -1 2870
box -12 -8 32 272
use FILL  FILL_3__1786_
timestamp 1701859473
transform -1 0 5070 0 -1 2350
box -12 -8 32 272
use FILL  FILL_3__1787_
timestamp 1701859473
transform 1 0 5050 0 1 2350
box -12 -8 32 272
use FILL  FILL_3__1788_
timestamp 1701859473
transform -1 0 4850 0 -1 2350
box -12 -8 32 272
use FILL  FILL_3__1789_
timestamp 1701859473
transform 1 0 70 0 1 1830
box -12 -8 32 272
use FILL  FILL_3__1790_
timestamp 1701859473
transform -1 0 310 0 -1 2350
box -12 -8 32 272
use FILL  FILL_3__1791_
timestamp 1701859473
transform -1 0 2110 0 -1 2350
box -12 -8 32 272
use FILL  FILL_3__1792_
timestamp 1701859473
transform -1 0 3490 0 -1 2350
box -12 -8 32 272
use FILL  FILL_3__1793_
timestamp 1701859473
transform -1 0 4590 0 1 1830
box -12 -8 32 272
use FILL  FILL_3__1794_
timestamp 1701859473
transform 1 0 910 0 1 1830
box -12 -8 32 272
use FILL  FILL_3__1795_
timestamp 1701859473
transform -1 0 2170 0 1 2350
box -12 -8 32 272
use FILL  FILL_3__1796_
timestamp 1701859473
transform -1 0 1790 0 -1 1830
box -12 -8 32 272
use FILL  FILL_3__1797_
timestamp 1701859473
transform 1 0 2010 0 -1 1830
box -12 -8 32 272
use FILL  FILL_3__1798_
timestamp 1701859473
transform 1 0 930 0 -1 1310
box -12 -8 32 272
use FILL  FILL_3__1799_
timestamp 1701859473
transform 1 0 3750 0 1 3910
box -12 -8 32 272
use FILL  FILL_3__1800_
timestamp 1701859473
transform 1 0 3430 0 1 1830
box -12 -8 32 272
use FILL  FILL_3__1801_
timestamp 1701859473
transform -1 0 1170 0 1 1830
box -12 -8 32 272
use FILL  FILL_3__1802_
timestamp 1701859473
transform -1 0 3710 0 1 2350
box -12 -8 32 272
use FILL  FILL_3__1803_
timestamp 1701859473
transform -1 0 3930 0 1 2350
box -12 -8 32 272
use FILL  FILL_3__1804_
timestamp 1701859473
transform -1 0 4170 0 1 2350
box -12 -8 32 272
use FILL  FILL_3__1805_
timestamp 1701859473
transform 1 0 5470 0 1 2350
box -12 -8 32 272
use FILL  FILL_3__1806_
timestamp 1701859473
transform -1 0 4870 0 1 2350
box -12 -8 32 272
use FILL  FILL_3__1807_
timestamp 1701859473
transform -1 0 5270 0 1 2350
box -12 -8 32 272
use FILL  FILL_3__1808_
timestamp 1701859473
transform 1 0 4790 0 1 1830
box -12 -8 32 272
use FILL  FILL_3__1809_
timestamp 1701859473
transform -1 0 7150 0 -1 270
box -12 -8 32 272
use FILL  FILL_3__1810_
timestamp 1701859473
transform -1 0 7130 0 1 1310
box -12 -8 32 272
use FILL  FILL_3__1811_
timestamp 1701859473
transform 1 0 7470 0 -1 1830
box -12 -8 32 272
use FILL  FILL_3__1812_
timestamp 1701859473
transform -1 0 7550 0 -1 1310
box -12 -8 32 272
use FILL  FILL_3__1813_
timestamp 1701859473
transform 1 0 9130 0 1 790
box -12 -8 32 272
use FILL  FILL_3__1814_
timestamp 1701859473
transform -1 0 8170 0 -1 1830
box -12 -8 32 272
use FILL  FILL_3__1815_
timestamp 1701859473
transform 1 0 8370 0 1 2350
box -12 -8 32 272
use FILL  FILL_3__1816_
timestamp 1701859473
transform -1 0 9650 0 -1 2350
box -12 -8 32 272
use FILL  FILL_3__1817_
timestamp 1701859473
transform -1 0 9370 0 1 1310
box -12 -8 32 272
use FILL  FILL_3__1818_
timestamp 1701859473
transform -1 0 9570 0 1 270
box -12 -8 32 272
use FILL  FILL_3__1819_
timestamp 1701859473
transform -1 0 8390 0 -1 1830
box -12 -8 32 272
use FILL  FILL_3__1820_
timestamp 1701859473
transform -1 0 8470 0 1 1310
box -12 -8 32 272
use FILL  FILL_3__1821_
timestamp 1701859473
transform -1 0 4910 0 1 1310
box -12 -8 32 272
use FILL  FILL_3__1822_
timestamp 1701859473
transform -1 0 4710 0 -1 790
box -12 -8 32 272
use FILL  FILL_3__1823_
timestamp 1701859473
transform -1 0 4250 0 -1 790
box -12 -8 32 272
use FILL  FILL_3__1824_
timestamp 1701859473
transform 1 0 4630 0 1 2350
box -12 -8 32 272
use FILL  FILL_3__1825_
timestamp 1701859473
transform 1 0 5690 0 1 1830
box -12 -8 32 272
use FILL  FILL_3__1826_
timestamp 1701859473
transform 1 0 8190 0 -1 270
box -12 -8 32 272
use FILL  FILL_3__1827_
timestamp 1701859473
transform 1 0 9330 0 -1 790
box -12 -8 32 272
use FILL  FILL_3__1828_
timestamp 1701859473
transform 1 0 8490 0 1 270
box -12 -8 32 272
use FILL  FILL_3__1829_
timestamp 1701859473
transform 1 0 5790 0 1 270
box -12 -8 32 272
use FILL  FILL_3__1830_
timestamp 1701859473
transform 1 0 3230 0 1 4430
box -12 -8 32 272
use FILL  FILL_3__1831_
timestamp 1701859473
transform -1 0 8010 0 -1 790
box -12 -8 32 272
use FILL  FILL_3__1832_
timestamp 1701859473
transform 1 0 6510 0 -1 790
box -12 -8 32 272
use FILL  FILL_3__1833_
timestamp 1701859473
transform -1 0 710 0 1 270
box -12 -8 32 272
use FILL  FILL_3__1834_
timestamp 1701859473
transform 1 0 1150 0 -1 1310
box -12 -8 32 272
use FILL  FILL_3__1835_
timestamp 1701859473
transform -1 0 2530 0 -1 1310
box -12 -8 32 272
use FILL  FILL_3__1836_
timestamp 1701859473
transform 1 0 1090 0 1 790
box -12 -8 32 272
use FILL  FILL_3__1837_
timestamp 1701859473
transform -1 0 2490 0 1 790
box -12 -8 32 272
use FILL  FILL_3__1838_
timestamp 1701859473
transform 1 0 2230 0 1 790
box -12 -8 32 272
use FILL  FILL_3__1839_
timestamp 1701859473
transform -1 0 290 0 1 270
box -12 -8 32 272
use FILL  FILL_3__1840_
timestamp 1701859473
transform -1 0 930 0 1 2870
box -12 -8 32 272
use FILL  FILL_3__1841_
timestamp 1701859473
transform 1 0 3710 0 1 2870
box -12 -8 32 272
use FILL  FILL_3__1842_
timestamp 1701859473
transform -1 0 2970 0 -1 1830
box -12 -8 32 272
use FILL  FILL_3__1843_
timestamp 1701859473
transform -1 0 3930 0 -1 2350
box -12 -8 32 272
use FILL  FILL_3__1844_
timestamp 1701859473
transform 1 0 3830 0 -1 2870
box -12 -8 32 272
use FILL  FILL_3__1845_
timestamp 1701859473
transform -1 0 1770 0 -1 4950
box -12 -8 32 272
use FILL  FILL_3__1846_
timestamp 1701859473
transform 1 0 4130 0 1 4430
box -12 -8 32 272
use FILL  FILL_3__1847_
timestamp 1701859473
transform 1 0 3450 0 1 4430
box -12 -8 32 272
use FILL  FILL_3__1848_
timestamp 1701859473
transform 1 0 3890 0 1 4430
box -12 -8 32 272
use FILL  FILL_3__1849_
timestamp 1701859473
transform -1 0 4090 0 -1 2870
box -12 -8 32 272
use FILL  FILL_3__1850_
timestamp 1701859473
transform -1 0 910 0 1 790
box -12 -8 32 272
use FILL  FILL_3__1851_
timestamp 1701859473
transform 1 0 1570 0 -1 1830
box -12 -8 32 272
use FILL  FILL_3__1852_
timestamp 1701859473
transform -1 0 2390 0 1 2350
box -12 -8 32 272
use FILL  FILL_3__1853_
timestamp 1701859473
transform 1 0 70 0 -1 2350
box -12 -8 32 272
use FILL  FILL_3__1854_
timestamp 1701859473
transform 1 0 2310 0 -1 2350
box -12 -8 32 272
use FILL  FILL_3__1855_
timestamp 1701859473
transform -1 0 2570 0 -1 2350
box -12 -8 32 272
use FILL  FILL_3__1856_
timestamp 1701859473
transform 1 0 1470 0 -1 790
box -12 -8 32 272
use FILL  FILL_3__1857_
timestamp 1701859473
transform -1 0 2670 0 -1 790
box -12 -8 32 272
use FILL  FILL_3__1858_
timestamp 1701859473
transform 1 0 2410 0 -1 790
box -12 -8 32 272
use FILL  FILL_3__1859_
timestamp 1701859473
transform 1 0 2190 0 -1 790
box -12 -8 32 272
use FILL  FILL_3__1860_
timestamp 1701859473
transform -1 0 1730 0 -1 790
box -12 -8 32 272
use FILL  FILL_3__1861_
timestamp 1701859473
transform -1 0 1970 0 -1 790
box -12 -8 32 272
use FILL  FILL_3__1862_
timestamp 1701859473
transform -1 0 2050 0 1 270
box -12 -8 32 272
use FILL  FILL_3__1863_
timestamp 1701859473
transform 1 0 2270 0 1 270
box -12 -8 32 272
use FILL  FILL_3__1864_
timestamp 1701859473
transform 1 0 3510 0 1 270
box -12 -8 32 272
use FILL  FILL_3__1865_
timestamp 1701859473
transform 1 0 7310 0 -1 1310
box -12 -8 32 272
use FILL  FILL_3__1866_
timestamp 1701859473
transform 1 0 3670 0 -1 1310
box -12 -8 32 272
use FILL  FILL_3__1867_
timestamp 1701859473
transform 1 0 1130 0 -1 1830
box -12 -8 32 272
use FILL  FILL_3__1868_
timestamp 1701859473
transform 1 0 1570 0 1 1310
box -12 -8 32 272
use FILL  FILL_3__1869_
timestamp 1701859473
transform 1 0 1990 0 1 1310
box -12 -8 32 272
use FILL  FILL_3__1870_
timestamp 1701859473
transform -1 0 1610 0 -1 1310
box -12 -8 32 272
use FILL  FILL_3__1871_
timestamp 1701859473
transform -1 0 2730 0 -1 1310
box -12 -8 32 272
use FILL  FILL_3__1872_
timestamp 1701859473
transform -1 0 510 0 1 790
box -12 -8 32 272
use FILL  FILL_3__1873_
timestamp 1701859473
transform 1 0 690 0 1 790
box -12 -8 32 272
use FILL  FILL_3__1874_
timestamp 1701859473
transform -1 0 1330 0 1 790
box -12 -8 32 272
use FILL  FILL_3__1875_
timestamp 1701859473
transform 1 0 910 0 -1 790
box -12 -8 32 272
use FILL  FILL_3__1876_
timestamp 1701859473
transform 1 0 1230 0 -1 790
box -12 -8 32 272
use FILL  FILL_3__1877_
timestamp 1701859473
transform 1 0 2170 0 1 4950
box -12 -8 32 272
use FILL  FILL_3__1878_
timestamp 1701859473
transform 1 0 510 0 -1 1310
box -12 -8 32 272
use FILL  FILL_3__1879_
timestamp 1701859473
transform 1 0 730 0 1 1310
box -12 -8 32 272
use FILL  FILL_3__1880_
timestamp 1701859473
transform -1 0 1990 0 -1 4950
box -12 -8 32 272
use FILL  FILL_3__1881_
timestamp 1701859473
transform -1 0 2230 0 -1 4950
box -12 -8 32 272
use FILL  FILL_3__1882_
timestamp 1701859473
transform 1 0 1550 0 -1 3390
box -12 -8 32 272
use FILL  FILL_3__1883_
timestamp 1701859473
transform 1 0 1030 0 -1 3390
box -12 -8 32 272
use FILL  FILL_3__1884_
timestamp 1701859473
transform -1 0 4050 0 1 3390
box -12 -8 32 272
use FILL  FILL_3__1885_
timestamp 1701859473
transform -1 0 3770 0 -1 3390
box -12 -8 32 272
use FILL  FILL_3__1886_
timestamp 1701859473
transform 1 0 3510 0 -1 3390
box -12 -8 32 272
use FILL  FILL_3__1887_
timestamp 1701859473
transform -1 0 3490 0 1 2870
box -12 -8 32 272
use FILL  FILL_3__1888_
timestamp 1701859473
transform -1 0 2530 0 1 270
box -12 -8 32 272
use FILL  FILL_3__1889_
timestamp 1701859473
transform 1 0 1670 0 -1 2870
box -12 -8 32 272
use FILL  FILL_3__1890_
timestamp 1701859473
transform -1 0 310 0 -1 1830
box -12 -8 32 272
use FILL  FILL_3__1891_
timestamp 1701859473
transform 1 0 70 0 -1 1830
box -12 -8 32 272
use FILL  FILL_3__1892_
timestamp 1701859473
transform 1 0 4910 0 -1 3390
box -12 -8 32 272
use FILL  FILL_3__1893_
timestamp 1701859473
transform 1 0 3910 0 1 1830
box -12 -8 32 272
use FILL  FILL_3__1894_
timestamp 1701859473
transform 1 0 4110 0 1 1830
box -12 -8 32 272
use FILL  FILL_3__1895_
timestamp 1701859473
transform -1 0 1850 0 1 1830
box -12 -8 32 272
use FILL  FILL_3__1896_
timestamp 1701859473
transform 1 0 1870 0 -1 2350
box -12 -8 32 272
use FILL  FILL_3__1897_
timestamp 1701859473
transform 1 0 3490 0 1 2350
box -12 -8 32 272
use FILL  FILL_3__1898_
timestamp 1701859473
transform 1 0 3270 0 1 2350
box -12 -8 32 272
use FILL  FILL_3__1899_
timestamp 1701859473
transform -1 0 3250 0 -1 2350
box -12 -8 32 272
use FILL  FILL_3__1900_
timestamp 1701859473
transform -1 0 4090 0 -1 1830
box -12 -8 32 272
use FILL  FILL_3__1901_
timestamp 1701859473
transform -1 0 730 0 1 1830
box -12 -8 32 272
use FILL  FILL_3__1902_
timestamp 1701859473
transform 1 0 5030 0 1 1830
box -12 -8 32 272
use FILL  FILL_3__1903_
timestamp 1701859473
transform 1 0 3350 0 1 1310
box -12 -8 32 272
use FILL  FILL_3__1904_
timestamp 1701859473
transform -1 0 3450 0 -1 1310
box -12 -8 32 272
use FILL  FILL_3__1905_
timestamp 1701859473
transform 1 0 2990 0 1 270
box -12 -8 32 272
use FILL  FILL_3__1906_
timestamp 1701859473
transform 1 0 270 0 1 2350
box -12 -8 32 272
use FILL  FILL_3__1907_
timestamp 1701859473
transform -1 0 3030 0 -1 2350
box -12 -8 32 272
use FILL  FILL_3__1908_
timestamp 1701859473
transform 1 0 6450 0 -1 2350
box -12 -8 32 272
use FILL  FILL_3__1909_
timestamp 1701859473
transform -1 0 6050 0 -1 2350
box -12 -8 32 272
use FILL  FILL_3__1910_
timestamp 1701859473
transform -1 0 5550 0 -1 2350
box -12 -8 32 272
use FILL  FILL_3__1911_
timestamp 1701859473
transform -1 0 710 0 1 2870
box -12 -8 32 272
use FILL  FILL_3__1912_
timestamp 1701859473
transform -1 0 3310 0 1 3910
box -12 -8 32 272
use FILL  FILL_3__1913_
timestamp 1701859473
transform -1 0 1030 0 -1 2870
box -12 -8 32 272
use FILL  FILL_3__1914_
timestamp 1701859473
transform -1 0 1470 0 1 3390
box -12 -8 32 272
use FILL  FILL_3__1915_
timestamp 1701859473
transform 1 0 2550 0 1 3390
box -12 -8 32 272
use FILL  FILL_3__1916_
timestamp 1701859473
transform -1 0 3410 0 1 3390
box -12 -8 32 272
use FILL  FILL_3__1917_
timestamp 1701859473
transform -1 0 4690 0 -1 3390
box -12 -8 32 272
use FILL  FILL_3__1918_
timestamp 1701859473
transform 1 0 1730 0 1 4950
box -12 -8 32 272
use FILL  FILL_3__1919_
timestamp 1701859473
transform -1 0 1250 0 -1 2870
box -12 -8 32 272
use FILL  FILL_3__1920_
timestamp 1701859473
transform -1 0 5030 0 1 4430
box -12 -8 32 272
use FILL  FILL_3__1921_
timestamp 1701859473
transform 1 0 4790 0 1 4430
box -12 -8 32 272
use FILL  FILL_3__1922_
timestamp 1701859473
transform -1 0 4590 0 1 4430
box -12 -8 32 272
use FILL  FILL_3__1923_
timestamp 1701859473
transform 1 0 4450 0 -1 3390
box -12 -8 32 272
use FILL  FILL_3__1924_
timestamp 1701859473
transform 1 0 1950 0 1 4950
box -12 -8 32 272
use FILL  FILL_3__1925_
timestamp 1701859473
transform 1 0 6090 0 -1 4430
box -12 -8 32 272
use FILL  FILL_3__1926_
timestamp 1701859473
transform 1 0 710 0 -1 1310
box -12 -8 32 272
use FILL  FILL_3__1927_
timestamp 1701859473
transform 1 0 2950 0 -1 1310
box -12 -8 32 272
use FILL  FILL_3__1928_
timestamp 1701859473
transform -1 0 3210 0 -1 1310
box -12 -8 32 272
use FILL  FILL_3__1929_
timestamp 1701859473
transform 1 0 3390 0 1 790
box -12 -8 32 272
use FILL  FILL_3__1930_
timestamp 1701859473
transform 1 0 3210 0 1 270
box -12 -8 32 272
use FILL  FILL_3__1931_
timestamp 1701859473
transform 1 0 3810 0 1 270
box -12 -8 32 272
use FILL  FILL_3__1932_
timestamp 1701859473
transform -1 0 4050 0 1 270
box -12 -8 32 272
use FILL  FILL_3__1933_
timestamp 1701859473
transform -1 0 1850 0 1 270
box -12 -8 32 272
use FILL  FILL_3__1934_
timestamp 1701859473
transform -1 0 5470 0 1 790
box -12 -8 32 272
use FILL  FILL_3__1935_
timestamp 1701859473
transform 1 0 5590 0 -1 270
box -12 -8 32 272
use FILL  FILL_3__1936_
timestamp 1701859473
transform -1 0 8350 0 1 3390
box -12 -8 32 272
use FILL  FILL_3__1937_
timestamp 1701859473
transform -1 0 7570 0 -1 270
box -12 -8 32 272
use FILL  FILL_3__1938_
timestamp 1701859473
transform -1 0 7770 0 -1 270
box -12 -8 32 272
use FILL  FILL_3__1939_
timestamp 1701859473
transform -1 0 6690 0 -1 270
box -12 -8 32 272
use FILL  FILL_3__1940_
timestamp 1701859473
transform -1 0 5810 0 -1 270
box -12 -8 32 272
use FILL  FILL_3__1941_
timestamp 1701859473
transform 1 0 5830 0 -1 790
box -12 -8 32 272
use FILL  FILL_3__1942_
timestamp 1701859473
transform 1 0 4810 0 -1 1310
box -12 -8 32 272
use FILL  FILL_3__1943_
timestamp 1701859473
transform 1 0 8070 0 1 270
box -12 -8 32 272
use FILL  FILL_3__1944_
timestamp 1701859473
transform -1 0 8310 0 1 270
box -12 -8 32 272
use FILL  FILL_3__1945_
timestamp 1701859473
transform 1 0 7850 0 1 270
box -12 -8 32 272
use FILL  FILL_3__1946_
timestamp 1701859473
transform -1 0 6050 0 1 270
box -12 -8 32 272
use FILL  FILL_3__1947_
timestamp 1701859473
transform -1 0 6070 0 -1 790
box -12 -8 32 272
use FILL  FILL_3__1948_
timestamp 1701859473
transform 1 0 5350 0 -1 790
box -12 -8 32 272
use FILL  FILL_3__1949_
timestamp 1701859473
transform 1 0 4590 0 -1 1310
box -12 -8 32 272
use FILL  FILL_3__1950_
timestamp 1701859473
transform -1 0 8230 0 -1 790
box -12 -8 32 272
use FILL  FILL_3__1951_
timestamp 1701859473
transform 1 0 510 0 -1 2350
box -12 -8 32 272
use FILL  FILL_3__1952_
timestamp 1701859473
transform -1 0 5690 0 1 2350
box -12 -8 32 272
use FILL  FILL_3__1953_
timestamp 1701859473
transform 1 0 5790 0 -1 2350
box -12 -8 32 272
use FILL  FILL_3__1954_
timestamp 1701859473
transform 1 0 8170 0 -1 1310
box -12 -8 32 272
use FILL  FILL_3__1955_
timestamp 1701859473
transform -1 0 8710 0 1 1310
box -12 -8 32 272
use FILL  FILL_3__1956_
timestamp 1701859473
transform -1 0 6250 0 -1 1310
box -12 -8 32 272
use FILL  FILL_3__1957_
timestamp 1701859473
transform -1 0 6010 0 -1 1310
box -12 -8 32 272
use FILL  FILL_3__1958_
timestamp 1701859473
transform 1 0 5270 0 -1 1310
box -12 -8 32 272
use FILL  FILL_3__1959_
timestamp 1701859473
transform 1 0 5710 0 -1 2870
box -12 -8 32 272
use FILL  FILL_3__1960_
timestamp 1701859473
transform -1 0 6150 0 -1 2870
box -12 -8 32 272
use FILL  FILL_3__1961_
timestamp 1701859473
transform -1 0 4410 0 1 2350
box -12 -8 32 272
use FILL  FILL_3__1962_
timestamp 1701859473
transform 1 0 5870 0 1 2350
box -12 -8 32 272
use FILL  FILL_3__1963_
timestamp 1701859473
transform 1 0 5330 0 1 1310
box -12 -8 32 272
use FILL  FILL_3__1964_
timestamp 1701859473
transform 1 0 9150 0 1 1310
box -12 -8 32 272
use FILL  FILL_3__1965_
timestamp 1701859473
transform 1 0 7550 0 1 790
box -12 -8 32 272
use FILL  FILL_3__1966_
timestamp 1701859473
transform -1 0 7670 0 1 270
box -12 -8 32 272
use FILL  FILL_3__1967_
timestamp 1701859473
transform -1 0 6730 0 1 270
box -12 -8 32 272
use FILL  FILL_3__1968_
timestamp 1701859473
transform 1 0 5510 0 -1 1310
box -12 -8 32 272
use FILL  FILL_3__1969_
timestamp 1701859473
transform 1 0 5710 0 1 2870
box -12 -8 32 272
use FILL  FILL_3__1970_
timestamp 1701859473
transform 1 0 5350 0 -1 3390
box -12 -8 32 272
use FILL  FILL_3__1971_
timestamp 1701859473
transform 1 0 5790 0 1 3910
box -12 -8 32 272
use FILL  FILL_3__1972_
timestamp 1701859473
transform 1 0 5730 0 1 4950
box -12 -8 32 272
use FILL  FILL_3__1973_
timestamp 1701859473
transform -1 0 6070 0 -1 3910
box -12 -8 32 272
use FILL  FILL_3__1974_
timestamp 1701859473
transform 1 0 6250 0 -1 3910
box -12 -8 32 272
use FILL  FILL_3__1975_
timestamp 1701859473
transform -1 0 6050 0 1 3910
box -12 -8 32 272
use FILL  FILL_3__1976_
timestamp 1701859473
transform -1 0 6510 0 -1 3910
box -12 -8 32 272
use FILL  FILL_3__1977_
timestamp 1701859473
transform 1 0 6830 0 1 2870
box -12 -8 32 272
use FILL  FILL_3__1978_
timestamp 1701859473
transform -1 0 6370 0 -1 2870
box -12 -8 32 272
use FILL  FILL_3__1979_
timestamp 1701859473
transform 1 0 6410 0 1 2870
box -12 -8 32 272
use FILL  FILL_3__1980_
timestamp 1701859473
transform 1 0 6610 0 1 2870
box -12 -8 32 272
use FILL  FILL_3__1981_
timestamp 1701859473
transform 1 0 6190 0 1 2870
box -12 -8 32 272
use FILL  FILL_3__1982_
timestamp 1701859473
transform -1 0 5650 0 -1 1830
box -12 -8 32 272
use FILL  FILL_3__1983_
timestamp 1701859473
transform -1 0 4750 0 -1 270
box -12 -8 32 272
use FILL  FILL_3__1984_
timestamp 1701859473
transform -1 0 6450 0 -1 1310
box -12 -8 32 272
use FILL  FILL_3__1985_
timestamp 1701859473
transform 1 0 5010 0 -1 1310
box -12 -8 32 272
use FILL  FILL_3__1986_
timestamp 1701859473
transform 1 0 8210 0 1 790
box -12 -8 32 272
use FILL  FILL_3__1987_
timestamp 1701859473
transform 1 0 6890 0 1 1310
box -12 -8 32 272
use FILL  FILL_3__1988_
timestamp 1701859473
transform -1 0 7350 0 1 1310
box -12 -8 32 272
use FILL  FILL_3__1989_
timestamp 1701859473
transform 1 0 2710 0 -1 5470
box -12 -8 32 272
use FILL  FILL_3__1990_
timestamp 1701859473
transform 1 0 2030 0 1 1830
box -12 -8 32 272
use FILL  FILL_3__1991_
timestamp 1701859473
transform -1 0 2750 0 1 1830
box -12 -8 32 272
use FILL  FILL_3__1992_
timestamp 1701859473
transform -1 0 4150 0 -1 2350
box -12 -8 32 272
use FILL  FILL_3__1993_
timestamp 1701859473
transform -1 0 4390 0 -1 2350
box -12 -8 32 272
use FILL  FILL_3__1994_
timestamp 1701859473
transform 1 0 2490 0 1 1830
box -12 -8 32 272
use FILL  FILL_3__1995_
timestamp 1701859473
transform 1 0 2970 0 1 1830
box -12 -8 32 272
use FILL  FILL_3__1996_
timestamp 1701859473
transform -1 0 6650 0 1 790
box -12 -8 32 272
use FILL  FILL_3__1997_
timestamp 1701859473
transform -1 0 4990 0 1 790
box -12 -8 32 272
use FILL  FILL_3__1998_
timestamp 1701859473
transform 1 0 4250 0 1 270
box -12 -8 32 272
use FILL  FILL_3__1999_
timestamp 1701859473
transform -1 0 3850 0 -1 270
box -12 -8 32 272
use FILL  FILL_3__2000_
timestamp 1701859473
transform -1 0 4530 0 -1 270
box -12 -8 32 272
use FILL  FILL_3__2001_
timestamp 1701859473
transform -1 0 5910 0 -1 2870
box -12 -8 32 272
use FILL  FILL_3__2002_
timestamp 1701859473
transform -1 0 1850 0 1 2870
box -12 -8 32 272
use FILL  FILL_3__2003_
timestamp 1701859473
transform 1 0 1350 0 -1 3390
box -12 -8 32 272
use FILL  FILL_3__2004_
timestamp 1701859473
transform 1 0 2770 0 -1 3390
box -12 -8 32 272
use FILL  FILL_3__2005_
timestamp 1701859473
transform -1 0 3050 0 1 2870
box -12 -8 32 272
use FILL  FILL_3__2006_
timestamp 1701859473
transform 1 0 2790 0 1 2870
box -12 -8 32 272
use FILL  FILL_3__2007_
timestamp 1701859473
transform 1 0 6810 0 -1 2870
box -12 -8 32 272
use FILL  FILL_3__2008_
timestamp 1701859473
transform 1 0 490 0 -1 1830
box -12 -8 32 272
use FILL  FILL_3__2009_
timestamp 1701859473
transform -1 0 4010 0 -1 3390
box -12 -8 32 272
use FILL  FILL_3__2010_
timestamp 1701859473
transform -1 0 4310 0 -1 2870
box -12 -8 32 272
use FILL  FILL_3__2011_
timestamp 1701859473
transform -1 0 2050 0 1 790
box -12 -8 32 272
use FILL  FILL_3__2012_
timestamp 1701859473
transform 1 0 1550 0 1 790
box -12 -8 32 272
use FILL  FILL_3__2013_
timestamp 1701859473
transform -1 0 1810 0 1 790
box -12 -8 32 272
use FILL  FILL_3__2014_
timestamp 1701859473
transform 1 0 4470 0 1 1310
box -12 -8 32 272
use FILL  FILL_3__2015_
timestamp 1701859473
transform 1 0 3190 0 1 1830
box -12 -8 32 272
use FILL  FILL_3__2016_
timestamp 1701859473
transform -1 0 3690 0 1 1830
box -12 -8 32 272
use FILL  FILL_3__2017_
timestamp 1701859473
transform -1 0 5210 0 -1 1830
box -12 -8 32 272
use FILL  FILL_3__2018_
timestamp 1701859473
transform 1 0 4970 0 -1 1830
box -12 -8 32 272
use FILL  FILL_3__2019_
timestamp 1701859473
transform -1 0 5490 0 -1 2870
box -12 -8 32 272
use FILL  FILL_3__2020_
timestamp 1701859473
transform -1 0 5250 0 -1 2870
box -12 -8 32 272
use FILL  FILL_3__2021_
timestamp 1701859473
transform -1 0 6890 0 -1 1310
box -12 -8 32 272
use FILL  FILL_3__2022_
timestamp 1701859473
transform -1 0 7130 0 1 790
box -12 -8 32 272
use FILL  FILL_3__2023_
timestamp 1701859473
transform 1 0 8170 0 1 1830
box -12 -8 32 272
use FILL  FILL_3__2024_
timestamp 1701859473
transform -1 0 8390 0 1 1830
box -12 -8 32 272
use FILL  FILL_3__2025_
timestamp 1701859473
transform 1 0 9550 0 -1 790
box -12 -8 32 272
use FILL  FILL_3__2026_
timestamp 1701859473
transform -1 0 8690 0 1 790
box -12 -8 32 272
use FILL  FILL_3__2027_
timestamp 1701859473
transform -1 0 6890 0 1 790
box -12 -8 32 272
use FILL  FILL_3__2028_
timestamp 1701859473
transform 1 0 6990 0 -1 790
box -12 -8 32 272
use FILL  FILL_3__2029_
timestamp 1701859473
transform 1 0 7430 0 1 270
box -12 -8 32 272
use FILL  FILL_3__2030_
timestamp 1701859473
transform -1 0 7110 0 -1 1310
box -12 -8 32 272
use FILL  FILL_3__2031_
timestamp 1701859473
transform 1 0 7430 0 -1 790
box -12 -8 32 272
use FILL  FILL_3__2032_
timestamp 1701859473
transform -1 0 8730 0 1 270
box -12 -8 32 272
use FILL  FILL_3__2033_
timestamp 1701859473
transform 1 0 8210 0 1 1310
box -12 -8 32 272
use FILL  FILL_3__2034_
timestamp 1701859473
transform -1 0 8890 0 -1 1310
box -12 -8 32 272
use FILL  FILL_3__2035_
timestamp 1701859473
transform -1 0 8470 0 1 790
box -12 -8 32 272
use FILL  FILL_3__2036_
timestamp 1701859473
transform -1 0 8630 0 -1 1830
box -12 -8 32 272
use FILL  FILL_3__2037_
timestamp 1701859473
transform -1 0 8690 0 -1 790
box -12 -8 32 272
use FILL  FILL_3__2038_
timestamp 1701859473
transform 1 0 7990 0 1 790
box -12 -8 32 272
use FILL  FILL_3__2039_
timestamp 1701859473
transform 1 0 7770 0 1 790
box -12 -8 32 272
use FILL  FILL_3__2040_
timestamp 1701859473
transform -1 0 7690 0 -1 790
box -12 -8 32 272
use FILL  FILL_3__2041_
timestamp 1701859473
transform -1 0 6910 0 -1 270
box -12 -8 32 272
use FILL  FILL_3__2042_
timestamp 1701859473
transform 1 0 8890 0 -1 790
box -12 -8 32 272
use FILL  FILL_3__2043_
timestamp 1701859473
transform 1 0 7210 0 1 270
box -12 -8 32 272
use FILL  FILL_3__2044_
timestamp 1701859473
transform 1 0 6950 0 1 270
box -12 -8 32 272
use FILL  FILL_3__2045_
timestamp 1701859473
transform -1 0 6270 0 1 270
box -12 -8 32 272
use FILL  FILL_3__2046_
timestamp 1701859473
transform 1 0 6450 0 -1 270
box -12 -8 32 272
use FILL  FILL_3__2047_
timestamp 1701859473
transform -1 0 6230 0 -1 270
box -12 -8 32 272
use FILL  FILL_3__2048_
timestamp 1701859473
transform -1 0 6030 0 -1 270
box -12 -8 32 272
use FILL  FILL_3__2049_
timestamp 1701859473
transform -1 0 7210 0 -1 790
box -12 -8 32 272
use FILL  FILL_3__2050_
timestamp 1701859473
transform 1 0 1450 0 -1 2870
box -12 -8 32 272
use FILL  FILL_3__2051_
timestamp 1701859473
transform 1 0 6250 0 -1 2350
box -12 -8 32 272
use FILL  FILL_3__2052_
timestamp 1701859473
transform -1 0 6150 0 1 790
box -12 -8 32 272
use FILL  FILL_3__2053_
timestamp 1701859473
transform -1 0 4370 0 1 1830
box -12 -8 32 272
use FILL  FILL_3__2054_
timestamp 1701859473
transform 1 0 2870 0 1 1310
box -12 -8 32 272
use FILL  FILL_3__2055_
timestamp 1701859473
transform -1 0 3130 0 1 1310
box -12 -8 32 272
use FILL  FILL_3__2056_
timestamp 1701859473
transform -1 0 1850 0 -1 1310
box -12 -8 32 272
use FILL  FILL_3__2057_
timestamp 1701859473
transform 1 0 2710 0 1 790
box -12 -8 32 272
use FILL  FILL_3__2058_
timestamp 1701859473
transform 1 0 3630 0 1 790
box -12 -8 32 272
use FILL  FILL_3__2059_
timestamp 1701859473
transform 1 0 3870 0 1 790
box -12 -8 32 272
use FILL  FILL_3__2060_
timestamp 1701859473
transform -1 0 4110 0 1 790
box -12 -8 32 272
use FILL  FILL_3__2061_
timestamp 1701859473
transform -1 0 2970 0 -1 270
box -12 -8 32 272
use FILL  FILL_3__2062_
timestamp 1701859473
transform 1 0 2750 0 1 270
box -12 -8 32 272
use FILL  FILL_3__2063_
timestamp 1701859473
transform 1 0 3130 0 -1 270
box -12 -8 32 272
use FILL  FILL_3__2064_
timestamp 1701859473
transform 1 0 3370 0 -1 270
box -12 -8 32 272
use FILL  FILL_3__2065_
timestamp 1701859473
transform -1 0 3610 0 -1 270
box -12 -8 32 272
use FILL  FILL_3__2066_
timestamp 1701859473
transform -1 0 5390 0 -1 270
box -12 -8 32 272
use FILL  FILL_3__2067_
timestamp 1701859473
transform 1 0 7330 0 1 790
box -12 -8 32 272
use FILL  FILL_3__2068_
timestamp 1701859473
transform 1 0 5890 0 1 790
box -12 -8 32 272
use FILL  FILL_3__2069_
timestamp 1701859473
transform 1 0 3370 0 -1 1830
box -12 -8 32 272
use FILL  FILL_3__2070_
timestamp 1701859473
transform -1 0 3850 0 -1 1830
box -12 -8 32 272
use FILL  FILL_3__2071_
timestamp 1701859473
transform -1 0 5690 0 1 790
box -12 -8 32 272
use FILL  FILL_3__2072_
timestamp 1701859473
transform -1 0 7750 0 1 1310
box -12 -8 32 272
use FILL  FILL_3__2073_
timestamp 1701859473
transform 1 0 6630 0 1 1310
box -12 -8 32 272
use FILL  FILL_3__2074_
timestamp 1701859473
transform 1 0 1770 0 1 1310
box -12 -8 32 272
use FILL  FILL_3__2075_
timestamp 1701859473
transform -1 0 2250 0 1 1310
box -12 -8 32 272
use FILL  FILL_3__2076_
timestamp 1701859473
transform -1 0 2290 0 -1 1310
box -12 -8 32 272
use FILL  FILL_3__2077_
timestamp 1701859473
transform 1 0 4150 0 -1 1310
box -12 -8 32 272
use FILL  FILL_3__2078_
timestamp 1701859473
transform -1 0 2290 0 1 1830
box -12 -8 32 272
use FILL  FILL_3__2079_
timestamp 1701859473
transform -1 0 930 0 -1 1830
box -12 -8 32 272
use FILL  FILL_3__2080_
timestamp 1701859473
transform 1 0 2250 0 -1 1830
box -12 -8 32 272
use FILL  FILL_3__2081_
timestamp 1701859473
transform 1 0 2490 0 -1 1830
box -12 -8 32 272
use FILL  FILL_3__2082_
timestamp 1701859473
transform -1 0 2710 0 -1 1830
box -12 -8 32 272
use FILL  FILL_3__2083_
timestamp 1701859473
transform 1 0 4390 0 -1 1310
box -12 -8 32 272
use FILL  FILL_3__2084_
timestamp 1701859473
transform -1 0 5230 0 1 790
box -12 -8 32 272
use FILL  FILL_3__2085_
timestamp 1701859473
transform -1 0 5070 0 -1 270
box -12 -8 32 272
use FILL  FILL_3__2086_
timestamp 1701859473
transform -1 0 4290 0 -1 270
box -12 -8 32 272
use FILL  FILL_3__2087_
timestamp 1701859473
transform -1 0 4770 0 1 790
box -12 -8 32 272
use FILL  FILL_3__2088_
timestamp 1701859473
transform -1 0 5610 0 1 270
box -12 -8 32 272
use FILL  FILL_3__2089_
timestamp 1701859473
transform 1 0 5370 0 1 270
box -12 -8 32 272
use FILL  FILL_3__2090_
timestamp 1701859473
transform -1 0 4950 0 -1 790
box -12 -8 32 272
use FILL  FILL_3__2091_
timestamp 1701859473
transform 1 0 3170 0 1 790
box -12 -8 32 272
use FILL  FILL_3__2092_
timestamp 1701859473
transform 1 0 2730 0 -1 270
box -12 -8 32 272
use FILL  FILL_3__2093_
timestamp 1701859473
transform -1 0 2890 0 -1 790
box -12 -8 32 272
use FILL  FILL_3__2094_
timestamp 1701859473
transform 1 0 2290 0 -1 270
box -12 -8 32 272
use FILL  FILL_3__2095_
timestamp 1701859473
transform 1 0 2490 0 -1 270
box -12 -8 32 272
use FILL  FILL_3__2096_
timestamp 1701859473
transform -1 0 4950 0 1 270
box -12 -8 32 272
use FILL  FILL_3__2097_
timestamp 1701859473
transform -1 0 5170 0 1 270
box -12 -8 32 272
use FILL  FILL_3__2098_
timestamp 1701859473
transform 1 0 4710 0 1 270
box -12 -8 32 272
use FILL  FILL_3__2099_
timestamp 1701859473
transform 1 0 4030 0 -1 270
box -12 -8 32 272
use FILL  FILL_3__2100_
timestamp 1701859473
transform -1 0 5890 0 -1 1830
box -12 -8 32 272
use FILL  FILL_3__2101_
timestamp 1701859473
transform -1 0 5810 0 1 1310
box -12 -8 32 272
use FILL  FILL_3__2102_
timestamp 1701859473
transform -1 0 6210 0 1 1310
box -12 -8 32 272
use FILL  FILL_3__2103_
timestamp 1701859473
transform 1 0 5770 0 -1 1310
box -12 -8 32 272
use FILL  FILL_3__2104_
timestamp 1701859473
transform -1 0 6010 0 1 1310
box -12 -8 32 272
use FILL  FILL_3__2105_
timestamp 1701859473
transform -1 0 4310 0 -1 1830
box -12 -8 32 272
use FILL  FILL_3__2106_
timestamp 1701859473
transform 1 0 3990 0 -1 790
box -12 -8 32 272
use FILL  FILL_3__2107_
timestamp 1701859473
transform -1 0 3570 0 -1 790
box -12 -8 32 272
use FILL  FILL_3__2108_
timestamp 1701859473
transform 1 0 2930 0 1 790
box -12 -8 32 272
use FILL  FILL_3__2109_
timestamp 1701859473
transform -1 0 3350 0 -1 790
box -12 -8 32 272
use FILL  FILL_3__2110_
timestamp 1701859473
transform 1 0 3110 0 -1 790
box -12 -8 32 272
use FILL  FILL_3__2111_
timestamp 1701859473
transform -1 0 3790 0 -1 790
box -12 -8 32 272
use FILL  FILL_3__2112_
timestamp 1701859473
transform -1 0 5150 0 -1 790
box -12 -8 32 272
use FILL  FILL_3__2113_
timestamp 1701859473
transform -1 0 5130 0 1 1310
box -12 -8 32 272
use FILL  FILL_3__2114_
timestamp 1701859473
transform -1 0 5570 0 1 1310
box -12 -8 32 272
use FILL  FILL_3__2115_
timestamp 1701859473
transform -1 0 5610 0 -1 790
box -12 -8 32 272
use FILL  FILL_3__2116_
timestamp 1701859473
transform 1 0 2430 0 1 1310
box -12 -8 32 272
use FILL  FILL_3__2117_
timestamp 1701859473
transform 1 0 2630 0 1 1310
box -12 -8 32 272
use FILL  FILL_3__2118_
timestamp 1701859473
transform 1 0 3810 0 1 1310
box -12 -8 32 272
use FILL  FILL_3__2119_
timestamp 1701859473
transform -1 0 4070 0 1 1310
box -12 -8 32 272
use FILL  FILL_3__2120_
timestamp 1701859473
transform 1 0 3930 0 -1 1310
box -12 -8 32 272
use FILL  FILL_3__2121_
timestamp 1701859473
transform -1 0 4510 0 1 270
box -12 -8 32 272
use FILL  FILL_3__2122_
timestamp 1701859473
transform -1 0 2850 0 1 2350
box -12 -8 32 272
use FILL  FILL_3__2123_
timestamp 1701859473
transform 1 0 2790 0 -1 2350
box -12 -8 32 272
use FILL  FILL_3__2124_
timestamp 1701859473
transform -1 0 3690 0 -1 2350
box -12 -8 32 272
use FILL  FILL_3__2125_
timestamp 1701859473
transform 1 0 5810 0 -1 3390
box -12 -8 32 272
use FILL  FILL_3__2126_
timestamp 1701859473
transform 1 0 5490 0 1 2870
box -12 -8 32 272
use FILL  FILL_3__2127_
timestamp 1701859473
transform -1 0 5970 0 1 2870
box -12 -8 32 272
use FILL  FILL_3__2128_
timestamp 1701859473
transform 1 0 4590 0 1 2870
box -12 -8 32 272
use FILL  FILL_3__2129_
timestamp 1701859473
transform 1 0 5270 0 1 2870
box -12 -8 32 272
use FILL  FILL_3__2130_
timestamp 1701859473
transform -1 0 4630 0 -1 2350
box -12 -8 32 272
use FILL  FILL_3__2131_
timestamp 1701859473
transform 1 0 4670 0 1 1310
box -12 -8 32 272
use FILL  FILL_3__2132_
timestamp 1701859473
transform -1 0 4550 0 1 790
box -12 -8 32 272
use FILL  FILL_3__2133_
timestamp 1701859473
transform 1 0 4470 0 -1 790
box -12 -8 32 272
use FILL  FILL_3__2134_
timestamp 1701859473
transform 1 0 3590 0 -1 2870
box -12 -8 32 272
use FILL  FILL_3__2135_
timestamp 1701859473
transform 1 0 4210 0 -1 3390
box -12 -8 32 272
use FILL  FILL_3__2136_
timestamp 1701859473
transform -1 0 2750 0 1 3390
box -12 -8 32 272
use FILL  FILL_3__2137_
timestamp 1701859473
transform 1 0 2310 0 1 3390
box -12 -8 32 272
use FILL  FILL_3__2138_
timestamp 1701859473
transform 1 0 3110 0 -1 4430
box -12 -8 32 272
use FILL  FILL_3__2139_
timestamp 1701859473
transform -1 0 2890 0 -1 4430
box -12 -8 32 272
use FILL  FILL_3__2140_
timestamp 1701859473
transform 1 0 2810 0 1 4430
box -12 -8 32 272
use FILL  FILL_3__2141_
timestamp 1701859473
transform -1 0 3050 0 1 4430
box -12 -8 32 272
use FILL  FILL_3__2142_
timestamp 1701859473
transform 1 0 2930 0 1 3390
box -12 -8 32 272
use FILL  FILL_3__2143_
timestamp 1701859473
transform -1 0 7430 0 -1 3390
box -12 -8 32 272
use FILL  FILL_3__2144_
timestamp 1701859473
transform 1 0 2070 0 1 2870
box -12 -8 32 272
use FILL  FILL_3__2145_
timestamp 1701859473
transform -1 0 10050 0 -1 2870
box -12 -8 32 272
use FILL  FILL_3__2146_
timestamp 1701859473
transform -1 0 7630 0 -1 3390
box -12 -8 32 272
use FILL  FILL_3__2147_
timestamp 1701859473
transform 1 0 7590 0 -1 3910
box -12 -8 32 272
use FILL  FILL_3__2148_
timestamp 1701859473
transform 1 0 7430 0 1 3390
box -12 -8 32 272
use FILL  FILL_3__2149_
timestamp 1701859473
transform 1 0 7630 0 1 3390
box -12 -8 32 272
use FILL  FILL_3__2150_
timestamp 1701859473
transform -1 0 7890 0 1 3390
box -12 -8 32 272
use FILL  FILL_3__2151_
timestamp 1701859473
transform 1 0 7170 0 -1 3390
box -12 -8 32 272
use FILL  FILL_3__2152_
timestamp 1701859473
transform 1 0 6930 0 -1 3390
box -12 -8 32 272
use FILL  FILL_3__2153_
timestamp 1701859473
transform -1 0 6070 0 -1 3390
box -12 -8 32 272
use FILL  FILL_3__2154_
timestamp 1701859473
transform 1 0 2830 0 -1 7030
box -12 -8 32 272
use FILL  FILL_3__2155_
timestamp 1701859473
transform 1 0 6390 0 1 5990
box -12 -8 32 272
use FILL  FILL_3__2156_
timestamp 1701859473
transform -1 0 4610 0 1 3910
box -12 -8 32 272
use FILL  FILL_3__2157_
timestamp 1701859473
transform -1 0 4750 0 -1 4430
box -12 -8 32 272
use FILL  FILL_3__2158_
timestamp 1701859473
transform -1 0 2610 0 1 2350
box -12 -8 32 272
use FILL  FILL_3__2159_
timestamp 1701859473
transform 1 0 3510 0 1 3910
box -12 -8 32 272
use FILL  FILL_3__2160_
timestamp 1701859473
transform -1 0 3830 0 -1 4430
box -12 -8 32 272
use FILL  FILL_3__2161_
timestamp 1701859473
transform -1 0 3970 0 1 3910
box -12 -8 32 272
use FILL  FILL_3__2162_
timestamp 1701859473
transform -1 0 4410 0 1 3910
box -12 -8 32 272
use FILL  FILL_3__2163_
timestamp 1701859473
transform 1 0 3730 0 -1 3910
box -12 -8 32 272
use FILL  FILL_3__2164_
timestamp 1701859473
transform -1 0 550 0 -1 4950
box -12 -8 32 272
use FILL  FILL_3__2165_
timestamp 1701859473
transform -1 0 3250 0 -1 3910
box -12 -8 32 272
use FILL  FILL_3__2166_
timestamp 1701859473
transform 1 0 3950 0 -1 3910
box -12 -8 32 272
use FILL  FILL_3__2167_
timestamp 1701859473
transform 1 0 4150 0 1 3910
box -12 -8 32 272
use FILL  FILL_3__2168_
timestamp 1701859473
transform 1 0 3070 0 1 3910
box -12 -8 32 272
use FILL  FILL_3__2169_
timestamp 1701859473
transform 1 0 2430 0 -1 4430
box -12 -8 32 272
use FILL  FILL_3__2170_
timestamp 1701859473
transform -1 0 2690 0 -1 4430
box -12 -8 32 272
use FILL  FILL_3__2171_
timestamp 1701859473
transform 1 0 4030 0 -1 4430
box -12 -8 32 272
use FILL  FILL_3__2172_
timestamp 1701859473
transform 1 0 4270 0 -1 4430
box -12 -8 32 272
use FILL  FILL_3__2173_
timestamp 1701859473
transform -1 0 4510 0 -1 4430
box -12 -8 32 272
use FILL  FILL_3__2174_
timestamp 1701859473
transform 1 0 6010 0 1 7030
box -12 -8 32 272
use FILL  FILL_3__2175_
timestamp 1701859473
transform -1 0 2510 0 1 8070
box -12 -8 32 272
use FILL  FILL_3__2176_
timestamp 1701859473
transform -1 0 6430 0 -1 8070
box -12 -8 32 272
use FILL  FILL_3__2177_
timestamp 1701859473
transform 1 0 4950 0 1 8070
box -12 -8 32 272
use FILL  FILL_3__2178_
timestamp 1701859473
transform -1 0 4130 0 -1 8590
box -12 -8 32 272
use FILL  FILL_3__2179_
timestamp 1701859473
transform -1 0 5950 0 -1 8070
box -12 -8 32 272
use FILL  FILL_3__2180_
timestamp 1701859473
transform -1 0 2970 0 -1 9630
box -12 -8 32 272
use FILL  FILL_3__2181_
timestamp 1701859473
transform 1 0 5030 0 1 7550
box -12 -8 32 272
use FILL  FILL_3__2182_
timestamp 1701859473
transform 1 0 5550 0 -1 10150
box -12 -8 32 272
use FILL  FILL_3__2183_
timestamp 1701859473
transform -1 0 3530 0 1 10150
box -12 -8 32 272
use FILL  FILL_3__2184_
timestamp 1701859473
transform 1 0 4350 0 1 8070
box -12 -8 32 272
use FILL  FILL_3__2185_
timestamp 1701859473
transform 1 0 5950 0 1 10150
box -12 -8 32 272
use FILL  FILL_3__2186_
timestamp 1701859473
transform 1 0 3510 0 1 10670
box -12 -8 32 272
use FILL  FILL_3__2187_
timestamp 1701859473
transform -1 0 5430 0 -1 10670
box -12 -8 32 272
use FILL  FILL_3__2188_
timestamp 1701859473
transform 1 0 2110 0 -1 10670
box -12 -8 32 272
use FILL  FILL_3__2189_
timestamp 1701859473
transform 1 0 5670 0 -1 10670
box -12 -8 32 272
use FILL  FILL_3__2190_
timestamp 1701859473
transform -1 0 2830 0 1 10150
box -12 -8 32 272
use FILL  FILL_3__2191_
timestamp 1701859473
transform -1 0 5310 0 -1 10150
box -12 -8 32 272
use FILL  FILL_3__2192_
timestamp 1701859473
transform -1 0 11110 0 1 3910
box -12 -8 32 272
use FILL  FILL_3__2193_
timestamp 1701859473
transform 1 0 1230 0 -1 3910
box -12 -8 32 272
use FILL  FILL_3__2194_
timestamp 1701859473
transform 1 0 1030 0 -1 3910
box -12 -8 32 272
use FILL  FILL_3__2195_
timestamp 1701859473
transform 1 0 2610 0 1 3910
box -12 -8 32 272
use FILL  FILL_3__2196_
timestamp 1701859473
transform 1 0 2850 0 1 3910
box -12 -8 32 272
use FILL  FILL_3__2197_
timestamp 1701859473
transform 1 0 5330 0 1 3910
box -12 -8 32 272
use FILL  FILL_3__2198_
timestamp 1701859473
transform 1 0 270 0 1 1830
box -12 -8 32 272
use FILL  FILL_3__2199_
timestamp 1701859473
transform -1 0 2830 0 -1 3910
box -12 -8 32 272
use FILL  FILL_3__2200_
timestamp 1701859473
transform 1 0 5350 0 -1 3910
box -12 -8 32 272
use FILL  FILL_3__2201_
timestamp 1701859473
transform -1 0 5590 0 1 3910
box -12 -8 32 272
use FILL  FILL_3__2202_
timestamp 1701859473
transform -1 0 8170 0 -1 4430
box -12 -8 32 272
use FILL  FILL_3__2203_
timestamp 1701859473
transform -1 0 4890 0 -1 3910
box -12 -8 32 272
use FILL  FILL_3__2204_
timestamp 1701859473
transform 1 0 5110 0 -1 3910
box -12 -8 32 272
use FILL  FILL_3__2205_
timestamp 1701859473
transform -1 0 8970 0 -1 3910
box -12 -8 32 272
use FILL  FILL_3__2206_
timestamp 1701859473
transform 1 0 9050 0 1 3910
box -12 -8 32 272
use FILL  FILL_3__2207_
timestamp 1701859473
transform 1 0 9510 0 -1 3910
box -12 -8 32 272
use FILL  FILL_3__2208_
timestamp 1701859473
transform -1 0 9770 0 -1 3910
box -12 -8 32 272
use FILL  FILL_3__2209_
timestamp 1701859473
transform -1 0 9570 0 1 4430
box -12 -8 32 272
use FILL  FILL_3__2210_
timestamp 1701859473
transform -1 0 10570 0 -1 4950
box -12 -8 32 272
use FILL  FILL_3__2211_
timestamp 1701859473
transform 1 0 9270 0 -1 3910
box -12 -8 32 272
use FILL  FILL_3__2212_
timestamp 1701859473
transform -1 0 8850 0 1 3910
box -12 -8 32 272
use FILL  FILL_3__2213_
timestamp 1701859473
transform -1 0 9290 0 1 3910
box -12 -8 32 272
use FILL  FILL_3__2214_
timestamp 1701859473
transform -1 0 9490 0 -1 4430
box -12 -8 32 272
use FILL  FILL_3__2215_
timestamp 1701859473
transform 1 0 9690 0 -1 4430
box -12 -8 32 272
use FILL  FILL_3__2216_
timestamp 1701859473
transform -1 0 9450 0 -1 7030
box -12 -8 32 272
use FILL  FILL_3__2217_
timestamp 1701859473
transform 1 0 9230 0 -1 4430
box -12 -8 32 272
use FILL  FILL_3__2218_
timestamp 1701859473
transform -1 0 9750 0 1 3910
box -12 -8 32 272
use FILL  FILL_3__2219_
timestamp 1701859473
transform 1 0 9930 0 1 3910
box -12 -8 32 272
use FILL  FILL_3__2220_
timestamp 1701859473
transform 1 0 10310 0 -1 4950
box -12 -8 32 272
use FILL  FILL_3__2221_
timestamp 1701859473
transform -1 0 9690 0 -1 7030
box -12 -8 32 272
use FILL  FILL_3__2222_
timestamp 1701859473
transform 1 0 10050 0 1 4430
box -12 -8 32 272
use FILL  FILL_3__2223_
timestamp 1701859473
transform -1 0 9950 0 -1 4430
box -12 -8 32 272
use FILL  FILL_3__2224_
timestamp 1701859473
transform -1 0 9810 0 1 4430
box -12 -8 32 272
use FILL  FILL_3__2225_
timestamp 1701859473
transform 1 0 10050 0 -1 4950
box -12 -8 32 272
use FILL  FILL_3__2226_
timestamp 1701859473
transform 1 0 8930 0 -1 7030
box -12 -8 32 272
use FILL  FILL_3__2227_
timestamp 1701859473
transform -1 0 9210 0 -1 7030
box -12 -8 32 272
use FILL  FILL_3__2228_
timestamp 1701859473
transform -1 0 5750 0 -1 7030
box -12 -8 32 272
use FILL  FILL_3__2229_
timestamp 1701859473
transform 1 0 4310 0 1 3390
box -12 -8 32 272
use FILL  FILL_3__2230_
timestamp 1701859473
transform -1 0 4410 0 -1 3910
box -12 -8 32 272
use FILL  FILL_3__2231_
timestamp 1701859473
transform -1 0 4190 0 -1 3910
box -12 -8 32 272
use FILL  FILL_3__2232_
timestamp 1701859473
transform 1 0 1590 0 1 2870
box -12 -8 32 272
use FILL  FILL_3__2233_
timestamp 1701859473
transform 1 0 2310 0 1 2870
box -12 -8 32 272
use FILL  FILL_3__2234_
timestamp 1701859473
transform -1 0 2570 0 1 2870
box -12 -8 32 272
use FILL  FILL_3__2235_
timestamp 1701859473
transform 1 0 6330 0 1 3390
box -12 -8 32 272
use FILL  FILL_3__2236_
timestamp 1701859473
transform -1 0 5610 0 -1 3910
box -12 -8 32 272
use FILL  FILL_3__2237_
timestamp 1701859473
transform -1 0 4650 0 -1 3910
box -12 -8 32 272
use FILL  FILL_3__2238_
timestamp 1701859473
transform 1 0 4710 0 -1 4950
box -12 -8 32 272
use FILL  FILL_3__2239_
timestamp 1701859473
transform 1 0 2830 0 1 4950
box -12 -8 32 272
use FILL  FILL_3__2240_
timestamp 1701859473
transform 1 0 2390 0 1 3910
box -12 -8 32 272
use FILL  FILL_3__2241_
timestamp 1701859473
transform -1 0 2410 0 1 4950
box -12 -8 32 272
use FILL  FILL_3__2242_
timestamp 1701859473
transform 1 0 2450 0 -1 4950
box -12 -8 32 272
use FILL  FILL_3__2243_
timestamp 1701859473
transform 1 0 2630 0 1 4950
box -12 -8 32 272
use FILL  FILL_3__2244_
timestamp 1701859473
transform 1 0 3050 0 1 4950
box -12 -8 32 272
use FILL  FILL_3__2245_
timestamp 1701859473
transform 1 0 2890 0 1 5990
box -12 -8 32 272
use FILL  FILL_3__2246_
timestamp 1701859473
transform 1 0 2910 0 -1 4950
box -12 -8 32 272
use FILL  FILL_3__2247_
timestamp 1701859473
transform -1 0 3030 0 -1 6510
box -12 -8 32 272
use FILL  FILL_3__2248_
timestamp 1701859473
transform 1 0 3490 0 -1 7030
box -12 -8 32 272
use FILL  FILL_3__2249_
timestamp 1701859473
transform 1 0 6270 0 1 7030
box -12 -8 32 272
use FILL  FILL_3__2250_
timestamp 1701859473
transform -1 0 10570 0 -1 7550
box -12 -8 32 272
use FILL  FILL_3__2251_
timestamp 1701859473
transform -1 0 10630 0 1 8070
box -12 -8 32 272
use FILL  FILL_3__2252_
timestamp 1701859473
transform -1 0 10930 0 -1 8070
box -12 -8 32 272
use FILL  FILL_3__2253_
timestamp 1701859473
transform -1 0 10690 0 -1 8070
box -12 -8 32 272
use FILL  FILL_3__2254_
timestamp 1701859473
transform 1 0 5390 0 1 8070
box -12 -8 32 272
use FILL  FILL_3__2255_
timestamp 1701859473
transform 1 0 3010 0 1 7030
box -12 -8 32 272
use FILL  FILL_3__2256_
timestamp 1701859473
transform -1 0 5130 0 1 7030
box -12 -8 32 272
use FILL  FILL_3__2257_
timestamp 1701859473
transform 1 0 5070 0 -1 7550
box -12 -8 32 272
use FILL  FILL_3__2258_
timestamp 1701859473
transform 1 0 5710 0 -1 8590
box -12 -8 32 272
use FILL  FILL_3__2259_
timestamp 1701859473
transform 1 0 10330 0 -1 7550
box -12 -8 32 272
use FILL  FILL_3__2260_
timestamp 1701859473
transform 1 0 9910 0 1 8070
box -12 -8 32 272
use FILL  FILL_3__2261_
timestamp 1701859473
transform -1 0 10210 0 1 7550
box -12 -8 32 272
use FILL  FILL_3__2262_
timestamp 1701859473
transform -1 0 9970 0 1 7550
box -12 -8 32 272
use FILL  FILL_3__2263_
timestamp 1701859473
transform 1 0 5470 0 1 7550
box -12 -8 32 272
use FILL  FILL_3__2264_
timestamp 1701859473
transform 1 0 1630 0 -1 6510
box -12 -8 32 272
use FILL  FILL_3__2265_
timestamp 1701859473
transform 1 0 1810 0 -1 6510
box -12 -8 32 272
use FILL  FILL_3__2266_
timestamp 1701859473
transform 1 0 3910 0 1 6510
box -12 -8 32 272
use FILL  FILL_3__2267_
timestamp 1701859473
transform -1 0 3670 0 -1 7550
box -12 -8 32 272
use FILL  FILL_3__2268_
timestamp 1701859473
transform 1 0 4350 0 -1 7550
box -12 -8 32 272
use FILL  FILL_3__2269_
timestamp 1701859473
transform 1 0 5670 0 1 7550
box -12 -8 32 272
use FILL  FILL_3__2270_
timestamp 1701859473
transform 1 0 8590 0 1 7550
box -12 -8 32 272
use FILL  FILL_3__2271_
timestamp 1701859473
transform -1 0 8870 0 -1 8070
box -12 -8 32 272
use FILL  FILL_3__2272_
timestamp 1701859473
transform -1 0 9130 0 -1 8070
box -12 -8 32 272
use FILL  FILL_3__2273_
timestamp 1701859473
transform -1 0 8630 0 -1 8070
box -12 -8 32 272
use FILL  FILL_3__2274_
timestamp 1701859473
transform -1 0 5990 0 -1 9630
box -12 -8 32 272
use FILL  FILL_3__2275_
timestamp 1701859473
transform -1 0 2290 0 1 8070
box -12 -8 32 272
use FILL  FILL_3__2276_
timestamp 1701859473
transform -1 0 3170 0 1 8070
box -12 -8 32 272
use FILL  FILL_3__2277_
timestamp 1701859473
transform -1 0 3650 0 -1 8590
box -12 -8 32 272
use FILL  FILL_3__2278_
timestamp 1701859473
transform 1 0 6550 0 1 9110
box -12 -8 32 272
use FILL  FILL_3__2279_
timestamp 1701859473
transform -1 0 10250 0 1 5990
box -12 -8 32 272
use FILL  FILL_3__2280_
timestamp 1701859473
transform 1 0 10430 0 1 5990
box -12 -8 32 272
use FILL  FILL_3__2281_
timestamp 1701859473
transform -1 0 10710 0 -1 5990
box -12 -8 32 272
use FILL  FILL_3__2282_
timestamp 1701859473
transform -1 0 10490 0 -1 6510
box -12 -8 32 272
use FILL  FILL_3__2283_
timestamp 1701859473
transform 1 0 5950 0 -1 8590
box -12 -8 32 272
use FILL  FILL_3__2284_
timestamp 1701859473
transform -1 0 2070 0 1 8070
box -12 -8 32 272
use FILL  FILL_3__2285_
timestamp 1701859473
transform -1 0 4130 0 1 8070
box -12 -8 32 272
use FILL  FILL_3__2286_
timestamp 1701859473
transform 1 0 5030 0 -1 8590
box -12 -8 32 272
use FILL  FILL_3__2287_
timestamp 1701859473
transform -1 0 6110 0 1 8590
box -12 -8 32 272
use FILL  FILL_3__2288_
timestamp 1701859473
transform -1 0 8830 0 1 7550
box -12 -8 32 272
use FILL  FILL_3__2289_
timestamp 1701859473
transform 1 0 8490 0 1 8070
box -12 -8 32 272
use FILL  FILL_3__2290_
timestamp 1701859473
transform -1 0 9990 0 -1 8070
box -12 -8 32 272
use FILL  FILL_3__2291_
timestamp 1701859473
transform -1 0 8770 0 1 8070
box -12 -8 32 272
use FILL  FILL_3__2292_
timestamp 1701859473
transform -1 0 6210 0 -1 9110
box -12 -8 32 272
use FILL  FILL_3__2293_
timestamp 1701859473
transform -1 0 2530 0 -1 8590
box -12 -8 32 272
use FILL  FILL_3__2294_
timestamp 1701859473
transform -1 0 4010 0 1 8590
box -12 -8 32 272
use FILL  FILL_3__2295_
timestamp 1701859473
transform 1 0 4930 0 1 8590
box -12 -8 32 272
use FILL  FILL_3__2296_
timestamp 1701859473
transform 1 0 6650 0 -1 9110
box -12 -8 32 272
use FILL  FILL_3__2297_
timestamp 1701859473
transform -1 0 9550 0 -1 5990
box -12 -8 32 272
use FILL  FILL_3__2298_
timestamp 1701859473
transform -1 0 9990 0 -1 5470
box -12 -8 32 272
use FILL  FILL_3__2299_
timestamp 1701859473
transform -1 0 9330 0 -1 6510
box -12 -8 32 272
use FILL  FILL_3__2300_
timestamp 1701859473
transform 1 0 9530 0 1 5990
box -12 -8 32 272
use FILL  FILL_3__2301_
timestamp 1701859473
transform 1 0 5570 0 1 9630
box -12 -8 32 272
use FILL  FILL_3__2302_
timestamp 1701859473
transform -1 0 3470 0 -1 9110
box -12 -8 32 272
use FILL  FILL_3__2303_
timestamp 1701859473
transform 1 0 2590 0 1 9110
box -12 -8 32 272
use FILL  FILL_3__2304_
timestamp 1701859473
transform 1 0 2790 0 -1 9110
box -12 -8 32 272
use FILL  FILL_3__2305_
timestamp 1701859473
transform -1 0 3770 0 1 8590
box -12 -8 32 272
use FILL  FILL_3__2306_
timestamp 1701859473
transform 1 0 4450 0 1 8590
box -12 -8 32 272
use FILL  FILL_3__2307_
timestamp 1701859473
transform 1 0 6310 0 1 9110
box -12 -8 32 272
use FILL  FILL_3__2308_
timestamp 1701859473
transform -1 0 8890 0 -1 6510
box -12 -8 32 272
use FILL  FILL_3__2309_
timestamp 1701859473
transform -1 0 8590 0 1 5990
box -12 -8 32 272
use FILL  FILL_3__2310_
timestamp 1701859473
transform -1 0 9090 0 -1 6510
box -12 -8 32 272
use FILL  FILL_3__2311_
timestamp 1701859473
transform -1 0 8650 0 -1 6510
box -12 -8 32 272
use FILL  FILL_3__2312_
timestamp 1701859473
transform -1 0 5550 0 -1 9630
box -12 -8 32 272
use FILL  FILL_3__2313_
timestamp 1701859473
transform -1 0 1830 0 1 8590
box -12 -8 32 272
use FILL  FILL_3__2314_
timestamp 1701859473
transform 1 0 1430 0 -1 8590
box -12 -8 32 272
use FILL  FILL_3__2315_
timestamp 1701859473
transform 1 0 1870 0 -1 8590
box -12 -8 32 272
use FILL  FILL_3__2316_
timestamp 1701859473
transform -1 0 4230 0 1 8590
box -12 -8 32 272
use FILL  FILL_3__2317_
timestamp 1701859473
transform 1 0 4690 0 1 8590
box -12 -8 32 272
use FILL  FILL_3__2318_
timestamp 1701859473
transform 1 0 6790 0 1 9110
box -12 -8 32 272
use FILL  FILL_3__2319_
timestamp 1701859473
transform -1 0 11110 0 1 4430
box -12 -8 32 272
use FILL  FILL_3__2320_
timestamp 1701859473
transform 1 0 5090 0 1 3910
box -12 -8 32 272
use FILL  FILL_3__2321_
timestamp 1701859473
transform 1 0 6510 0 1 3910
box -12 -8 32 272
use FILL  FILL_3__2322_
timestamp 1701859473
transform -1 0 7890 0 1 3910
box -12 -8 32 272
use FILL  FILL_3__2323_
timestamp 1701859473
transform 1 0 7930 0 -1 4430
box -12 -8 32 272
use FILL  FILL_3__2324_
timestamp 1701859473
transform -1 0 11150 0 -1 2870
box -12 -8 32 272
use FILL  FILL_3__2325_
timestamp 1701859473
transform -1 0 8130 0 1 3910
box -12 -8 32 272
use FILL  FILL_3__2326_
timestamp 1701859473
transform -1 0 3170 0 -1 4950
box -12 -8 32 272
use FILL  FILL_3__2327_
timestamp 1701859473
transform -1 0 3370 0 -1 4950
box -12 -8 32 272
use FILL  FILL_3__2328_
timestamp 1701859473
transform 1 0 3850 0 -1 5470
box -12 -8 32 272
use FILL  FILL_3__2329_
timestamp 1701859473
transform 1 0 3610 0 -1 5470
box -12 -8 32 272
use FILL  FILL_3__2330_
timestamp 1701859473
transform 1 0 3750 0 1 4950
box -12 -8 32 272
use FILL  FILL_3__2331_
timestamp 1701859473
transform 1 0 4830 0 1 3910
box -12 -8 32 272
use FILL  FILL_3__2332_
timestamp 1701859473
transform -1 0 4170 0 1 4950
box -12 -8 32 272
use FILL  FILL_3__2333_
timestamp 1701859473
transform -1 0 11130 0 -1 4430
box -12 -8 32 272
use FILL  FILL_3__2334_
timestamp 1701859473
transform 1 0 9010 0 -1 4430
box -12 -8 32 272
use FILL  FILL_3__2335_
timestamp 1701859473
transform 1 0 5190 0 -1 5470
box -12 -8 32 272
use FILL  FILL_3__2336_
timestamp 1701859473
transform -1 0 5050 0 1 5990
box -12 -8 32 272
use FILL  FILL_3__2337_
timestamp 1701859473
transform 1 0 4550 0 1 3390
box -12 -8 32 272
use FILL  FILL_3__2338_
timestamp 1701859473
transform 1 0 3150 0 1 3390
box -12 -8 32 272
use FILL  FILL_3__2339_
timestamp 1701859473
transform 1 0 4730 0 1 3390
box -12 -8 32 272
use FILL  FILL_3__2340_
timestamp 1701859473
transform 1 0 4970 0 1 3390
box -12 -8 32 272
use FILL  FILL_3__2341_
timestamp 1701859473
transform -1 0 550 0 1 5990
box -12 -8 32 272
use FILL  FILL_3__2342_
timestamp 1701859473
transform 1 0 2650 0 1 5470
box -12 -8 32 272
use FILL  FILL_3__2343_
timestamp 1701859473
transform -1 0 4590 0 1 6510
box -12 -8 32 272
use FILL  FILL_3__2344_
timestamp 1701859473
transform -1 0 4870 0 1 5470
box -12 -8 32 272
use FILL  FILL_3__2345_
timestamp 1701859473
transform -1 0 4670 0 1 5470
box -12 -8 32 272
use FILL  FILL_3__2346_
timestamp 1701859473
transform -1 0 4830 0 -1 5990
box -12 -8 32 272
use FILL  FILL_3__2347_
timestamp 1701859473
transform -1 0 5690 0 -1 5990
box -12 -8 32 272
use FILL  FILL_3__2348_
timestamp 1701859473
transform 1 0 5250 0 -1 6510
box -12 -8 32 272
use FILL  FILL_3__2349_
timestamp 1701859473
transform -1 0 5030 0 -1 6510
box -12 -8 32 272
use FILL  FILL_3__2350_
timestamp 1701859473
transform -1 0 4450 0 -1 6510
box -12 -8 32 272
use FILL  FILL_3__2351_
timestamp 1701859473
transform 1 0 5590 0 1 7030
box -12 -8 32 272
use FILL  FILL_3__2352_
timestamp 1701859473
transform -1 0 5810 0 1 7030
box -12 -8 32 272
use FILL  FILL_3__2353_
timestamp 1701859473
transform -1 0 750 0 1 7030
box -12 -8 32 272
use FILL  FILL_3__2354_
timestamp 1701859473
transform 1 0 5450 0 -1 5990
box -12 -8 32 272
use FILL  FILL_3__2355_
timestamp 1701859473
transform 1 0 5350 0 1 7030
box -12 -8 32 272
use FILL  FILL_3__2356_
timestamp 1701859473
transform -1 0 4850 0 -1 7550
box -12 -8 32 272
use FILL  FILL_3__2357_
timestamp 1701859473
transform 1 0 4710 0 1 8070
box -12 -8 32 272
use FILL  FILL_3__2358_
timestamp 1701859473
transform 1 0 5190 0 1 8070
box -12 -8 32 272
use FILL  FILL_3__2359_
timestamp 1701859473
transform -1 0 5510 0 -1 8590
box -12 -8 32 272
use FILL  FILL_3__2360_
timestamp 1701859473
transform -1 0 750 0 -1 6510
box -12 -8 32 272
use FILL  FILL_3__2361_
timestamp 1701859473
transform -1 0 5250 0 1 5990
box -12 -8 32 272
use FILL  FILL_3__2362_
timestamp 1701859473
transform 1 0 5250 0 1 6510
box -12 -8 32 272
use FILL  FILL_3__2363_
timestamp 1701859473
transform 1 0 5270 0 -1 7030
box -12 -8 32 272
use FILL  FILL_3__2364_
timestamp 1701859473
transform 1 0 5270 0 -1 8070
box -12 -8 32 272
use FILL  FILL_3__2365_
timestamp 1701859473
transform 1 0 5510 0 -1 8070
box -12 -8 32 272
use FILL  FILL_3__2366_
timestamp 1701859473
transform -1 0 5730 0 -1 8070
box -12 -8 32 272
use FILL  FILL_3__2367_
timestamp 1701859473
transform 1 0 2690 0 -1 7550
box -12 -8 32 272
use FILL  FILL_3__2368_
timestamp 1701859473
transform -1 0 5530 0 -1 7030
box -12 -8 32 272
use FILL  FILL_3__2369_
timestamp 1701859473
transform 1 0 5230 0 1 7550
box -12 -8 32 272
use FILL  FILL_3__2370_
timestamp 1701859473
transform -1 0 5270 0 -1 8590
box -12 -8 32 272
use FILL  FILL_3__2371_
timestamp 1701859473
transform 1 0 5950 0 -1 9110
box -12 -8 32 272
use FILL  FILL_3__2372_
timestamp 1701859473
transform 1 0 6110 0 1 9110
box -12 -8 32 272
use FILL  FILL_3__2373_
timestamp 1701859473
transform -1 0 6190 0 -1 9630
box -12 -8 32 272
use FILL  FILL_3__2374_
timestamp 1701859473
transform 1 0 70 0 -1 9110
box -12 -8 32 272
use FILL  FILL_3__2375_
timestamp 1701859473
transform -1 0 4210 0 1 5470
box -12 -8 32 272
use FILL  FILL_3__2376_
timestamp 1701859473
transform 1 0 4550 0 -1 5990
box -12 -8 32 272
use FILL  FILL_3__2377_
timestamp 1701859473
transform -1 0 3970 0 -1 6510
box -12 -8 32 272
use FILL  FILL_3__2378_
timestamp 1701859473
transform 1 0 3710 0 -1 6510
box -12 -8 32 272
use FILL  FILL_3__2379_
timestamp 1701859473
transform -1 0 5030 0 1 6510
box -12 -8 32 272
use FILL  FILL_3__2380_
timestamp 1701859473
transform -1 0 4810 0 -1 8590
box -12 -8 32 272
use FILL  FILL_3__2381_
timestamp 1701859473
transform 1 0 3870 0 -1 8590
box -12 -8 32 272
use FILL  FILL_3__2382_
timestamp 1701859473
transform -1 0 4570 0 -1 8590
box -12 -8 32 272
use FILL  FILL_3__2383_
timestamp 1701859473
transform -1 0 5650 0 1 8590
box -12 -8 32 272
use FILL  FILL_3__2384_
timestamp 1701859473
transform -1 0 5870 0 1 8590
box -12 -8 32 272
use FILL  FILL_3__2385_
timestamp 1701859473
transform 1 0 1250 0 -1 10150
box -12 -8 32 272
use FILL  FILL_3__2386_
timestamp 1701859473
transform 1 0 5510 0 -1 7550
box -12 -8 32 272
use FILL  FILL_3__2387_
timestamp 1701859473
transform 1 0 5490 0 -1 9110
box -12 -8 32 272
use FILL  FILL_3__2388_
timestamp 1701859473
transform -1 0 5290 0 -1 9110
box -12 -8 32 272
use FILL  FILL_3__2389_
timestamp 1701859473
transform -1 0 5070 0 -1 9630
box -12 -8 32 272
use FILL  FILL_3__2390_
timestamp 1701859473
transform 1 0 5130 0 1 9630
box -12 -8 32 272
use FILL  FILL_3__2391_
timestamp 1701859473
transform -1 0 5350 0 1 9630
box -12 -8 32 272
use FILL  FILL_3__2392_
timestamp 1701859473
transform 1 0 1450 0 -1 10150
box -12 -8 32 272
use FILL  FILL_3__2393_
timestamp 1701859473
transform -1 0 5310 0 -1 7550
box -12 -8 32 272
use FILL  FILL_3__2394_
timestamp 1701859473
transform 1 0 5390 0 1 8590
box -12 -8 32 272
use FILL  FILL_3__2395_
timestamp 1701859473
transform -1 0 5750 0 -1 9110
box -12 -8 32 272
use FILL  FILL_3__2396_
timestamp 1701859473
transform 1 0 5670 0 1 9110
box -12 -8 32 272
use FILL  FILL_3__2397_
timestamp 1701859473
transform 1 0 5910 0 1 9110
box -12 -8 32 272
use FILL  FILL_3__2398_
timestamp 1701859473
transform 1 0 5730 0 -1 9630
box -12 -8 32 272
use FILL  FILL_3__2399_
timestamp 1701859473
transform -1 0 3170 0 -1 5470
box -12 -8 32 272
use FILL  FILL_3__2400_
timestamp 1701859473
transform -1 0 3350 0 1 5990
box -12 -8 32 272
use FILL  FILL_3__2401_
timestamp 1701859473
transform 1 0 3270 0 -1 6510
box -12 -8 32 272
use FILL  FILL_3__2402_
timestamp 1701859473
transform -1 0 2210 0 -1 4430
box -12 -8 32 272
use FILL  FILL_3__2403_
timestamp 1701859473
transform -1 0 2610 0 1 4430
box -12 -8 32 272
use FILL  FILL_3__2404_
timestamp 1701859473
transform -1 0 2930 0 -1 5470
box -12 -8 32 272
use FILL  FILL_3__2405_
timestamp 1701859473
transform 1 0 2310 0 -1 2870
box -12 -8 32 272
use FILL  FILL_3__2406_
timestamp 1701859473
transform 1 0 3010 0 -1 3390
box -12 -8 32 272
use FILL  FILL_3__2407_
timestamp 1701859473
transform -1 0 3150 0 1 5470
box -12 -8 32 272
use FILL  FILL_3__2408_
timestamp 1701859473
transform 1 0 770 0 -1 2870
box -12 -8 32 272
use FILL  FILL_3__2409_
timestamp 1701859473
transform 1 0 790 0 -1 3910
box -12 -8 32 272
use FILL  FILL_3__2410_
timestamp 1701859473
transform 1 0 1190 0 1 4430
box -12 -8 32 272
use FILL  FILL_3__2411_
timestamp 1701859473
transform -1 0 750 0 -1 4950
box -12 -8 32 272
use FILL  FILL_3__2412_
timestamp 1701859473
transform 1 0 2430 0 -1 5990
box -12 -8 32 272
use FILL  FILL_3__2413_
timestamp 1701859473
transform 1 0 2890 0 1 5470
box -12 -8 32 272
use FILL  FILL_3__2414_
timestamp 1701859473
transform 1 0 4050 0 -1 5470
box -12 -8 32 272
use FILL  FILL_3__2415_
timestamp 1701859473
transform -1 0 3990 0 1 7030
box -12 -8 32 272
use FILL  FILL_3__2416_
timestamp 1701859473
transform 1 0 3950 0 1 4950
box -12 -8 32 272
use FILL  FILL_3__2417_
timestamp 1701859473
transform 1 0 4290 0 -1 5470
box -12 -8 32 272
use FILL  FILL_3__2418_
timestamp 1701859473
transform -1 0 1550 0 -1 4950
box -12 -8 32 272
use FILL  FILL_3__2419_
timestamp 1701859473
transform 1 0 2130 0 1 4430
box -12 -8 32 272
use FILL  FILL_3__2420_
timestamp 1701859473
transform 1 0 3790 0 1 5990
box -12 -8 32 272
use FILL  FILL_3__2421_
timestamp 1701859473
transform -1 0 3570 0 1 5990
box -12 -8 32 272
use FILL  FILL_3__2422_
timestamp 1701859473
transform -1 0 3450 0 -1 5990
box -12 -8 32 272
use FILL  FILL_3__2423_
timestamp 1701859473
transform -1 0 3670 0 -1 5990
box -12 -8 32 272
use FILL  FILL_3__2424_
timestamp 1701859473
transform 1 0 3210 0 -1 5990
box -12 -8 32 272
use FILL  FILL_3__2425_
timestamp 1701859473
transform 1 0 4350 0 1 5990
box -12 -8 32 272
use FILL  FILL_3__2426_
timestamp 1701859473
transform 1 0 3950 0 -1 7030
box -12 -8 32 272
use FILL  FILL_3__2427_
timestamp 1701859473
transform 1 0 4770 0 1 5990
box -12 -8 32 272
use FILL  FILL_3__2428_
timestamp 1701859473
transform 1 0 4530 0 1 5990
box -12 -8 32 272
use FILL  FILL_3__2429_
timestamp 1701859473
transform -1 0 4210 0 -1 6510
box -12 -8 32 272
use FILL  FILL_3__2430_
timestamp 1701859473
transform 1 0 4770 0 1 6510
box -12 -8 32 272
use FILL  FILL_3__2431_
timestamp 1701859473
transform -1 0 4870 0 -1 7030
box -12 -8 32 272
use FILL  FILL_3__2432_
timestamp 1701859473
transform 1 0 5090 0 -1 7030
box -12 -8 32 272
use FILL  FILL_3__2433_
timestamp 1701859473
transform -1 0 4350 0 -1 8070
box -12 -8 32 272
use FILL  FILL_3__2434_
timestamp 1701859473
transform 1 0 4830 0 1 7550
box -12 -8 32 272
use FILL  FILL_3__2435_
timestamp 1701859473
transform 1 0 4170 0 1 7030
box -12 -8 32 272
use FILL  FILL_3__2436_
timestamp 1701859473
transform -1 0 4610 0 -1 7550
box -12 -8 32 272
use FILL  FILL_3__2437_
timestamp 1701859473
transform -1 0 4590 0 -1 8070
box -12 -8 32 272
use FILL  FILL_3__2438_
timestamp 1701859473
transform -1 0 4830 0 -1 8070
box -12 -8 32 272
use FILL  FILL_3__2439_
timestamp 1701859473
transform -1 0 5070 0 -1 8070
box -12 -8 32 272
use FILL  FILL_3__2440_
timestamp 1701859473
transform 1 0 4610 0 1 10150
box -12 -8 32 272
use FILL  FILL_3__2441_
timestamp 1701859473
transform 1 0 3890 0 -1 7550
box -12 -8 32 272
use FILL  FILL_3__2442_
timestamp 1701859473
transform -1 0 4110 0 -1 8070
box -12 -8 32 272
use FILL  FILL_3__2443_
timestamp 1701859473
transform -1 0 3890 0 1 8070
box -12 -8 32 272
use FILL  FILL_3__2444_
timestamp 1701859473
transform 1 0 3630 0 1 8070
box -12 -8 32 272
use FILL  FILL_3__2445_
timestamp 1701859473
transform -1 0 4610 0 1 7550
box -12 -8 32 272
use FILL  FILL_3__2446_
timestamp 1701859473
transform 1 0 4530 0 1 8070
box -12 -8 32 272
use FILL  FILL_3__2447_
timestamp 1701859473
transform 1 0 4270 0 1 9110
box -12 -8 32 272
use FILL  FILL_3__2448_
timestamp 1701859473
transform 1 0 4930 0 1 9110
box -12 -8 32 272
use FILL  FILL_3__2449_
timestamp 1701859473
transform 1 0 5190 0 1 9110
box -12 -8 32 272
use FILL  FILL_3__2450_
timestamp 1701859473
transform 1 0 5430 0 1 9110
box -12 -8 32 272
use FILL  FILL_3__2451_
timestamp 1701859473
transform -1 0 5310 0 -1 9630
box -12 -8 32 272
use FILL  FILL_3__2452_
timestamp 1701859473
transform -1 0 5230 0 -1 10670
box -12 -8 32 272
use FILL  FILL_3__2453_
timestamp 1701859473
transform 1 0 3770 0 -1 10150
box -12 -8 32 272
use FILL  FILL_3__2454_
timestamp 1701859473
transform 1 0 3890 0 1 7550
box -12 -8 32 272
use FILL  FILL_3__2455_
timestamp 1701859473
transform 1 0 3850 0 -1 8070
box -12 -8 32 272
use FILL  FILL_3__2456_
timestamp 1701859473
transform -1 0 3630 0 -1 8070
box -12 -8 32 272
use FILL  FILL_3__2457_
timestamp 1701859473
transform 1 0 3390 0 1 8070
box -12 -8 32 272
use FILL  FILL_3__2458_
timestamp 1701859473
transform -1 0 4330 0 -1 8590
box -12 -8 32 272
use FILL  FILL_3__2459_
timestamp 1701859473
transform -1 0 4490 0 -1 11190
box -12 -8 32 272
use FILL  FILL_3__2460_
timestamp 1701859473
transform 1 0 4130 0 -1 10670
box -12 -8 32 272
use FILL  FILL_3__2461_
timestamp 1701859473
transform 1 0 4310 0 -1 9110
box -12 -8 32 272
use FILL  FILL_3__2462_
timestamp 1701859473
transform -1 0 4570 0 -1 9110
box -12 -8 32 272
use FILL  FILL_3__2463_
timestamp 1701859473
transform -1 0 4810 0 -1 9110
box -12 -8 32 272
use FILL  FILL_3__2464_
timestamp 1701859473
transform -1 0 5050 0 -1 9110
box -12 -8 32 272
use FILL  FILL_3__2465_
timestamp 1701859473
transform -1 0 4910 0 -1 11190
box -12 -8 32 272
use FILL  FILL_3__2466_
timestamp 1701859473
transform -1 0 3990 0 -1 10150
box -12 -8 32 272
use FILL  FILL_3__2467_
timestamp 1701859473
transform -1 0 4090 0 -1 9630
box -12 -8 32 272
use FILL  FILL_3__2468_
timestamp 1701859473
transform -1 0 4350 0 -1 9630
box -12 -8 32 272
use FILL  FILL_3__2469_
timestamp 1701859473
transform -1 0 4210 0 1 9630
box -12 -8 32 272
use FILL  FILL_3__2470_
timestamp 1701859473
transform -1 0 4450 0 1 9630
box -12 -8 32 272
use FILL  FILL_3__2471_
timestamp 1701859473
transform -1 0 5030 0 -1 10670
box -12 -8 32 272
use FILL  FILL_3__2472_
timestamp 1701859473
transform 1 0 3990 0 1 9630
box -12 -8 32 272
use FILL  FILL_3__2473_
timestamp 1701859473
transform 1 0 4550 0 -1 9630
box -12 -8 32 272
use FILL  FILL_3__2474_
timestamp 1701859473
transform -1 0 4830 0 -1 9630
box -12 -8 32 272
use FILL  FILL_3__2475_
timestamp 1701859473
transform 1 0 4670 0 1 9630
box -12 -8 32 272
use FILL  FILL_3__2476_
timestamp 1701859473
transform -1 0 4910 0 1 9630
box -12 -8 32 272
use FILL  FILL_3__2477_
timestamp 1701859473
transform 1 0 4850 0 1 10670
box -12 -8 32 272
use FILL  FILL_3__2478_
timestamp 1701859473
transform 1 0 3090 0 1 5990
box -12 -8 32 272
use FILL  FILL_3__2479_
timestamp 1701859473
transform -1 0 2650 0 1 5990
box -12 -8 32 272
use FILL  FILL_3__2480_
timestamp 1701859473
transform -1 0 2670 0 -1 5990
box -12 -8 32 272
use FILL  FILL_3__2481_
timestamp 1701859473
transform -1 0 2910 0 -1 5990
box -12 -8 32 272
use FILL  FILL_3__2482_
timestamp 1701859473
transform 1 0 1490 0 -1 5990
box -12 -8 32 272
use FILL  FILL_3__2483_
timestamp 1701859473
transform 1 0 2310 0 1 6510
box -12 -8 32 272
use FILL  FILL_3__2484_
timestamp 1701859473
transform -1 0 1930 0 1 6510
box -12 -8 32 272
use FILL  FILL_3__2485_
timestamp 1701859473
transform -1 0 2130 0 1 6510
box -12 -8 32 272
use FILL  FILL_3__2486_
timestamp 1701859473
transform 1 0 2330 0 -1 7030
box -12 -8 32 272
use FILL  FILL_3__2487_
timestamp 1701859473
transform 1 0 2090 0 -1 7030
box -12 -8 32 272
use FILL  FILL_3__2488_
timestamp 1701859473
transform -1 0 1890 0 -1 7030
box -12 -8 32 272
use FILL  FILL_3__2489_
timestamp 1701859473
transform 1 0 1390 0 -1 7030
box -12 -8 32 272
use FILL  FILL_3__2490_
timestamp 1701859473
transform -1 0 990 0 1 5470
box -12 -8 32 272
use FILL  FILL_3__2491_
timestamp 1701859473
transform 1 0 1190 0 1 5470
box -12 -8 32 272
use FILL  FILL_3__2492_
timestamp 1701859473
transform -1 0 2050 0 -1 6510
box -12 -8 32 272
use FILL  FILL_3__2493_
timestamp 1701859473
transform 1 0 1930 0 1 5990
box -12 -8 32 272
use FILL  FILL_3__2494_
timestamp 1701859473
transform -1 0 1490 0 1 5990
box -12 -8 32 272
use FILL  FILL_3__2495_
timestamp 1701859473
transform 1 0 1230 0 1 5990
box -12 -8 32 272
use FILL  FILL_3__2496_
timestamp 1701859473
transform 1 0 1630 0 -1 7030
box -12 -8 32 272
use FILL  FILL_3__2497_
timestamp 1701859473
transform -1 0 1830 0 -1 7550
box -12 -8 32 272
use FILL  FILL_3__2498_
timestamp 1701859473
transform 1 0 770 0 1 8070
box -12 -8 32 272
use FILL  FILL_3__2499_
timestamp 1701859473
transform 1 0 2450 0 1 7550
box -12 -8 32 272
use FILL  FILL_3__2500_
timestamp 1701859473
transform 1 0 1870 0 1 7550
box -12 -8 32 272
use FILL  FILL_3__2501_
timestamp 1701859473
transform 1 0 1650 0 1 7550
box -12 -8 32 272
use FILL  FILL_3__2502_
timestamp 1701859473
transform -1 0 1190 0 1 7550
box -12 -8 32 272
use FILL  FILL_3__2503_
timestamp 1701859473
transform -1 0 1430 0 1 8070
box -12 -8 32 272
use FILL  FILL_3__2504_
timestamp 1701859473
transform -1 0 1850 0 1 8070
box -12 -8 32 272
use FILL  FILL_3__2505_
timestamp 1701859473
transform 1 0 1190 0 1 8070
box -12 -8 32 272
use FILL  FILL_3__2506_
timestamp 1701859473
transform -1 0 1710 0 -1 8070
box -12 -8 32 272
use FILL  FILL_3__2507_
timestamp 1701859473
transform 1 0 1450 0 -1 8070
box -12 -8 32 272
use FILL  FILL_3__2508_
timestamp 1701859473
transform 1 0 970 0 1 8070
box -12 -8 32 272
use FILL  FILL_3__2509_
timestamp 1701859473
transform 1 0 530 0 -1 8590
box -12 -8 32 272
use FILL  FILL_3__2510_
timestamp 1701859473
transform -1 0 1470 0 1 9110
box -12 -8 32 272
use FILL  FILL_3__2511_
timestamp 1701859473
transform -1 0 1410 0 -1 9630
box -12 -8 32 272
use FILL  FILL_3__2512_
timestamp 1701859473
transform 1 0 970 0 -1 9630
box -12 -8 32 272
use FILL  FILL_3__2513_
timestamp 1701859473
transform -1 0 970 0 1 8590
box -12 -8 32 272
use FILL  FILL_3__2514_
timestamp 1701859473
transform 1 0 2050 0 -1 8590
box -12 -8 32 272
use FILL  FILL_3__2515_
timestamp 1701859473
transform 1 0 1170 0 -1 9110
box -12 -8 32 272
use FILL  FILL_3__2516_
timestamp 1701859473
transform -1 0 1010 0 1 9110
box -12 -8 32 272
use FILL  FILL_3__2517_
timestamp 1701859473
transform -1 0 770 0 1 9110
box -12 -8 32 272
use FILL  FILL_3__2518_
timestamp 1701859473
transform 1 0 1630 0 -1 9630
box -12 -8 32 272
use FILL  FILL_3__2519_
timestamp 1701859473
transform 1 0 1730 0 1 9630
box -12 -8 32 272
use FILL  FILL_3__2520_
timestamp 1701859473
transform -1 0 2570 0 -1 9110
box -12 -8 32 272
use FILL  FILL_3__2521_
timestamp 1701859473
transform 1 0 2310 0 -1 9110
box -12 -8 32 272
use FILL  FILL_3__2522_
timestamp 1701859473
transform -1 0 1930 0 1 9630
box -12 -8 32 272
use FILL  FILL_3__2523_
timestamp 1701859473
transform -1 0 2150 0 1 9630
box -12 -8 32 272
use FILL  FILL_3__2524_
timestamp 1701859473
transform -1 0 1890 0 -1 9110
box -12 -8 32 272
use FILL  FILL_3__2525_
timestamp 1701859473
transform 1 0 770 0 -1 8590
box -12 -8 32 272
use FILL  FILL_3__2526_
timestamp 1701859473
transform -1 0 1670 0 -1 8590
box -12 -8 32 272
use FILL  FILL_3__2527_
timestamp 1701859473
transform -1 0 1210 0 -1 8590
box -12 -8 32 272
use FILL  FILL_3__2528_
timestamp 1701859473
transform -1 0 990 0 -1 8590
box -12 -8 32 272
use FILL  FILL_3__2529_
timestamp 1701859473
transform -1 0 1230 0 1 9110
box -12 -8 32 272
use FILL  FILL_3__2530_
timestamp 1701859473
transform -1 0 7490 0 -1 6510
box -12 -8 32 272
use FILL  FILL_3__2531_
timestamp 1701859473
transform 1 0 7910 0 1 7550
box -12 -8 32 272
use FILL  FILL_3__2532_
timestamp 1701859473
transform -1 0 9810 0 1 2870
box -12 -8 32 272
use FILL  FILL_3__2533_
timestamp 1701859473
transform -1 0 8890 0 1 4430
box -12 -8 32 272
use FILL  FILL_3__2534_
timestamp 1701859473
transform -1 0 9290 0 -1 5470
box -12 -8 32 272
use FILL  FILL_3__2535_
timestamp 1701859473
transform 1 0 70 0 -1 4950
box -12 -8 32 272
use FILL  FILL_3__2536_
timestamp 1701859473
transform 1 0 630 0 1 4950
box -12 -8 32 272
use FILL  FILL_3__2537_
timestamp 1701859473
transform 1 0 770 0 1 3390
box -12 -8 32 272
use FILL  FILL_3__2538_
timestamp 1701859473
transform -1 0 330 0 -1 3910
box -12 -8 32 272
use FILL  FILL_3__2539_
timestamp 1701859473
transform -1 0 90 0 1 4950
box -12 -8 32 272
use FILL  FILL_3__2540_
timestamp 1701859473
transform 1 0 3030 0 1 2350
box -12 -8 32 272
use FILL  FILL_3__2541_
timestamp 1701859473
transform -1 0 3290 0 1 2870
box -12 -8 32 272
use FILL  FILL_3__2542_
timestamp 1701859473
transform -1 0 2290 0 -1 6510
box -12 -8 32 272
use FILL  FILL_3__2543_
timestamp 1701859473
transform 1 0 850 0 1 4950
box -12 -8 32 272
use FILL  FILL_3__2544_
timestamp 1701859473
transform 1 0 1410 0 1 4430
box -12 -8 32 272
use FILL  FILL_3__2545_
timestamp 1701859473
transform 1 0 1270 0 -1 5470
box -12 -8 32 272
use FILL  FILL_3__2546_
timestamp 1701859473
transform -1 0 2010 0 -1 5470
box -12 -8 32 272
use FILL  FILL_3__2547_
timestamp 1701859473
transform 1 0 1950 0 -1 4430
box -12 -8 32 272
use FILL  FILL_3__2548_
timestamp 1701859473
transform 1 0 1070 0 1 4950
box -12 -8 32 272
use FILL  FILL_3__2549_
timestamp 1701859473
transform 1 0 1290 0 1 4950
box -12 -8 32 272
use FILL  FILL_3__2550_
timestamp 1701859473
transform -1 0 1770 0 -1 5470
box -12 -8 32 272
use FILL  FILL_3__2551_
timestamp 1701859473
transform 1 0 2550 0 -1 9630
box -12 -8 32 272
use FILL  FILL_3__2552_
timestamp 1701859473
transform 1 0 3390 0 -1 5470
box -12 -8 32 272
use FILL  FILL_3__2553_
timestamp 1701859473
transform -1 0 2770 0 -1 6510
box -12 -8 32 272
use FILL  FILL_3__2554_
timestamp 1701859473
transform -1 0 3230 0 1 6510
box -12 -8 32 272
use FILL  FILL_3__2555_
timestamp 1701859473
transform -1 0 3470 0 1 6510
box -12 -8 32 272
use FILL  FILL_3__2556_
timestamp 1701859473
transform -1 0 2790 0 1 6510
box -12 -8 32 272
use FILL  FILL_3__2557_
timestamp 1701859473
transform 1 0 2490 0 -1 6510
box -12 -8 32 272
use FILL  FILL_3__2558_
timestamp 1701859473
transform 1 0 3230 0 -1 7550
box -12 -8 32 272
use FILL  FILL_3__2559_
timestamp 1701859473
transform 1 0 3430 0 -1 7550
box -12 -8 32 272
use FILL  FILL_3__2560_
timestamp 1701859473
transform -1 0 3490 0 1 7030
box -12 -8 32 272
use FILL  FILL_3__2561_
timestamp 1701859473
transform -1 0 1510 0 1 4950
box -12 -8 32 272
use FILL  FILL_3__2562_
timestamp 1701859473
transform 1 0 3230 0 1 7030
box -12 -8 32 272
use FILL  FILL_3__2563_
timestamp 1701859473
transform 1 0 3790 0 1 5470
box -12 -8 32 272
use FILL  FILL_3__2564_
timestamp 1701859473
transform -1 0 3670 0 1 6510
box -12 -8 32 272
use FILL  FILL_3__2565_
timestamp 1701859473
transform 1 0 3730 0 1 7030
box -12 -8 32 272
use FILL  FILL_3__2566_
timestamp 1701859473
transform 1 0 3190 0 1 7550
box -12 -8 32 272
use FILL  FILL_3__2567_
timestamp 1701859473
transform 1 0 3150 0 -1 8070
box -12 -8 32 272
use FILL  FILL_3__2568_
timestamp 1701859473
transform -1 0 2970 0 -1 8590
box -12 -8 32 272
use FILL  FILL_3__2569_
timestamp 1701859473
transform 1 0 2730 0 -1 8590
box -12 -8 32 272
use FILL  FILL_3__2570_
timestamp 1701859473
transform 1 0 2910 0 -1 8070
box -12 -8 32 272
use FILL  FILL_3__2571_
timestamp 1701859473
transform -1 0 3870 0 -1 9630
box -12 -8 32 272
use FILL  FILL_3__2572_
timestamp 1701859473
transform -1 0 3890 0 -1 5990
box -12 -8 32 272
use FILL  FILL_3__2573_
timestamp 1701859473
transform -1 0 3750 0 -1 7030
box -12 -8 32 272
use FILL  FILL_3__2574_
timestamp 1701859473
transform 1 0 3470 0 -1 6510
box -12 -8 32 272
use FILL  FILL_3__2575_
timestamp 1701859473
transform 1 0 3370 0 -1 8070
box -12 -8 32 272
use FILL  FILL_3__2576_
timestamp 1701859473
transform -1 0 3410 0 -1 8590
box -12 -8 32 272
use FILL  FILL_3__2577_
timestamp 1701859473
transform 1 0 3290 0 1 9110
box -12 -8 32 272
use FILL  FILL_3__2578_
timestamp 1701859473
transform 1 0 3790 0 1 9110
box -12 -8 32 272
use FILL  FILL_3__2579_
timestamp 1701859473
transform -1 0 2770 0 -1 9630
box -12 -8 32 272
use FILL  FILL_3__2580_
timestamp 1701859473
transform -1 0 4130 0 -1 9110
box -12 -8 32 272
use FILL  FILL_3__2581_
timestamp 1701859473
transform -1 0 4050 0 1 9110
box -12 -8 32 272
use FILL  FILL_3__2582_
timestamp 1701859473
transform 1 0 3550 0 1 9110
box -12 -8 32 272
use FILL  FILL_3__2583_
timestamp 1701859473
transform 1 0 3050 0 1 9110
box -12 -8 32 272
use FILL  FILL_3__2584_
timestamp 1701859473
transform 1 0 2810 0 1 9110
box -12 -8 32 272
use FILL  FILL_3__2585_
timestamp 1701859473
transform 1 0 3910 0 -1 9110
box -12 -8 32 272
use FILL  FILL_3__2586_
timestamp 1701859473
transform 1 0 3070 0 1 9630
box -12 -8 32 272
use FILL  FILL_3__2587_
timestamp 1701859473
transform 1 0 3650 0 -1 9110
box -12 -8 32 272
use FILL  FILL_3__2588_
timestamp 1701859473
transform 1 0 3250 0 1 8590
box -12 -8 32 272
use FILL  FILL_3__2589_
timestamp 1701859473
transform 1 0 3090 0 -1 10150
box -12 -8 32 272
use FILL  FILL_3__2590_
timestamp 1701859473
transform 1 0 2830 0 -1 10150
box -12 -8 32 272
use FILL  FILL_3__2591_
timestamp 1701859473
transform -1 0 3590 0 -1 11190
box -12 -8 32 272
use FILL  FILL_3__2592_
timestamp 1701859473
transform -1 0 3650 0 -1 9630
box -12 -8 32 272
use FILL  FILL_3__2593_
timestamp 1701859473
transform -1 0 3170 0 -1 9630
box -12 -8 32 272
use FILL  FILL_3__2594_
timestamp 1701859473
transform -1 0 3330 0 -1 10150
box -12 -8 32 272
use FILL  FILL_3__2595_
timestamp 1701859473
transform 1 0 3050 0 -1 11190
box -12 -8 32 272
use FILL  FILL_3__2596_
timestamp 1701859473
transform 1 0 3330 0 -1 11190
box -12 -8 32 272
use FILL  FILL_3__2597_
timestamp 1701859473
transform 1 0 2790 0 -1 10670
box -12 -8 32 272
use FILL  FILL_3__2598_
timestamp 1701859473
transform -1 0 3530 0 1 9630
box -12 -8 32 272
use FILL  FILL_3__2599_
timestamp 1701859473
transform -1 0 3310 0 1 9630
box -12 -8 32 272
use FILL  FILL_3__2600_
timestamp 1701859473
transform -1 0 3030 0 1 10150
box -12 -8 32 272
use FILL  FILL_3__2601_
timestamp 1701859473
transform 1 0 2990 0 -1 10670
box -12 -8 32 272
use FILL  FILL_3__2602_
timestamp 1701859473
transform -1 0 3250 0 -1 10670
box -12 -8 32 272
use FILL  FILL_3__2603_
timestamp 1701859473
transform 1 0 3450 0 -1 10670
box -12 -8 32 272
use FILL  FILL_3__2604_
timestamp 1701859473
transform 1 0 3250 0 1 10150
box -12 -8 32 272
use FILL  FILL_3__2605_
timestamp 1701859473
transform 1 0 2370 0 1 10670
box -12 -8 32 272
use FILL  FILL_3__2606_
timestamp 1701859473
transform 1 0 2570 0 1 10670
box -12 -8 32 272
use FILL  FILL_3__2607_
timestamp 1701859473
transform -1 0 2810 0 1 10670
box -12 -8 32 272
use FILL  FILL_3__2608_
timestamp 1701859473
transform -1 0 3770 0 1 9630
box -12 -8 32 272
use FILL  FILL_3__2609_
timestamp 1701859473
transform -1 0 2390 0 1 9630
box -12 -8 32 272
use FILL  FILL_3__2610_
timestamp 1701859473
transform -1 0 2610 0 -1 10150
box -12 -8 32 272
use FILL  FILL_3__2611_
timestamp 1701859473
transform -1 0 2330 0 -1 10670
box -12 -8 32 272
use FILL  FILL_3__2612_
timestamp 1701859473
transform 1 0 2550 0 -1 10670
box -12 -8 32 272
use FILL  FILL_3__2613_
timestamp 1701859473
transform 1 0 1870 0 1 10670
box -12 -8 32 272
use FILL  FILL_3__2614_
timestamp 1701859473
transform 1 0 1870 0 -1 10670
box -12 -8 32 272
use FILL  FILL_3__2615_
timestamp 1701859473
transform -1 0 2390 0 -1 11190
box -12 -8 32 272
use FILL  FILL_3__2616_
timestamp 1701859473
transform -1 0 3410 0 -1 9630
box -12 -8 32 272
use FILL  FILL_3__2617_
timestamp 1701859473
transform 1 0 2310 0 -1 9630
box -12 -8 32 272
use FILL  FILL_3__2618_
timestamp 1701859473
transform -1 0 2590 0 1 10150
box -12 -8 32 272
use FILL  FILL_3__2619_
timestamp 1701859473
transform 1 0 2090 0 1 10670
box -12 -8 32 272
use FILL  FILL_3__2620_
timestamp 1701859473
transform 1 0 2130 0 -1 11190
box -12 -8 32 272
use FILL  FILL_3__2621_
timestamp 1701859473
transform -1 0 1410 0 1 5470
box -12 -8 32 272
use FILL  FILL_3__2622_
timestamp 1701859473
transform -1 0 1250 0 -1 5990
box -12 -8 32 272
use FILL  FILL_3__2623_
timestamp 1701859473
transform 1 0 2470 0 -1 5470
box -12 -8 32 272
use FILL  FILL_3__2624_
timestamp 1701859473
transform -1 0 2430 0 1 5470
box -12 -8 32 272
use FILL  FILL_3__2625_
timestamp 1701859473
transform 1 0 2230 0 -1 5470
box -12 -8 32 272
use FILL  FILL_3__2626_
timestamp 1701859473
transform -1 0 970 0 -1 5470
box -12 -8 32 272
use FILL  FILL_3__2627_
timestamp 1701859473
transform -1 0 1490 0 1 3910
box -12 -8 32 272
use FILL  FILL_3__2628_
timestamp 1701859473
transform 1 0 1170 0 1 3910
box -12 -8 32 272
use FILL  FILL_3__2629_
timestamp 1701859473
transform -1 0 770 0 -1 5470
box -12 -8 32 272
use FILL  FILL_3__2630_
timestamp 1701859473
transform 1 0 750 0 -1 5990
box -12 -8 32 272
use FILL  FILL_3__2631_
timestamp 1701859473
transform -1 0 750 0 1 5990
box -12 -8 32 272
use FILL  FILL_3__2632_
timestamp 1701859473
transform 1 0 2130 0 1 10150
box -12 -8 32 272
use FILL  FILL_3__2633_
timestamp 1701859473
transform -1 0 2370 0 1 10150
box -12 -8 32 272
use FILL  FILL_3__2634_
timestamp 1701859473
transform 1 0 2330 0 -1 10150
box -12 -8 32 272
use FILL  FILL_3__2635_
timestamp 1701859473
transform 1 0 2110 0 -1 10150
box -12 -8 32 272
use FILL  FILL_3__2636_
timestamp 1701859473
transform -1 0 750 0 -1 10150
box -12 -8 32 272
use FILL  FILL_3__2637_
timestamp 1701859473
transform -1 0 550 0 1 6510
box -12 -8 32 272
use FILL  FILL_3__2638_
timestamp 1701859473
transform -1 0 330 0 1 6510
box -12 -8 32 272
use FILL  FILL_3__2639_
timestamp 1701859473
transform -1 0 310 0 -1 6510
box -12 -8 32 272
use FILL  FILL_3__2640_
timestamp 1701859473
transform -1 0 310 0 1 5990
box -12 -8 32 272
use FILL  FILL_3__2641_
timestamp 1701859473
transform 1 0 70 0 -1 7550
box -12 -8 32 272
use FILL  FILL_3__2642_
timestamp 1701859473
transform -1 0 410 0 1 4950
box -12 -8 32 272
use FILL  FILL_3__2643_
timestamp 1701859473
transform -1 0 2550 0 1 6510
box -12 -8 32 272
use FILL  FILL_3__2644_
timestamp 1701859473
transform 1 0 2590 0 -1 7030
box -12 -8 32 272
use FILL  FILL_3__2645_
timestamp 1701859473
transform 1 0 2770 0 1 7030
box -12 -8 32 272
use FILL  FILL_3__2646_
timestamp 1701859473
transform 1 0 2070 0 1 7030
box -12 -8 32 272
use FILL  FILL_3__2647_
timestamp 1701859473
transform 1 0 750 0 1 7550
box -12 -8 32 272
use FILL  FILL_3__2648_
timestamp 1701859473
transform 1 0 290 0 1 7550
box -12 -8 32 272
use FILL  FILL_3__2649_
timestamp 1701859473
transform 1 0 270 0 -1 7550
box -12 -8 32 272
use FILL  FILL_3__2650_
timestamp 1701859473
transform -1 0 750 0 -1 7550
box -12 -8 32 272
use FILL  FILL_3__2651_
timestamp 1701859473
transform 1 0 490 0 -1 7550
box -12 -8 32 272
use FILL  FILL_3__2652_
timestamp 1701859473
transform 1 0 490 0 1 7030
box -12 -8 32 272
use FILL  FILL_3__2653_
timestamp 1701859473
transform 1 0 70 0 1 7550
box -12 -8 32 272
use FILL  FILL_3__2654_
timestamp 1701859473
transform -1 0 550 0 1 7550
box -12 -8 32 272
use FILL  FILL_3__2655_
timestamp 1701859473
transform 1 0 1870 0 1 7030
box -12 -8 32 272
use FILL  FILL_3__2656_
timestamp 1701859473
transform 1 0 1510 0 -1 5470
box -12 -8 32 272
use FILL  FILL_3__2657_
timestamp 1701859473
transform -1 0 1710 0 1 5990
box -12 -8 32 272
use FILL  FILL_3__2658_
timestamp 1701859473
transform -1 0 2190 0 1 5470
box -12 -8 32 272
use FILL  FILL_3__2659_
timestamp 1701859473
transform 1 0 1950 0 -1 5990
box -12 -8 32 272
use FILL  FILL_3__2660_
timestamp 1701859473
transform -1 0 1950 0 1 5470
box -12 -8 32 272
use FILL  FILL_3__2661_
timestamp 1701859473
transform -1 0 1630 0 1 5470
box -12 -8 32 272
use FILL  FILL_3__2662_
timestamp 1701859473
transform 1 0 730 0 1 5470
box -12 -8 32 272
use FILL  FILL_3__2663_
timestamp 1701859473
transform -1 0 1010 0 -1 5990
box -12 -8 32 272
use FILL  FILL_3__2664_
timestamp 1701859473
transform 1 0 730 0 -1 7030
box -12 -8 32 272
use FILL  FILL_3__2665_
timestamp 1701859473
transform 1 0 1190 0 -1 7030
box -12 -8 32 272
use FILL  FILL_3__2666_
timestamp 1701859473
transform 1 0 1390 0 1 7030
box -12 -8 32 272
use FILL  FILL_3__2667_
timestamp 1701859473
transform 1 0 930 0 -1 7030
box -12 -8 32 272
use FILL  FILL_3__2668_
timestamp 1701859473
transform -1 0 2730 0 1 7550
box -12 -8 32 272
use FILL  FILL_3__2669_
timestamp 1701859473
transform 1 0 2670 0 -1 8070
box -12 -8 32 272
use FILL  FILL_3__2670_
timestamp 1701859473
transform 1 0 1930 0 -1 8070
box -12 -8 32 272
use FILL  FILL_3__2671_
timestamp 1701859473
transform -1 0 1430 0 1 7550
box -12 -8 32 272
use FILL  FILL_3__2672_
timestamp 1701859473
transform 1 0 1150 0 -1 7550
box -12 -8 32 272
use FILL  FILL_3__2673_
timestamp 1701859473
transform -1 0 1350 0 -1 7550
box -12 -8 32 272
use FILL  FILL_3__2674_
timestamp 1701859473
transform 1 0 1630 0 1 7030
box -12 -8 32 272
use FILL  FILL_3__2675_
timestamp 1701859473
transform 1 0 1570 0 -1 7550
box -12 -8 32 272
use FILL  FILL_3__2676_
timestamp 1701859473
transform -1 0 2010 0 -1 7550
box -12 -8 32 272
use FILL  FILL_3__2677_
timestamp 1701859473
transform 1 0 2410 0 -1 8070
box -12 -8 32 272
use FILL  FILL_3__2678_
timestamp 1701859473
transform -1 0 2190 0 -1 8070
box -12 -8 32 272
use FILL  FILL_3__2679_
timestamp 1701859473
transform -1 0 1630 0 1 8070
box -12 -8 32 272
use FILL  FILL_3__2680_
timestamp 1701859473
transform -1 0 310 0 -1 8590
box -12 -8 32 272
use FILL  FILL_3__2681_
timestamp 1701859473
transform 1 0 930 0 -1 7550
box -12 -8 32 272
use FILL  FILL_3__2682_
timestamp 1701859473
transform -1 0 310 0 -1 8070
box -12 -8 32 272
use FILL  FILL_3__2683_
timestamp 1701859473
transform -1 0 90 0 -1 9630
box -12 -8 32 272
use FILL  FILL_3__2684_
timestamp 1701859473
transform -1 0 90 0 1 10150
box -12 -8 32 272
use FILL  FILL_3__2685_
timestamp 1701859473
transform 1 0 970 0 1 5990
box -12 -8 32 272
use FILL  FILL_3__2686_
timestamp 1701859473
transform 1 0 950 0 1 7550
box -12 -8 32 272
use FILL  FILL_3__2687_
timestamp 1701859473
transform -1 0 950 0 -1 10150
box -12 -8 32 272
use FILL  FILL_3__2688_
timestamp 1701859473
transform 1 0 70 0 -1 10150
box -12 -8 32 272
use FILL  FILL_3__2689_
timestamp 1701859473
transform 1 0 290 0 -1 9630
box -12 -8 32 272
use FILL  FILL_3__2690_
timestamp 1701859473
transform 1 0 290 0 1 9110
box -12 -8 32 272
use FILL  FILL_3__2691_
timestamp 1701859473
transform 1 0 2750 0 1 8590
box -12 -8 32 272
use FILL  FILL_3__2692_
timestamp 1701859473
transform 1 0 2510 0 1 8590
box -12 -8 32 272
use FILL  FILL_3__2693_
timestamp 1701859473
transform -1 0 1170 0 -1 9630
box -12 -8 32 272
use FILL  FILL_3__2694_
timestamp 1701859473
transform 1 0 750 0 -1 9630
box -12 -8 32 272
use FILL  FILL_3__2695_
timestamp 1701859473
transform 1 0 70 0 1 9630
box -12 -8 32 272
use FILL  FILL_3__2696_
timestamp 1701859473
transform -1 0 550 0 -1 10150
box -12 -8 32 272
use FILL  FILL_3__2697_
timestamp 1701859473
transform 1 0 290 0 -1 10150
box -12 -8 32 272
use FILL  FILL_3__2698_
timestamp 1701859473
transform 1 0 310 0 1 9630
box -12 -8 32 272
use FILL  FILL_3__2699_
timestamp 1701859473
transform 1 0 530 0 -1 9630
box -12 -8 32 272
use FILL  FILL_3__2700_
timestamp 1701859473
transform 1 0 550 0 1 9630
box -12 -8 32 272
use FILL  FILL_3__2701_
timestamp 1701859473
transform -1 0 770 0 -1 10670
box -12 -8 32 272
use FILL  FILL_3__2702_
timestamp 1701859473
transform 1 0 3490 0 1 8590
box -12 -8 32 272
use FILL  FILL_3__2703_
timestamp 1701859473
transform -1 0 3030 0 1 8590
box -12 -8 32 272
use FILL  FILL_3__2704_
timestamp 1701859473
transform -1 0 1510 0 1 9630
box -12 -8 32 272
use FILL  FILL_3__2705_
timestamp 1701859473
transform 1 0 1250 0 1 9630
box -12 -8 32 272
use FILL  FILL_3__2706_
timestamp 1701859473
transform 1 0 270 0 1 10150
box -12 -8 32 272
use FILL  FILL_3__2707_
timestamp 1701859473
transform -1 0 510 0 1 10150
box -12 -8 32 272
use FILL  FILL_3__2708_
timestamp 1701859473
transform 1 0 710 0 1 10150
box -12 -8 32 272
use FILL  FILL_3__2709_
timestamp 1701859473
transform -1 0 530 0 -1 10670
box -12 -8 32 272
use FILL  FILL_3__2710_
timestamp 1701859473
transform 1 0 1710 0 1 10150
box -12 -8 32 272
use FILL  FILL_3__2711_
timestamp 1701859473
transform 1 0 2250 0 1 8590
box -12 -8 32 272
use FILL  FILL_3__2712_
timestamp 1701859473
transform -1 0 2030 0 1 8590
box -12 -8 32 272
use FILL  FILL_3__2713_
timestamp 1701859473
transform -1 0 1890 0 -1 9630
box -12 -8 32 272
use FILL  FILL_3__2714_
timestamp 1701859473
transform 1 0 1650 0 -1 10150
box -12 -8 32 272
use FILL  FILL_3__2715_
timestamp 1701859473
transform 1 0 970 0 1 10150
box -12 -8 32 272
use FILL  FILL_3__2716_
timestamp 1701859473
transform 1 0 1210 0 1 10150
box -12 -8 32 272
use FILL  FILL_3__2717_
timestamp 1701859473
transform 1 0 1470 0 1 10150
box -12 -8 32 272
use FILL  FILL_3__2718_
timestamp 1701859473
transform -1 0 10050 0 1 4950
box -12 -8 32 272
use FILL  FILL_3__2719_
timestamp 1701859473
transform -1 0 9810 0 1 4950
box -12 -8 32 272
use FILL  FILL_3__2720_
timestamp 1701859473
transform -1 0 4590 0 1 4950
box -12 -8 32 272
use FILL  FILL_3__2721_
timestamp 1701859473
transform -1 0 7350 0 -1 2350
box -12 -8 32 272
use FILL  FILL_3__2722_
timestamp 1701859473
transform 1 0 9990 0 -1 790
box -12 -8 32 272
use FILL  FILL_3__2723_
timestamp 1701859473
transform -1 0 7110 0 1 1830
box -12 -8 32 272
use FILL  FILL_3__2724_
timestamp 1701859473
transform -1 0 7110 0 -1 2350
box -12 -8 32 272
use FILL  FILL_3__2725_
timestamp 1701859473
transform 1 0 6970 0 1 3390
box -12 -8 32 272
use FILL  FILL_3__2726_
timestamp 1701859473
transform -1 0 7210 0 1 3390
box -12 -8 32 272
use FILL  FILL_3__2727_
timestamp 1701859473
transform -1 0 5430 0 1 3390
box -12 -8 32 272
use FILL  FILL_3__2728_
timestamp 1701859473
transform -1 0 5650 0 1 3390
box -12 -8 32 272
use FILL  FILL_3__2729_
timestamp 1701859473
transform -1 0 6750 0 -1 3910
box -12 -8 32 272
use FILL  FILL_3__2730_
timestamp 1701859473
transform 1 0 8250 0 -1 3910
box -12 -8 32 272
use FILL  FILL_3__2731_
timestamp 1701859473
transform 1 0 9270 0 1 1830
box -12 -8 32 272
use FILL  FILL_3__2732_
timestamp 1701859473
transform 1 0 7710 0 1 1830
box -12 -8 32 272
use FILL  FILL_3__2733_
timestamp 1701859473
transform 1 0 8590 0 1 2350
box -12 -8 32 272
use FILL  FILL_3__2734_
timestamp 1701859473
transform 1 0 7170 0 -1 5470
box -12 -8 32 272
use FILL  FILL_3__2735_
timestamp 1701859473
transform 1 0 7250 0 -1 2870
box -12 -8 32 272
use FILL  FILL_3__2736_
timestamp 1701859473
transform -1 0 7530 0 1 1310
box -12 -8 32 272
use FILL  FILL_3__2737_
timestamp 1701859473
transform 1 0 8590 0 1 1830
box -12 -8 32 272
use FILL  FILL_3__2738_
timestamp 1701859473
transform -1 0 7970 0 -1 2870
box -12 -8 32 272
use FILL  FILL_3__2739_
timestamp 1701859473
transform -1 0 7790 0 1 2870
box -12 -8 32 272
use FILL  FILL_3__2740_
timestamp 1701859473
transform -1 0 6570 0 -1 1830
box -12 -8 32 272
use FILL  FILL_3__2741_
timestamp 1701859473
transform 1 0 6770 0 -1 1830
box -12 -8 32 272
use FILL  FILL_3__2742_
timestamp 1701859473
transform -1 0 8210 0 -1 2870
box -12 -8 32 272
use FILL  FILL_3__2743_
timestamp 1701859473
transform -1 0 8230 0 1 2870
box -12 -8 32 272
use FILL  FILL_3__2744_
timestamp 1701859473
transform -1 0 7350 0 -1 270
box -12 -8 32 272
use FILL  FILL_3__2745_
timestamp 1701859473
transform -1 0 7310 0 1 1830
box -12 -8 32 272
use FILL  FILL_3__2746_
timestamp 1701859473
transform 1 0 7970 0 1 2870
box -12 -8 32 272
use FILL  FILL_3__2747_
timestamp 1701859473
transform -1 0 7770 0 -1 2350
box -12 -8 32 272
use FILL  FILL_3__2748_
timestamp 1701859473
transform 1 0 7950 0 -1 2350
box -12 -8 32 272
use FILL  FILL_3__2749_
timestamp 1701859473
transform 1 0 5910 0 1 1830
box -12 -8 32 272
use FILL  FILL_3__2750_
timestamp 1701859473
transform -1 0 6670 0 -1 1310
box -12 -8 32 272
use FILL  FILL_3__2751_
timestamp 1701859473
transform -1 0 6390 0 1 1830
box -12 -8 32 272
use FILL  FILL_3__2752_
timestamp 1701859473
transform -1 0 7750 0 1 2350
box -12 -8 32 272
use FILL  FILL_3__2753_
timestamp 1701859473
transform -1 0 7490 0 1 2350
box -12 -8 32 272
use FILL  FILL_3__2754_
timestamp 1701859473
transform 1 0 8830 0 -1 4950
box -12 -8 32 272
use FILL  FILL_3__2755_
timestamp 1701859473
transform 1 0 9730 0 1 790
box -12 -8 32 272
use FILL  FILL_3__2756_
timestamp 1701859473
transform -1 0 9970 0 1 790
box -12 -8 32 272
use FILL  FILL_3__2757_
timestamp 1701859473
transform 1 0 10670 0 -1 2870
box -12 -8 32 272
use FILL  FILL_3__2758_
timestamp 1701859473
transform -1 0 9170 0 -1 2870
box -12 -8 32 272
use FILL  FILL_3__2759_
timestamp 1701859473
transform 1 0 9090 0 1 4430
box -12 -8 32 272
use FILL  FILL_3__2760_
timestamp 1701859473
transform 1 0 10430 0 -1 790
box -12 -8 32 272
use FILL  FILL_3__2761_
timestamp 1701859473
transform 1 0 10190 0 -1 790
box -12 -8 32 272
use FILL  FILL_3__2762_
timestamp 1701859473
transform -1 0 10870 0 -1 1830
box -12 -8 32 272
use FILL  FILL_3__2763_
timestamp 1701859473
transform 1 0 6610 0 1 1830
box -12 -8 32 272
use FILL  FILL_3__2764_
timestamp 1701859473
transform -1 0 6870 0 1 1830
box -12 -8 32 272
use FILL  FILL_3__2765_
timestamp 1701859473
transform -1 0 10170 0 1 1830
box -12 -8 32 272
use FILL  FILL_3__2766_
timestamp 1701859473
transform -1 0 9990 0 -1 1830
box -12 -8 32 272
use FILL  FILL_3__2767_
timestamp 1701859473
transform -1 0 10410 0 -1 1830
box -12 -8 32 272
use FILL  FILL_3__2768_
timestamp 1701859473
transform -1 0 10390 0 1 1830
box -12 -8 32 272
use FILL  FILL_3__2769_
timestamp 1701859473
transform -1 0 10850 0 1 2350
box -12 -8 32 272
use FILL  FILL_3__2770_
timestamp 1701859473
transform -1 0 10630 0 -1 1830
box -12 -8 32 272
use FILL  FILL_3__2771_
timestamp 1701859473
transform 1 0 11050 0 1 2350
box -12 -8 32 272
use FILL  FILL_3__2772_
timestamp 1701859473
transform -1 0 10710 0 1 4950
box -12 -8 32 272
use FILL  FILL_3__2773_
timestamp 1701859473
transform 1 0 10450 0 -1 3910
box -12 -8 32 272
use FILL  FILL_3__2774_
timestamp 1701859473
transform -1 0 10750 0 -1 2350
box -12 -8 32 272
use FILL  FILL_3__2775_
timestamp 1701859473
transform -1 0 9110 0 -1 1310
box -12 -8 32 272
use FILL  FILL_3__2776_
timestamp 1701859473
transform 1 0 10650 0 -1 790
box -12 -8 32 272
use FILL  FILL_3__2777_
timestamp 1701859473
transform -1 0 8410 0 -1 270
box -12 -8 32 272
use FILL  FILL_3__2778_
timestamp 1701859473
transform 1 0 10950 0 1 270
box -12 -8 32 272
use FILL  FILL_3__2779_
timestamp 1701859473
transform 1 0 9030 0 -1 1830
box -12 -8 32 272
use FILL  FILL_3__2780_
timestamp 1701859473
transform -1 0 10050 0 1 1310
box -12 -8 32 272
use FILL  FILL_3__2781_
timestamp 1701859473
transform 1 0 10190 0 -1 1310
box -12 -8 32 272
use FILL  FILL_3__2782_
timestamp 1701859473
transform 1 0 8810 0 1 1830
box -12 -8 32 272
use FILL  FILL_3__2783_
timestamp 1701859473
transform 1 0 8370 0 -1 1310
box -12 -8 32 272
use FILL  FILL_3__2784_
timestamp 1701859473
transform 1 0 8610 0 -1 1310
box -12 -8 32 272
use FILL  FILL_3__2785_
timestamp 1701859473
transform 1 0 8830 0 -1 1830
box -12 -8 32 272
use FILL  FILL_3__2786_
timestamp 1701859473
transform -1 0 9310 0 -1 1310
box -12 -8 32 272
use FILL  FILL_3__2787_
timestamp 1701859473
transform -1 0 9510 0 -1 1830
box -12 -8 32 272
use FILL  FILL_3__2788_
timestamp 1701859473
transform 1 0 10190 0 -1 1830
box -12 -8 32 272
use FILL  FILL_3__2789_
timestamp 1701859473
transform 1 0 10270 0 1 1310
box -12 -8 32 272
use FILL  FILL_3__2790_
timestamp 1701859473
transform -1 0 10070 0 -1 2350
box -12 -8 32 272
use FILL  FILL_3__2791_
timestamp 1701859473
transform 1 0 9830 0 -1 2350
box -12 -8 32 272
use FILL  FILL_3__2792_
timestamp 1701859473
transform -1 0 10290 0 -1 2350
box -12 -8 32 272
use FILL  FILL_3__2793_
timestamp 1701859473
transform -1 0 10530 0 -1 2350
box -12 -8 32 272
use FILL  FILL_3__2794_
timestamp 1701859473
transform -1 0 10950 0 -1 2350
box -12 -8 32 272
use FILL  FILL_3__2795_
timestamp 1701859473
transform -1 0 10910 0 -1 2870
box -12 -8 32 272
use FILL  FILL_3__2796_
timestamp 1701859473
transform -1 0 10250 0 -1 2870
box -12 -8 32 272
use FILL  FILL_3__2797_
timestamp 1701859473
transform -1 0 9750 0 -1 1830
box -12 -8 32 272
use FILL  FILL_3__2798_
timestamp 1701859473
transform -1 0 10630 0 1 2350
box -12 -8 32 272
use FILL  FILL_3__2799_
timestamp 1701859473
transform 1 0 10410 0 -1 2870
box -12 -8 32 272
use FILL  FILL_3__2800_
timestamp 1701859473
transform -1 0 10430 0 -1 4430
box -12 -8 32 272
use FILL  FILL_3__2801_
timestamp 1701859473
transform -1 0 9390 0 -1 2870
box -12 -8 32 272
use FILL  FILL_3__2802_
timestamp 1701859473
transform -1 0 7250 0 -1 1830
box -12 -8 32 272
use FILL  FILL_3__2803_
timestamp 1701859473
transform 1 0 8450 0 -1 2870
box -12 -8 32 272
use FILL  FILL_3__2804_
timestamp 1701859473
transform -1 0 9510 0 -1 3390
box -12 -8 32 272
use FILL  FILL_3__2805_
timestamp 1701859473
transform -1 0 9810 0 -1 2870
box -12 -8 32 272
use FILL  FILL_3__2806_
timestamp 1701859473
transform 1 0 9570 0 -1 2870
box -12 -8 32 272
use FILL  FILL_3__2807_
timestamp 1701859473
transform 1 0 8910 0 -1 2350
box -12 -8 32 272
use FILL  FILL_3__2808_
timestamp 1701859473
transform 1 0 8670 0 -1 2350
box -12 -8 32 272
use FILL  FILL_3__2809_
timestamp 1701859473
transform 1 0 10390 0 1 2350
box -12 -8 32 272
use FILL  FILL_3__2810_
timestamp 1701859473
transform -1 0 10170 0 1 2350
box -12 -8 32 272
use FILL  FILL_3__2811_
timestamp 1701859473
transform 1 0 4950 0 -1 4430
box -12 -8 32 272
use FILL  FILL_3__2812_
timestamp 1701859473
transform -1 0 8910 0 1 4950
box -12 -8 32 272
use FILL  FILL_3__2813_
timestamp 1701859473
transform 1 0 9010 0 1 3390
box -12 -8 32 272
use FILL  FILL_3__2814_
timestamp 1701859473
transform -1 0 8830 0 -1 4430
box -12 -8 32 272
use FILL  FILL_3__2815_
timestamp 1701859473
transform -1 0 8610 0 1 3910
box -12 -8 32 272
use FILL  FILL_3__2816_
timestamp 1701859473
transform -1 0 8230 0 1 4950
box -12 -8 32 272
use FILL  FILL_3__2817_
timestamp 1701859473
transform 1 0 8670 0 1 4950
box -12 -8 32 272
use FILL  FILL_3__2818_
timestamp 1701859473
transform 1 0 8370 0 -1 4430
box -12 -8 32 272
use FILL  FILL_3__2819_
timestamp 1701859473
transform 1 0 8570 0 -1 4430
box -12 -8 32 272
use FILL  FILL_3__2820_
timestamp 1701859473
transform -1 0 9530 0 1 2350
box -12 -8 32 272
use FILL  FILL_3__2821_
timestamp 1701859473
transform 1 0 9050 0 1 2350
box -12 -8 32 272
use FILL  FILL_3__2822_
timestamp 1701859473
transform -1 0 9050 0 1 1830
box -12 -8 32 272
use FILL  FILL_3__2823_
timestamp 1701859473
transform -1 0 8830 0 1 2350
box -12 -8 32 272
use FILL  FILL_3__2824_
timestamp 1701859473
transform 1 0 9950 0 -1 3390
box -12 -8 32 272
use FILL  FILL_3__2825_
timestamp 1701859473
transform -1 0 10670 0 -1 3390
box -12 -8 32 272
use FILL  FILL_3__2826_
timestamp 1701859473
transform 1 0 9530 0 1 790
box -12 -8 32 272
use FILL  FILL_3__2827_
timestamp 1701859473
transform -1 0 9270 0 -1 1830
box -12 -8 32 272
use FILL  FILL_3__2828_
timestamp 1701859473
transform 1 0 6990 0 -1 1830
box -12 -8 32 272
use FILL  FILL_3__2829_
timestamp 1701859473
transform -1 0 10010 0 1 2870
box -12 -8 32 272
use FILL  FILL_3__2830_
timestamp 1701859473
transform 1 0 8310 0 -1 3390
box -12 -8 32 272
use FILL  FILL_3__2831_
timestamp 1701859473
transform 1 0 8350 0 1 3910
box -12 -8 32 272
use FILL  FILL_3__2832_
timestamp 1701859473
transform -1 0 9330 0 1 2350
box -12 -8 32 272
use FILL  FILL_3__2833_
timestamp 1701859473
transform -1 0 9270 0 -1 3390
box -12 -8 32 272
use FILL  FILL_3__2834_
timestamp 1701859473
transform -1 0 9030 0 -1 3390
box -12 -8 32 272
use FILL  FILL_3__2835_
timestamp 1701859473
transform -1 0 9330 0 1 790
box -12 -8 32 272
use FILL  FILL_3__2836_
timestamp 1701859473
transform 1 0 8910 0 1 1310
box -12 -8 32 272
use FILL  FILL_3__2837_
timestamp 1701859473
transform -1 0 9590 0 1 1310
box -12 -8 32 272
use FILL  FILL_3__2838_
timestamp 1701859473
transform -1 0 9710 0 1 3390
box -12 -8 32 272
use FILL  FILL_3__2839_
timestamp 1701859473
transform -1 0 9750 0 -1 3390
box -12 -8 32 272
use FILL  FILL_3__2840_
timestamp 1701859473
transform 1 0 9070 0 -1 270
box -12 -8 32 272
use FILL  FILL_3__2841_
timestamp 1701859473
transform -1 0 8870 0 -1 270
box -12 -8 32 272
use FILL  FILL_3__2842_
timestamp 1701859473
transform 1 0 9290 0 -1 270
box -12 -8 32 272
use FILL  FILL_3__2843_
timestamp 1701859473
transform 1 0 9530 0 -1 270
box -12 -8 32 272
use FILL  FILL_3__2844_
timestamp 1701859473
transform 1 0 9330 0 1 270
box -12 -8 32 272
use FILL  FILL_3__2845_
timestamp 1701859473
transform -1 0 10010 0 1 270
box -12 -8 32 272
use FILL  FILL_3__2846_
timestamp 1701859473
transform 1 0 9750 0 1 270
box -12 -8 32 272
use FILL  FILL_3__2847_
timestamp 1701859473
transform -1 0 11150 0 -1 10670
box -12 -8 32 272
use FILL  FILL_3__2848_
timestamp 1701859473
transform -1 0 10630 0 -1 1310
box -12 -8 32 272
use FILL  FILL_3__2849_
timestamp 1701859473
transform -1 0 10970 0 1 1310
box -12 -8 32 272
use FILL  FILL_3__2850_
timestamp 1701859473
transform -1 0 11110 0 -1 1830
box -12 -8 32 272
use FILL  FILL_3__2851_
timestamp 1701859473
transform 1 0 10710 0 -1 3910
box -12 -8 32 272
use FILL  FILL_3__2852_
timestamp 1701859473
transform -1 0 8910 0 1 270
box -12 -8 32 272
use FILL  FILL_3__2853_
timestamp 1701859473
transform -1 0 9130 0 1 270
box -12 -8 32 272
use FILL  FILL_3__2854_
timestamp 1701859473
transform 1 0 10630 0 1 790
box -12 -8 32 272
use FILL  FILL_3__2855_
timestamp 1701859473
transform -1 0 9830 0 1 1310
box -12 -8 32 272
use FILL  FILL_3__2856_
timestamp 1701859473
transform -1 0 10490 0 1 1310
box -12 -8 32 272
use FILL  FILL_3__2857_
timestamp 1701859473
transform -1 0 10730 0 1 1310
box -12 -8 32 272
use FILL  FILL_3__2858_
timestamp 1701859473
transform -1 0 11090 0 1 1830
box -12 -8 32 272
use FILL  FILL_3__2859_
timestamp 1701859473
transform 1 0 10950 0 -1 3910
box -12 -8 32 272
use FILL  FILL_3__2860_
timestamp 1701859473
transform 1 0 10870 0 -1 3390
box -12 -8 32 272
use FILL  FILL_3__2861_
timestamp 1701859473
transform 1 0 9750 0 -1 270
box -12 -8 32 272
use FILL  FILL_3__2862_
timestamp 1701859473
transform 1 0 8610 0 -1 270
box -12 -8 32 272
use FILL  FILL_3__2863_
timestamp 1701859473
transform -1 0 10250 0 1 270
box -12 -8 32 272
use FILL  FILL_3__2864_
timestamp 1701859473
transform 1 0 10490 0 1 270
box -12 -8 32 272
use FILL  FILL_3__2865_
timestamp 1701859473
transform -1 0 10730 0 1 270
box -12 -8 32 272
use FILL  FILL_3__2866_
timestamp 1701859473
transform -1 0 11110 0 -1 790
box -12 -8 32 272
use FILL  FILL_3__2867_
timestamp 1701859473
transform 1 0 11070 0 -1 3390
box -12 -8 32 272
use FILL  FILL_3__2868_
timestamp 1701859473
transform 1 0 11050 0 1 790
box -12 -8 32 272
use FILL  FILL_3__2869_
timestamp 1701859473
transform 1 0 10170 0 1 790
box -12 -8 32 272
use FILL  FILL_3__2870_
timestamp 1701859473
transform -1 0 10390 0 1 790
box -12 -8 32 272
use FILL  FILL_3__2871_
timestamp 1701859473
transform -1 0 10830 0 1 790
box -12 -8 32 272
use FILL  FILL_3__2872_
timestamp 1701859473
transform -1 0 11170 0 1 1310
box -12 -8 32 272
use FILL  FILL_3__2873_
timestamp 1701859473
transform -1 0 9950 0 1 3390
box -12 -8 32 272
use FILL  FILL_3__2874_
timestamp 1701859473
transform -1 0 10190 0 1 3390
box -12 -8 32 272
use FILL  FILL_3__2875_
timestamp 1701859473
transform -1 0 10770 0 -1 4950
box -12 -8 32 272
use FILL  FILL_3__2876_
timestamp 1701859473
transform -1 0 9730 0 1 1830
box -12 -8 32 272
use FILL  FILL_3__2877_
timestamp 1701859473
transform 1 0 9910 0 1 1830
box -12 -8 32 272
use FILL  FILL_3__2878_
timestamp 1701859473
transform 1 0 9730 0 -1 1310
box -12 -8 32 272
use FILL  FILL_3__2879_
timestamp 1701859473
transform -1 0 9970 0 -1 1310
box -12 -8 32 272
use FILL  FILL_3__2880_
timestamp 1701859473
transform 1 0 9470 0 1 1830
box -12 -8 32 272
use FILL  FILL_3__2881_
timestamp 1701859473
transform 1 0 10850 0 -1 790
box -12 -8 32 272
use FILL  FILL_3__2882_
timestamp 1701859473
transform -1 0 9530 0 -1 1310
box -12 -8 32 272
use FILL  FILL_3__2883_
timestamp 1701859473
transform -1 0 10430 0 -1 1310
box -12 -8 32 272
use FILL  FILL_3__2884_
timestamp 1701859473
transform 1 0 11070 0 -1 1310
box -12 -8 32 272
use FILL  FILL_3__2885_
timestamp 1701859473
transform -1 0 10850 0 -1 1310
box -12 -8 32 272
use FILL  FILL_3__2886_
timestamp 1701859473
transform 1 0 10610 0 1 1830
box -12 -8 32 272
use FILL  FILL_3__2887_
timestamp 1701859473
transform 1 0 10170 0 -1 4430
box -12 -8 32 272
use FILL  FILL_3__2888_
timestamp 1701859473
transform -1 0 3990 0 1 5470
box -12 -8 32 272
use FILL  FILL_3__2889_
timestamp 1701859473
transform 1 0 6110 0 1 2350
box -12 -8 32 272
use FILL  FILL_3__2890_
timestamp 1701859473
transform -1 0 8390 0 1 5990
box -12 -8 32 272
use FILL  FILL_3__2891_
timestamp 1701859473
transform -1 0 8190 0 1 5990
box -12 -8 32 272
use FILL  FILL_3__2892_
timestamp 1701859473
transform 1 0 7410 0 -1 5470
box -12 -8 32 272
use FILL  FILL_3__2893_
timestamp 1701859473
transform 1 0 7230 0 1 5470
box -12 -8 32 272
use FILL  FILL_3__2894_
timestamp 1701859473
transform 1 0 6510 0 -1 6510
box -12 -8 32 272
use FILL  FILL_3__2895_
timestamp 1701859473
transform 1 0 6650 0 1 6510
box -12 -8 32 272
use FILL  FILL_3__2896_
timestamp 1701859473
transform -1 0 7910 0 -1 5470
box -12 -8 32 272
use FILL  FILL_3__2897_
timestamp 1701859473
transform 1 0 7710 0 1 5470
box -12 -8 32 272
use FILL  FILL_3__2898_
timestamp 1701859473
transform 1 0 7230 0 -1 6510
box -12 -8 32 272
use FILL  FILL_3__2899_
timestamp 1701859473
transform 1 0 6750 0 -1 6510
box -12 -8 32 272
use FILL  FILL_3__2900_
timestamp 1701859473
transform -1 0 6290 0 -1 6510
box -12 -8 32 272
use FILL  FILL_3__2901_
timestamp 1701859473
transform 1 0 6030 0 -1 6510
box -12 -8 32 272
use FILL  FILL_3__2902_
timestamp 1701859473
transform -1 0 7950 0 1 5990
box -12 -8 32 272
use FILL  FILL_3__2903_
timestamp 1701859473
transform 1 0 7230 0 1 5990
box -12 -8 32 272
use FILL  FILL_3__2904_
timestamp 1701859473
transform 1 0 8350 0 -1 5470
box -12 -8 32 272
use FILL  FILL_3__2905_
timestamp 1701859473
transform 1 0 8370 0 1 5470
box -12 -8 32 272
use FILL  FILL_3__2906_
timestamp 1701859473
transform 1 0 8110 0 -1 5990
box -12 -8 32 272
use FILL  FILL_3__2907_
timestamp 1701859473
transform -1 0 7890 0 -1 5990
box -12 -8 32 272
use FILL  FILL_3__2908_
timestamp 1701859473
transform -1 0 8210 0 -1 4950
box -12 -8 32 272
use FILL  FILL_3__2909_
timestamp 1701859473
transform 1 0 3350 0 -1 4430
box -12 -8 32 272
use FILL  FILL_3__2910_
timestamp 1701859473
transform -1 0 6510 0 -1 4430
box -12 -8 32 272
use FILL  FILL_3__2911_
timestamp 1701859473
transform -1 0 6850 0 1 4430
box -12 -8 32 272
use FILL  FILL_3__2912_
timestamp 1701859473
transform 1 0 8630 0 -1 4950
box -12 -8 32 272
use FILL  FILL_3__2913_
timestamp 1701859473
transform -1 0 6810 0 -1 4950
box -12 -8 32 272
use FILL  FILL_3__2914_
timestamp 1701859473
transform 1 0 7070 0 -1 8070
box -12 -8 32 272
use FILL  FILL_3__2915_
timestamp 1701859473
transform 1 0 7190 0 -1 5990
box -12 -8 32 272
use FILL  FILL_3__2916_
timestamp 1701859473
transform 1 0 6950 0 -1 5990
box -12 -8 32 272
use FILL  FILL_3__2917_
timestamp 1701859473
transform -1 0 6330 0 -1 5990
box -12 -8 32 272
use FILL  FILL_3__2918_
timestamp 1701859473
transform 1 0 6250 0 1 5470
box -12 -8 32 272
use FILL  FILL_3__2919_
timestamp 1701859473
transform 1 0 6170 0 1 4950
box -12 -8 32 272
use FILL  FILL_3__2920_
timestamp 1701859473
transform 1 0 5930 0 1 4950
box -12 -8 32 272
use FILL  FILL_3__2921_
timestamp 1701859473
transform -1 0 7390 0 -1 3910
box -12 -8 32 272
use FILL  FILL_3__2922_
timestamp 1701859473
transform -1 0 7430 0 1 3910
box -12 -8 32 272
use FILL  FILL_3__2923_
timestamp 1701859473
transform -1 0 6750 0 -1 4430
box -12 -8 32 272
use FILL  FILL_3__2924_
timestamp 1701859473
transform 1 0 6370 0 1 4950
box -12 -8 32 272
use FILL  FILL_3__2925_
timestamp 1701859473
transform 1 0 7270 0 1 7550
box -12 -8 32 272
use FILL  FILL_3__2926_
timestamp 1701859473
transform -1 0 7510 0 1 4430
box -12 -8 32 272
use FILL  FILL_3__2927_
timestamp 1701859473
transform 1 0 7290 0 -1 4950
box -12 -8 32 272
use FILL  FILL_3__2928_
timestamp 1701859473
transform 1 0 7030 0 -1 4950
box -12 -8 32 272
use FILL  FILL_3__2929_
timestamp 1701859473
transform -1 0 6610 0 1 4950
box -12 -8 32 272
use FILL  FILL_3__2930_
timestamp 1701859473
transform 1 0 6150 0 1 1830
box -12 -8 32 272
use FILL  FILL_3__2931_
timestamp 1701859473
transform 1 0 7030 0 -1 2870
box -12 -8 32 272
use FILL  FILL_3__2932_
timestamp 1701859473
transform 1 0 5190 0 -1 4430
box -12 -8 32 272
use FILL  FILL_3__2933_
timestamp 1701859473
transform 1 0 5390 0 -1 4430
box -12 -8 32 272
use FILL  FILL_3__2934_
timestamp 1701859473
transform 1 0 5630 0 -1 4430
box -12 -8 32 272
use FILL  FILL_3__2935_
timestamp 1701859473
transform 1 0 6450 0 1 6510
box -12 -8 32 272
use FILL  FILL_3__2936_
timestamp 1701859473
transform 1 0 6330 0 -1 4950
box -12 -8 32 272
use FILL  FILL_3__2937_
timestamp 1701859473
transform 1 0 6550 0 -1 4950
box -12 -8 32 272
use FILL  FILL_3__2938_
timestamp 1701859473
transform 1 0 5030 0 1 4950
box -12 -8 32 272
use FILL  FILL_3__2939_
timestamp 1701859473
transform 1 0 4810 0 1 4950
box -12 -8 32 272
use FILL  FILL_3__2940_
timestamp 1701859473
transform -1 0 5870 0 -1 5470
box -12 -8 32 272
use FILL  FILL_3__2941_
timestamp 1701859473
transform 1 0 5630 0 -1 5470
box -12 -8 32 272
use FILL  FILL_3__2942_
timestamp 1701859473
transform -1 0 9330 0 1 4430
box -12 -8 32 272
use FILL  FILL_3__2943_
timestamp 1701859473
transform 1 0 6290 0 -1 4430
box -12 -8 32 272
use FILL  FILL_3__2944_
timestamp 1701859473
transform -1 0 6310 0 1 3910
box -12 -8 32 272
use FILL  FILL_3__2945_
timestamp 1701859473
transform -1 0 6390 0 1 4430
box -12 -8 32 272
use FILL  FILL_3__2946_
timestamp 1701859473
transform 1 0 6150 0 1 4430
box -12 -8 32 272
use FILL  FILL_3__2947_
timestamp 1701859473
transform -1 0 6550 0 -1 5990
box -12 -8 32 272
use FILL  FILL_3__2948_
timestamp 1701859473
transform 1 0 6090 0 -1 5990
box -12 -8 32 272
use FILL  FILL_3__2949_
timestamp 1701859473
transform -1 0 5910 0 -1 5990
box -12 -8 32 272
use FILL  FILL_3__2950_
timestamp 1701859473
transform 1 0 5770 0 1 5470
box -12 -8 32 272
use FILL  FILL_3__2951_
timestamp 1701859473
transform -1 0 6030 0 1 5470
box -12 -8 32 272
use FILL  FILL_3__2952_
timestamp 1701859473
transform -1 0 6110 0 -1 4950
box -12 -8 32 272
use FILL  FILL_3__2953_
timestamp 1701859473
transform -1 0 4390 0 1 4950
box -12 -8 32 272
use FILL  FILL_3__2954_
timestamp 1701859473
transform -1 0 6650 0 1 4430
box -12 -8 32 272
use FILL  FILL_3__2955_
timestamp 1701859473
transform -1 0 5930 0 1 4430
box -12 -8 32 272
use FILL  FILL_3__2956_
timestamp 1701859473
transform 1 0 5210 0 1 4430
box -12 -8 32 272
use FILL  FILL_3__2957_
timestamp 1701859473
transform 1 0 5150 0 -1 4950
box -12 -8 32 272
use FILL  FILL_3__2958_
timestamp 1701859473
transform -1 0 5470 0 1 4430
box -12 -8 32 272
use FILL  FILL_3__2959_
timestamp 1701859473
transform 1 0 6970 0 -1 5470
box -12 -8 32 272
use FILL  FILL_3__2960_
timestamp 1701859473
transform -1 0 6510 0 1 5470
box -12 -8 32 272
use FILL  FILL_3__2961_
timestamp 1701859473
transform 1 0 6270 0 -1 5470
box -12 -8 32 272
use FILL  FILL_3__2962_
timestamp 1701859473
transform -1 0 6530 0 -1 5470
box -12 -8 32 272
use FILL  FILL_3__2963_
timestamp 1701859473
transform -1 0 6770 0 -1 5470
box -12 -8 32 272
use FILL  FILL_3__2964_
timestamp 1701859473
transform -1 0 5410 0 -1 4950
box -12 -8 32 272
use FILL  FILL_3__2965_
timestamp 1701859473
transform 1 0 4910 0 -1 4950
box -12 -8 32 272
use FILL  FILL_3__2966_
timestamp 1701859473
transform -1 0 6370 0 1 2350
box -12 -8 32 272
use FILL  FILL_3__2967_
timestamp 1701859473
transform 1 0 7630 0 1 3910
box -12 -8 32 272
use FILL  FILL_3__2968_
timestamp 1701859473
transform -1 0 6950 0 -1 3910
box -12 -8 32 272
use FILL  FILL_3__2969_
timestamp 1701859473
transform -1 0 7170 0 -1 3910
box -12 -8 32 272
use FILL  FILL_3__2970_
timestamp 1701859473
transform -1 0 7210 0 1 3910
box -12 -8 32 272
use FILL  FILL_3__2971_
timestamp 1701859473
transform -1 0 6730 0 1 3910
box -12 -8 32 272
use FILL  FILL_3__2972_
timestamp 1701859473
transform 1 0 6950 0 1 3910
box -12 -8 32 272
use FILL  FILL_3__2973_
timestamp 1701859473
transform -1 0 7070 0 1 4430
box -12 -8 32 272
use FILL  FILL_3__2974_
timestamp 1701859473
transform 1 0 6970 0 -1 4430
box -12 -8 32 272
use FILL  FILL_3__2975_
timestamp 1701859473
transform -1 0 7730 0 -1 4430
box -12 -8 32 272
use FILL  FILL_3__2976_
timestamp 1701859473
transform -1 0 7490 0 -1 4430
box -12 -8 32 272
use FILL  FILL_3__2977_
timestamp 1701859473
transform 1 0 7210 0 -1 4430
box -12 -8 32 272
use FILL  FILL_3__2978_
timestamp 1701859473
transform 1 0 7270 0 1 4430
box -12 -8 32 272
use FILL  FILL_3__2979_
timestamp 1701859473
transform -1 0 3610 0 -1 4950
box -12 -8 32 272
use FILL  FILL_3__2980_
timestamp 1701859473
transform -1 0 2990 0 1 7550
box -12 -8 32 272
use FILL  FILL_3__2981_
timestamp 1701859473
transform 1 0 3510 0 1 4950
box -12 -8 32 272
use FILL  FILL_3__2982_
timestamp 1701859473
transform 1 0 9570 0 1 6510
box -12 -8 32 272
use FILL  FILL_3__2983_
timestamp 1701859473
transform 1 0 1890 0 1 4430
box -12 -8 32 272
use FILL  FILL_3__2984_
timestamp 1701859473
transform -1 0 3510 0 -1 3910
box -12 -8 32 272
use FILL  FILL_3__2985_
timestamp 1701859473
transform 1 0 3670 0 1 4430
box -12 -8 32 272
use FILL  FILL_3__2986_
timestamp 1701859473
transform -1 0 5870 0 -1 4430
box -12 -8 32 272
use FILL  FILL_3__2987_
timestamp 1701859473
transform -1 0 5690 0 1 4430
box -12 -8 32 272
use FILL  FILL_3__2988_
timestamp 1701859473
transform 1 0 9350 0 1 6510
box -12 -8 32 272
use FILL  FILL_3__2989_
timestamp 1701859473
transform 1 0 5970 0 1 6510
box -12 -8 32 272
use FILL  FILL_3__2990_
timestamp 1701859473
transform -1 0 6230 0 1 6510
box -12 -8 32 272
use FILL  FILL_3__2991_
timestamp 1701859473
transform 1 0 7130 0 1 6510
box -12 -8 32 272
use FILL  FILL_3__2992_
timestamp 1701859473
transform 1 0 9650 0 1 7030
box -12 -8 32 272
use FILL  FILL_3__2993_
timestamp 1701859473
transform 1 0 9850 0 1 7030
box -12 -8 32 272
use FILL  FILL_3__2994_
timestamp 1701859473
transform -1 0 10770 0 -1 7550
box -12 -8 32 272
use FILL  FILL_3__2995_
timestamp 1701859473
transform -1 0 7570 0 -1 7550
box -12 -8 32 272
use FILL  FILL_3__2996_
timestamp 1701859473
transform 1 0 7470 0 1 7550
box -12 -8 32 272
use FILL  FILL_3__2997_
timestamp 1701859473
transform -1 0 7350 0 -1 7550
box -12 -8 32 272
use FILL  FILL_3__2998_
timestamp 1701859473
transform -1 0 6410 0 -1 7550
box -12 -8 32 272
use FILL  FILL_3__2999_
timestamp 1701859473
transform 1 0 6130 0 1 7550
box -12 -8 32 272
use FILL  FILL_3__3000_
timestamp 1701859473
transform -1 0 5970 0 -1 7550
box -12 -8 32 272
use FILL  FILL_3__3001_
timestamp 1701859473
transform -1 0 5750 0 -1 7550
box -12 -8 32 272
use FILL  FILL_3__3002_
timestamp 1701859473
transform -1 0 6170 0 -1 7550
box -12 -8 32 272
use FILL  FILL_3__3003_
timestamp 1701859473
transform -1 0 6350 0 1 7550
box -12 -8 32 272
use FILL  FILL_3__3004_
timestamp 1701859473
transform 1 0 8150 0 1 7550
box -12 -8 32 272
use FILL  FILL_3__3005_
timestamp 1701859473
transform 1 0 10970 0 -1 7550
box -12 -8 32 272
use FILL  FILL_3__3006_
timestamp 1701859473
transform -1 0 10450 0 1 7550
box -12 -8 32 272
use FILL  FILL_3__3007_
timestamp 1701859473
transform 1 0 6970 0 1 7030
box -12 -8 32 272
use FILL  FILL_3__3008_
timestamp 1701859473
transform -1 0 6530 0 1 7030
box -12 -8 32 272
use FILL  FILL_3__3009_
timestamp 1701859473
transform -1 0 5930 0 -1 7030
box -12 -8 32 272
use FILL  FILL_3__3010_
timestamp 1701859473
transform 1 0 6150 0 -1 7030
box -12 -8 32 272
use FILL  FILL_3__3011_
timestamp 1701859473
transform 1 0 6730 0 1 7030
box -12 -8 32 272
use FILL  FILL_3__3012_
timestamp 1701859473
transform -1 0 7850 0 -1 7030
box -12 -8 32 272
use FILL  FILL_3__3013_
timestamp 1701859473
transform 1 0 8290 0 -1 7030
box -12 -8 32 272
use FILL  FILL_3__3014_
timestamp 1701859473
transform 1 0 10650 0 1 7550
box -12 -8 32 272
use FILL  FILL_3__3015_
timestamp 1701859473
transform -1 0 6370 0 -1 7030
box -12 -8 32 272
use FILL  FILL_3__3016_
timestamp 1701859473
transform -1 0 7250 0 1 7030
box -12 -8 32 272
use FILL  FILL_3__3017_
timestamp 1701859473
transform 1 0 6590 0 -1 7030
box -12 -8 32 272
use FILL  FILL_3__3018_
timestamp 1701859473
transform -1 0 6890 0 -1 7030
box -12 -8 32 272
use FILL  FILL_3__3019_
timestamp 1701859473
transform -1 0 7130 0 -1 7030
box -12 -8 32 272
use FILL  FILL_3__3020_
timestamp 1701859473
transform 1 0 8290 0 1 7030
box -12 -8 32 272
use FILL  FILL_3__3021_
timestamp 1701859473
transform -1 0 9350 0 -1 8070
box -12 -8 32 272
use FILL  FILL_3__3022_
timestamp 1701859473
transform 1 0 9530 0 -1 8070
box -12 -8 32 272
use FILL  FILL_3__3023_
timestamp 1701859473
transform -1 0 5750 0 1 6510
box -12 -8 32 272
use FILL  FILL_3__3024_
timestamp 1701859473
transform 1 0 5490 0 1 6510
box -12 -8 32 272
use FILL  FILL_3__3025_
timestamp 1701859473
transform -1 0 5510 0 -1 6510
box -12 -8 32 272
use FILL  FILL_3__3026_
timestamp 1701859473
transform 1 0 10930 0 -1 5990
box -12 -8 32 272
use FILL  FILL_3__3027_
timestamp 1701859473
transform -1 0 11170 0 -1 5990
box -12 -8 32 272
use FILL  FILL_3__3028_
timestamp 1701859473
transform -1 0 9790 0 -1 8070
box -12 -8 32 272
use FILL  FILL_3__3029_
timestamp 1701859473
transform -1 0 7110 0 -1 7550
box -12 -8 32 272
use FILL  FILL_3__3030_
timestamp 1701859473
transform -1 0 8090 0 -1 7030
box -12 -8 32 272
use FILL  FILL_3__3031_
timestamp 1701859473
transform 1 0 8070 0 1 7030
box -12 -8 32 272
use FILL  FILL_3__3032_
timestamp 1701859473
transform 1 0 7690 0 1 7550
box -12 -8 32 272
use FILL  FILL_3__3033_
timestamp 1701859473
transform -1 0 6770 0 1 8070
box -12 -8 32 272
use FILL  FILL_3__3034_
timestamp 1701859473
transform -1 0 7750 0 -1 8070
box -12 -8 32 272
use FILL  FILL_3__3035_
timestamp 1701859473
transform 1 0 7490 0 -1 8070
box -12 -8 32 272
use FILL  FILL_3__3036_
timestamp 1701859473
transform -1 0 6970 0 1 8070
box -12 -8 32 272
use FILL  FILL_3__3037_
timestamp 1701859473
transform -1 0 6530 0 1 8070
box -12 -8 32 272
use FILL  FILL_3__3038_
timestamp 1701859473
transform -1 0 7150 0 1 8070
box -12 -8 32 272
use FILL  FILL_3__3039_
timestamp 1701859473
transform 1 0 7370 0 1 8070
box -12 -8 32 272
use FILL  FILL_3__3040_
timestamp 1701859473
transform 1 0 9710 0 1 7550
box -12 -8 32 272
use FILL  FILL_3__3041_
timestamp 1701859473
transform -1 0 9570 0 -1 6510
box -12 -8 32 272
use FILL  FILL_3__3042_
timestamp 1701859473
transform 1 0 7270 0 -1 8070
box -12 -8 32 272
use FILL  FILL_3__3043_
timestamp 1701859473
transform -1 0 6590 0 1 7550
box -12 -8 32 272
use FILL  FILL_3__3044_
timestamp 1701859473
transform -1 0 6630 0 -1 7550
box -12 -8 32 272
use FILL  FILL_3__3045_
timestamp 1701859473
transform 1 0 6850 0 -1 7550
box -12 -8 32 272
use FILL  FILL_3__3046_
timestamp 1701859473
transform -1 0 7810 0 1 6510
box -12 -8 32 272
use FILL  FILL_3__3047_
timestamp 1701859473
transform 1 0 9150 0 1 6510
box -12 -8 32 272
use FILL  FILL_3__3048_
timestamp 1701859473
transform 1 0 9770 0 -1 6510
box -12 -8 32 272
use FILL  FILL_3__3049_
timestamp 1701859473
transform -1 0 6850 0 1 7550
box -12 -8 32 272
use FILL  FILL_3__3050_
timestamp 1701859473
transform -1 0 7070 0 1 7550
box -12 -8 32 272
use FILL  FILL_3__3051_
timestamp 1701859473
transform -1 0 7810 0 1 7030
box -12 -8 32 272
use FILL  FILL_3__3052_
timestamp 1701859473
transform 1 0 7510 0 1 7030
box -12 -8 32 272
use FILL  FILL_3__3053_
timestamp 1701859473
transform 1 0 7350 0 -1 7030
box -12 -8 32 272
use FILL  FILL_3__3054_
timestamp 1701859473
transform -1 0 7610 0 -1 7030
box -12 -8 32 272
use FILL  FILL_3__3055_
timestamp 1701859473
transform 1 0 8030 0 1 6510
box -12 -8 32 272
use FILL  FILL_3__3056_
timestamp 1701859473
transform -1 0 9550 0 1 5470
box -12 -8 32 272
use FILL  FILL_3__3057_
timestamp 1701859473
transform -1 0 9310 0 1 5470
box -12 -8 32 272
use FILL  FILL_3__3058_
timestamp 1701859473
transform 1 0 8730 0 -1 7550
box -12 -8 32 272
use FILL  FILL_3__3059_
timestamp 1701859473
transform -1 0 8610 0 -1 5990
box -12 -8 32 272
use FILL  FILL_3__3060_
timestamp 1701859473
transform 1 0 9790 0 1 6510
box -12 -8 32 272
use FILL  FILL_3__3061_
timestamp 1701859473
transform 1 0 10030 0 1 6510
box -12 -8 32 272
use FILL  FILL_3__3062_
timestamp 1701859473
transform -1 0 9650 0 -1 7550
box -12 -8 32 272
use FILL  FILL_3__3063_
timestamp 1701859473
transform 1 0 9390 0 -1 7550
box -12 -8 32 272
use FILL  FILL_3__3064_
timestamp 1701859473
transform -1 0 10350 0 -1 7030
box -12 -8 32 272
use FILL  FILL_3__3065_
timestamp 1701859473
transform -1 0 10590 0 -1 7030
box -12 -8 32 272
use FILL  FILL_3__3066_
timestamp 1701859473
transform -1 0 8510 0 -1 7550
box -12 -8 32 272
use FILL  FILL_3__3067_
timestamp 1701859473
transform 1 0 8250 0 -1 7550
box -12 -8 32 272
use FILL  FILL_3__3068_
timestamp 1701859473
transform 1 0 10210 0 -1 5990
box -12 -8 32 272
use FILL  FILL_3__3069_
timestamp 1701859473
transform 1 0 10450 0 -1 5990
box -12 -8 32 272
use FILL  FILL_3__3070_
timestamp 1701859473
transform 1 0 8910 0 -1 7550
box -12 -8 32 272
use FILL  FILL_3__3071_
timestamp 1701859473
transform -1 0 9170 0 -1 7550
box -12 -8 32 272
use FILL  FILL_3__3072_
timestamp 1701859473
transform -1 0 9790 0 1 5990
box -12 -8 32 272
use FILL  FILL_3__3073_
timestamp 1701859473
transform -1 0 10010 0 1 5990
box -12 -8 32 272
use FILL  FILL_3__3074_
timestamp 1701859473
transform 1 0 8830 0 1 5990
box -12 -8 32 272
use FILL  FILL_3__3075_
timestamp 1701859473
transform 1 0 8830 0 -1 5990
box -12 -8 32 272
use FILL  FILL_3__3076_
timestamp 1701859473
transform 1 0 10730 0 1 6510
box -12 -8 32 272
use FILL  FILL_3__3077_
timestamp 1701859473
transform 1 0 10930 0 1 6510
box -12 -8 32 272
use FILL  FILL_3__3078_
timestamp 1701859473
transform -1 0 8730 0 -1 7030
box -12 -8 32 272
use FILL  FILL_3__3079_
timestamp 1701859473
transform -1 0 8510 0 -1 7030
box -12 -8 32 272
use FILL  FILL_3__3080_
timestamp 1701859473
transform 1 0 10990 0 -1 8590
box -12 -8 32 272
use FILL  FILL_3__3081_
timestamp 1701859473
transform -1 0 10990 0 -1 270
box -12 -8 32 272
use FILL  FILL_3__3082_
timestamp 1701859473
transform 1 0 10090 0 -1 8590
box -12 -8 32 272
use FILL  FILL_3__3083_
timestamp 1701859473
transform -1 0 9870 0 -1 8590
box -12 -8 32 272
use FILL  FILL_3__3084_
timestamp 1701859473
transform -1 0 9050 0 1 7550
box -12 -8 32 272
use FILL  FILL_3__3085_
timestamp 1701859473
transform 1 0 8950 0 1 7030
box -12 -8 32 272
use FILL  FILL_3__3086_
timestamp 1701859473
transform -1 0 10710 0 1 5990
box -12 -8 32 272
use FILL  FILL_3__3087_
timestamp 1701859473
transform 1 0 10910 0 1 5990
box -12 -8 32 272
use FILL  FILL_3__3088_
timestamp 1701859473
transform 1 0 8270 0 1 8070
box -12 -8 32 272
use FILL  FILL_3__3089_
timestamp 1701859473
transform -1 0 8050 0 1 8070
box -12 -8 32 272
use FILL  FILL_3__3090_
timestamp 1701859473
transform -1 0 11150 0 1 4950
box -12 -8 32 272
use FILL  FILL_3__3091_
timestamp 1701859473
transform 1 0 10890 0 1 4950
box -12 -8 32 272
use FILL  FILL_3__3092_
timestamp 1701859473
transform 1 0 8810 0 -1 5470
box -12 -8 32 272
use FILL  FILL_3__3093_
timestamp 1701859473
transform -1 0 9050 0 -1 5470
box -12 -8 32 272
use FILL  FILL_3__3094_
timestamp 1701859473
transform -1 0 10250 0 -1 5470
box -12 -8 32 272
use FILL  FILL_3__3095_
timestamp 1701859473
transform 1 0 10190 0 1 5470
box -12 -8 32 272
use FILL  FILL_3__3096_
timestamp 1701859473
transform 1 0 8930 0 1 6510
box -12 -8 32 272
use FILL  FILL_3__3097_
timestamp 1701859473
transform -1 0 8710 0 1 6510
box -12 -8 32 272
use FILL  FILL_3__3098_
timestamp 1701859473
transform -1 0 10410 0 1 8070
box -12 -8 32 272
use FILL  FILL_3__3099_
timestamp 1701859473
transform -1 0 11170 0 -1 8070
box -12 -8 32 272
use FILL  FILL_3__3100_
timestamp 1701859473
transform 1 0 10170 0 1 8070
box -12 -8 32 272
use FILL  FILL_3__3101_
timestamp 1701859473
transform 1 0 10310 0 -1 8590
box -12 -8 32 272
use FILL  FILL_3__3102_
timestamp 1701859473
transform 1 0 8390 0 -1 8070
box -12 -8 32 272
use FILL  FILL_3__3103_
timestamp 1701859473
transform -1 0 8370 0 1 7550
box -12 -8 32 272
use FILL  FILL_3__3104_
timestamp 1701859473
transform -1 0 11170 0 1 6510
box -12 -8 32 272
use FILL  FILL_3__3105_
timestamp 1701859473
transform -1 0 10970 0 -1 4950
box -12 -8 32 272
use FILL  FILL_3__3106_
timestamp 1701859473
transform 1 0 9390 0 -1 8590
box -12 -8 32 272
use FILL  FILL_3__3107_
timestamp 1701859473
transform -1 0 9630 0 -1 8590
box -12 -8 32 272
use FILL  FILL_3__3108_
timestamp 1701859473
transform 1 0 9990 0 1 5470
box -12 -8 32 272
use FILL  FILL_3__3109_
timestamp 1701859473
transform -1 0 9770 0 1 5470
box -12 -8 32 272
use FILL  FILL_3__3110_
timestamp 1701859473
transform 1 0 8410 0 -1 6510
box -12 -8 32 272
use FILL  FILL_3__3111_
timestamp 1701859473
transform -1 0 8190 0 -1 6510
box -12 -8 32 272
use FILL  FILL_3__3112_
timestamp 1701859473
transform 1 0 530 0 -1 2870
box -12 -8 32 272
use FILL  FILL_3__3113_
timestamp 1701859473
transform 1 0 70 0 -1 2870
box -12 -8 32 272
use FILL  FILL_3__3114_
timestamp 1701859473
transform -1 0 330 0 -1 2870
box -12 -8 32 272
use FILL  FILL_3__3115_
timestamp 1701859473
transform -1 0 1210 0 1 2350
box -12 -8 32 272
use FILL  FILL_3__3116_
timestamp 1701859473
transform 1 0 970 0 -1 2350
box -12 -8 32 272
use FILL  FILL_3__3117_
timestamp 1701859473
transform 1 0 2050 0 -1 1310
box -12 -8 32 272
use FILL  FILL_3__3118_
timestamp 1701859473
transform -1 0 1430 0 -1 2350
box -12 -8 32 272
use FILL  FILL_3__3119_
timestamp 1701859473
transform -1 0 1190 0 -1 2350
box -12 -8 32 272
use FILL  FILL_3__3120_
timestamp 1701859473
transform -1 0 490 0 1 2350
box -12 -8 32 272
use FILL  FILL_3__3121_
timestamp 1701859473
transform 1 0 270 0 1 2870
box -12 -8 32 272
use FILL  FILL_3__3122_
timestamp 1701859473
transform 1 0 2530 0 -1 3390
box -12 -8 32 272
use FILL  FILL_3__3123_
timestamp 1701859473
transform 1 0 550 0 1 3390
box -12 -8 32 272
use FILL  FILL_3__3124_
timestamp 1701859473
transform -1 0 330 0 1 3390
box -12 -8 32 272
use FILL  FILL_3__3125_
timestamp 1701859473
transform -1 0 750 0 -1 2350
box -12 -8 32 272
use FILL  FILL_3__3126_
timestamp 1701859473
transform -1 0 1450 0 1 2350
box -12 -8 32 272
use FILL  FILL_3__3127_
timestamp 1701859473
transform -1 0 970 0 1 2350
box -12 -8 32 272
use FILL  FILL_3__3128_
timestamp 1701859473
transform -1 0 1910 0 1 2350
box -12 -8 32 272
use FILL  FILL_3__3129_
timestamp 1701859473
transform -1 0 1670 0 -1 2350
box -12 -8 32 272
use FILL  FILL_3__3130_
timestamp 1701859473
transform -1 0 1690 0 1 2350
box -12 -8 32 272
use FILL  FILL_3__3131_
timestamp 1701859473
transform -1 0 730 0 1 2350
box -12 -8 32 272
use FILL  FILL_3__3132_
timestamp 1701859473
transform 1 0 490 0 1 2870
box -12 -8 32 272
use FILL  FILL_3__3133_
timestamp 1701859473
transform 1 0 550 0 -1 3910
box -12 -8 32 272
use FILL  FILL_3__3134_
timestamp 1701859473
transform -1 0 1230 0 1 3390
box -12 -8 32 272
use FILL  FILL_3__3135_
timestamp 1701859473
transform 1 0 990 0 1 3390
box -12 -8 32 272
use FILL  FILL_3__3136_
timestamp 1701859473
transform -1 0 570 0 -1 3390
box -12 -8 32 272
use FILL  FILL_3__3137_
timestamp 1701859473
transform 1 0 290 0 -1 3390
box -12 -8 32 272
use FILL  FILL_3__3138_
timestamp 1701859473
transform -1 0 1690 0 1 4430
box -12 -8 32 272
use FILL  FILL_3__3139_
timestamp 1701859473
transform -1 0 1890 0 -1 3390
box -12 -8 32 272
use FILL  FILL_3__3140_
timestamp 1701859473
transform -1 0 310 0 1 3910
box -12 -8 32 272
use FILL  FILL_3__3141_
timestamp 1701859473
transform 1 0 750 0 1 4430
box -12 -8 32 272
use FILL  FILL_3__3142_
timestamp 1701859473
transform 1 0 990 0 1 4430
box -12 -8 32 272
use FILL  FILL_3__3143_
timestamp 1701859473
transform 1 0 1010 0 -1 4430
box -12 -8 32 272
use FILL  FILL_3__3144_
timestamp 1701859473
transform -1 0 1250 0 -1 4430
box -12 -8 32 272
use FILL  FILL_3__3145_
timestamp 1701859473
transform -1 0 530 0 1 3910
box -12 -8 32 272
use FILL  FILL_3__3146_
timestamp 1701859473
transform -1 0 750 0 1 3910
box -12 -8 32 272
use FILL  FILL_3__3147_
timestamp 1701859473
transform 1 0 530 0 -1 4430
box -12 -8 32 272
use FILL  FILL_3__3148_
timestamp 1701859473
transform -1 0 790 0 -1 4430
box -12 -8 32 272
use FILL  FILL_3__3149_
timestamp 1701859473
transform -1 0 90 0 -1 3910
box -12 -8 32 272
use FILL  FILL_3__3150_
timestamp 1701859473
transform -1 0 950 0 1 3910
box -12 -8 32 272
use FILL  FILL_3__3151_
timestamp 1701859473
transform 1 0 70 0 1 3910
box -12 -8 32 272
use FILL  FILL_3__3152_
timestamp 1701859473
transform 1 0 70 0 -1 4430
box -12 -8 32 272
use FILL  FILL_3__3153_
timestamp 1701859473
transform -1 0 310 0 -1 4430
box -12 -8 32 272
use FILL  FILL_3__3154_
timestamp 1701859473
transform -1 0 810 0 -1 3390
box -12 -8 32 272
use FILL  FILL_3__3155_
timestamp 1701859473
transform -1 0 90 0 1 2870
box -12 -8 32 272
use FILL  FILL_3__3156_
timestamp 1701859473
transform 1 0 70 0 -1 3390
box -12 -8 32 272
use FILL  FILL_3__3157_
timestamp 1701859473
transform -1 0 90 0 1 3390
box -12 -8 32 272
use FILL  FILL_3__3158_
timestamp 1701859473
transform 1 0 70 0 1 4430
box -12 -8 32 272
use FILL  FILL_3__3159_
timestamp 1701859473
transform 1 0 290 0 1 4430
box -12 -8 32 272
use FILL  FILL_3__3160_
timestamp 1701859473
transform -1 0 530 0 1 4430
box -12 -8 32 272
use FILL  FILL_3__3161_
timestamp 1701859473
transform 1 0 4170 0 -1 7030
box -12 -8 32 272
use FILL  FILL_3__3162_
timestamp 1701859473
transform -1 0 4410 0 -1 7030
box -12 -8 32 272
use FILL  FILL_3__3163_
timestamp 1701859473
transform 1 0 4630 0 -1 7030
box -12 -8 32 272
use FILL  FILL_3__3164_
timestamp 1701859473
transform 1 0 4870 0 1 7030
box -12 -8 32 272
use FILL  FILL_3__3165_
timestamp 1701859473
transform 1 0 4130 0 1 7550
box -12 -8 32 272
use FILL  FILL_3__3166_
timestamp 1701859473
transform -1 0 4370 0 1 7550
box -12 -8 32 272
use FILL  FILL_3__3167_
timestamp 1701859473
transform 1 0 4850 0 -1 10150
box -12 -8 32 272
use FILL  FILL_3__3168_
timestamp 1701859473
transform 1 0 5050 0 -1 10150
box -12 -8 32 272
use FILL  FILL_3__3169_
timestamp 1701859473
transform -1 0 3690 0 -1 10670
box -12 -8 32 272
use FILL  FILL_3__3170_
timestamp 1701859473
transform -1 0 3910 0 -1 10670
box -12 -8 32 272
use FILL  FILL_3__3171_
timestamp 1701859473
transform 1 0 4330 0 -1 10670
box -12 -8 32 272
use FILL  FILL_3__3172_
timestamp 1701859473
transform -1 0 4570 0 -1 10670
box -12 -8 32 272
use FILL  FILL_3__3173_
timestamp 1701859473
transform 1 0 4170 0 1 10150
box -12 -8 32 272
use FILL  FILL_3__3174_
timestamp 1701859473
transform -1 0 4410 0 1 10150
box -12 -8 32 272
use FILL  FILL_3__3175_
timestamp 1701859473
transform 1 0 5510 0 1 10150
box -12 -8 32 272
use FILL  FILL_3__3176_
timestamp 1701859473
transform 1 0 5270 0 1 10150
box -12 -8 32 272
use FILL  FILL_3__3177_
timestamp 1701859473
transform -1 0 1750 0 -1 5990
box -12 -8 32 272
use FILL  FILL_3__3178_
timestamp 1701859473
transform 1 0 2190 0 -1 5990
box -12 -8 32 272
use FILL  FILL_3__3179_
timestamp 1701859473
transform -1 0 1470 0 1 6510
box -12 -8 32 272
use FILL  FILL_3__3180_
timestamp 1701859473
transform -1 0 1690 0 1 6510
box -12 -8 32 272
use FILL  FILL_3__3181_
timestamp 1701859473
transform -1 0 550 0 -1 6510
box -12 -8 32 272
use FILL  FILL_3__3182_
timestamp 1701859473
transform -1 0 950 0 -1 6510
box -12 -8 32 272
use FILL  FILL_3__3183_
timestamp 1701859473
transform 1 0 310 0 1 8070
box -12 -8 32 272
use FILL  FILL_3__3184_
timestamp 1701859473
transform -1 0 550 0 1 8070
box -12 -8 32 272
use FILL  FILL_3__3185_
timestamp 1701859473
transform -1 0 90 0 -1 8590
box -12 -8 32 272
use FILL  FILL_3__3186_
timestamp 1701859473
transform -1 0 90 0 1 8070
box -12 -8 32 272
use FILL  FILL_3__3187_
timestamp 1701859473
transform 1 0 710 0 -1 9110
box -12 -8 32 272
use FILL  FILL_3__3188_
timestamp 1701859473
transform 1 0 930 0 -1 9110
box -12 -8 32 272
use FILL  FILL_3__3189_
timestamp 1701859473
transform 1 0 2110 0 -1 9630
box -12 -8 32 272
use FILL  FILL_3__3190_
timestamp 1701859473
transform 1 0 2350 0 1 9110
box -12 -8 32 272
use FILL  FILL_3__3191_
timestamp 1701859473
transform 1 0 1410 0 -1 9110
box -12 -8 32 272
use FILL  FILL_3__3192_
timestamp 1701859473
transform -1 0 1650 0 -1 9110
box -12 -8 32 272
use FILL  FILL_3__3324_
timestamp 1701859473
transform 1 0 5590 0 1 8070
box -12 -8 32 272
use FILL  FILL_3__3325_
timestamp 1701859473
transform -1 0 6310 0 1 8070
box -12 -8 32 272
use FILL  FILL_3__3326_
timestamp 1701859473
transform -1 0 6210 0 -1 8070
box -12 -8 32 272
use FILL  FILL_3__3327_
timestamp 1701859473
transform -1 0 6170 0 -1 8590
box -12 -8 32 272
use FILL  FILL_3__3328_
timestamp 1701859473
transform -1 0 6070 0 1 8070
box -12 -8 32 272
use FILL  FILL_3__3329_
timestamp 1701859473
transform 1 0 5830 0 1 8070
box -12 -8 32 272
use FILL  FILL_3__3330_
timestamp 1701859473
transform -1 0 7010 0 1 8590
box -12 -8 32 272
use FILL  FILL_3__3331_
timestamp 1701859473
transform 1 0 7290 0 -1 8590
box -12 -8 32 272
use FILL  FILL_3__3332_
timestamp 1701859473
transform 1 0 7010 0 -1 8590
box -12 -8 32 272
use FILL  FILL_3__3333_
timestamp 1701859473
transform 1 0 10210 0 1 8590
box -12 -8 32 272
use FILL  FILL_3__3334_
timestamp 1701859473
transform 1 0 9330 0 1 8590
box -12 -8 32 272
use FILL  FILL_3__3335_
timestamp 1701859473
transform 1 0 7870 0 -1 10150
box -12 -8 32 272
use FILL  FILL_3__3336_
timestamp 1701859473
transform -1 0 6710 0 1 9630
box -12 -8 32 272
use FILL  FILL_3__3337_
timestamp 1701859473
transform -1 0 6230 0 1 9630
box -12 -8 32 272
use FILL  FILL_3__3338_
timestamp 1701859473
transform 1 0 7190 0 -1 10150
box -12 -8 32 272
use FILL  FILL_3__3339_
timestamp 1701859473
transform -1 0 8070 0 1 10150
box -12 -8 32 272
use FILL  FILL_3__3340_
timestamp 1701859473
transform 1 0 7830 0 1 10150
box -12 -8 32 272
use FILL  FILL_3__3341_
timestamp 1701859473
transform 1 0 7590 0 1 10150
box -12 -8 32 272
use FILL  FILL_3__3342_
timestamp 1701859473
transform 1 0 6810 0 -1 11190
box -12 -8 32 272
use FILL  FILL_3__3343_
timestamp 1701859473
transform -1 0 7410 0 -1 10150
box -12 -8 32 272
use FILL  FILL_3__3344_
timestamp 1701859473
transform 1 0 7630 0 -1 10150
box -12 -8 32 272
use FILL  FILL_3__3345_
timestamp 1701859473
transform -1 0 9010 0 1 9630
box -12 -8 32 272
use FILL  FILL_3__3346_
timestamp 1701859473
transform 1 0 8530 0 1 10150
box -12 -8 32 272
use FILL  FILL_3__3347_
timestamp 1701859473
transform -1 0 8310 0 1 10150
box -12 -8 32 272
use FILL  FILL_3__3348_
timestamp 1701859473
transform 1 0 9130 0 -1 10670
box -12 -8 32 272
use FILL  FILL_3__3349_
timestamp 1701859473
transform 1 0 7870 0 1 9630
box -12 -8 32 272
use FILL  FILL_3__3350_
timestamp 1701859473
transform 1 0 7570 0 -1 8590
box -12 -8 32 272
use FILL  FILL_3__3351_
timestamp 1701859473
transform -1 0 7750 0 1 8590
box -12 -8 32 272
use FILL  FILL_3__3352_
timestamp 1701859473
transform -1 0 8210 0 -1 9110
box -12 -8 32 272
use FILL  FILL_3__3353_
timestamp 1701859473
transform 1 0 8090 0 -1 10150
box -12 -8 32 272
use FILL  FILL_3__3354_
timestamp 1701859473
transform 1 0 7770 0 -1 10670
box -12 -8 32 272
use FILL  FILL_3__3355_
timestamp 1701859473
transform -1 0 7550 0 -1 10670
box -12 -8 32 272
use FILL  FILL_3__3356_
timestamp 1701859473
transform 1 0 7330 0 -1 10670
box -12 -8 32 272
use FILL  FILL_3__3357_
timestamp 1701859473
transform 1 0 7150 0 1 10670
box -12 -8 32 272
use FILL  FILL_3__3358_
timestamp 1701859473
transform 1 0 7410 0 1 10670
box -12 -8 32 272
use FILL  FILL_3__3359_
timestamp 1701859473
transform 1 0 7650 0 1 10670
box -12 -8 32 272
use FILL  FILL_3__3360_
timestamp 1701859473
transform -1 0 7910 0 1 10670
box -12 -8 32 272
use FILL  FILL_3__3361_
timestamp 1701859473
transform 1 0 8930 0 -1 10670
box -12 -8 32 272
use FILL  FILL_3__3362_
timestamp 1701859473
transform 1 0 7990 0 -1 10670
box -12 -8 32 272
use FILL  FILL_3__3363_
timestamp 1701859473
transform 1 0 8110 0 1 10670
box -12 -8 32 272
use FILL  FILL_3__3364_
timestamp 1701859473
transform 1 0 7950 0 -1 11190
box -12 -8 32 272
use FILL  FILL_3__3365_
timestamp 1701859473
transform -1 0 7490 0 -1 11190
box -12 -8 32 272
use FILL  FILL_3__3366_
timestamp 1701859473
transform 1 0 7010 0 -1 11190
box -12 -8 32 272
use FILL  FILL_3__3367_
timestamp 1701859473
transform 1 0 6890 0 1 10670
box -12 -8 32 272
use FILL  FILL_3__3368_
timestamp 1701859473
transform 1 0 7230 0 -1 11190
box -12 -8 32 272
use FILL  FILL_3__3369_
timestamp 1701859473
transform 1 0 7710 0 -1 11190
box -12 -8 32 272
use FILL  FILL_3__3370_
timestamp 1701859473
transform 1 0 8230 0 -1 10670
box -12 -8 32 272
use FILL  FILL_3__3371_
timestamp 1701859473
transform 1 0 8330 0 1 10670
box -12 -8 32 272
use FILL  FILL_3__3372_
timestamp 1701859473
transform 1 0 9510 0 1 10670
box -12 -8 32 272
use FILL  FILL_3__3373_
timestamp 1701859473
transform -1 0 6610 0 -1 11190
box -12 -8 32 272
use FILL  FILL_3__3374_
timestamp 1701859473
transform 1 0 5710 0 1 10670
box -12 -8 32 272
use FILL  FILL_3__3375_
timestamp 1701859473
transform -1 0 5970 0 1 10670
box -12 -8 32 272
use FILL  FILL_3__3376_
timestamp 1701859473
transform -1 0 6190 0 1 10670
box -12 -8 32 272
use FILL  FILL_3__3377_
timestamp 1701859473
transform 1 0 6430 0 1 10670
box -12 -8 32 272
use FILL  FILL_3__3378_
timestamp 1701859473
transform 1 0 6370 0 -1 11190
box -12 -8 32 272
use FILL  FILL_3__3379_
timestamp 1701859473
transform 1 0 8690 0 -1 10670
box -12 -8 32 272
use FILL  FILL_3__3380_
timestamp 1701859473
transform 1 0 8810 0 1 10670
box -12 -8 32 272
use FILL  FILL_3__3381_
timestamp 1701859473
transform -1 0 6690 0 1 10670
box -12 -8 32 272
use FILL  FILL_3__3382_
timestamp 1701859473
transform 1 0 6150 0 -1 10670
box -12 -8 32 272
use FILL  FILL_3__3383_
timestamp 1701859473
transform -1 0 6410 0 -1 10670
box -12 -8 32 272
use FILL  FILL_3__3384_
timestamp 1701859473
transform -1 0 6850 0 -1 10670
box -12 -8 32 272
use FILL  FILL_3__3385_
timestamp 1701859473
transform 1 0 6610 0 -1 10670
box -12 -8 32 272
use FILL  FILL_3__3386_
timestamp 1701859473
transform 1 0 7090 0 -1 10670
box -12 -8 32 272
use FILL  FILL_3__3387_
timestamp 1701859473
transform 1 0 8450 0 -1 10670
box -12 -8 32 272
use FILL  FILL_3__3388_
timestamp 1701859473
transform 1 0 8570 0 1 10670
box -12 -8 32 272
use FILL  FILL_3__3389_
timestamp 1701859473
transform 1 0 10230 0 -1 10670
box -12 -8 32 272
use FILL  FILL_3__3390_
timestamp 1701859473
transform 1 0 9790 0 -1 10670
box -12 -8 32 272
use FILL  FILL_3__3391_
timestamp 1701859473
transform 1 0 9990 0 -1 10670
box -12 -8 32 272
use FILL  FILL_3__3392_
timestamp 1701859473
transform 1 0 10450 0 -1 10670
box -12 -8 32 272
use FILL  FILL_3__3393_
timestamp 1701859473
transform -1 0 11190 0 -1 10150
box -12 -8 32 272
use FILL  FILL_3__3394_
timestamp 1701859473
transform 1 0 7370 0 1 10150
box -12 -8 32 272
use FILL  FILL_3__3395_
timestamp 1701859473
transform 1 0 6430 0 1 10150
box -12 -8 32 272
use FILL  FILL_3__3396_
timestamp 1701859473
transform -1 0 6690 0 1 10150
box -12 -8 32 272
use FILL  FILL_3__3397_
timestamp 1701859473
transform -1 0 7010 0 -1 10150
box -12 -8 32 272
use FILL  FILL_3__3398_
timestamp 1701859473
transform 1 0 6290 0 -1 10150
box -12 -8 32 272
use FILL  FILL_3__3399_
timestamp 1701859473
transform -1 0 6770 0 -1 10150
box -12 -8 32 272
use FILL  FILL_3__3400_
timestamp 1701859473
transform -1 0 6950 0 1 10150
box -12 -8 32 272
use FILL  FILL_3__3401_
timestamp 1701859473
transform 1 0 7130 0 1 10150
box -12 -8 32 272
use FILL  FILL_3__3402_
timestamp 1701859473
transform -1 0 9070 0 1 10150
box -12 -8 32 272
use FILL  FILL_3__3403_
timestamp 1701859473
transform 1 0 9510 0 1 10150
box -12 -8 32 272
use FILL  FILL_3__3404_
timestamp 1701859473
transform -1 0 5770 0 1 9630
box -12 -8 32 272
use FILL  FILL_3__3405_
timestamp 1701859473
transform -1 0 6050 0 -1 10150
box -12 -8 32 272
use FILL  FILL_3__3406_
timestamp 1701859473
transform 1 0 6410 0 -1 9630
box -12 -8 32 272
use FILL  FILL_3__3407_
timestamp 1701859473
transform -1 0 6630 0 -1 9630
box -12 -8 32 272
use FILL  FILL_3__3408_
timestamp 1701859473
transform 1 0 6890 0 1 9630
box -12 -8 32 272
use FILL  FILL_3__3409_
timestamp 1701859473
transform -1 0 6510 0 -1 10150
box -12 -8 32 272
use FILL  FILL_3__3410_
timestamp 1701859473
transform 1 0 9250 0 -1 10150
box -12 -8 32 272
use FILL  FILL_3__3411_
timestamp 1701859473
transform 1 0 9270 0 1 10150
box -12 -8 32 272
use FILL  FILL_3__3412_
timestamp 1701859473
transform 1 0 9990 0 1 10150
box -12 -8 32 272
use FILL  FILL_3__3413_
timestamp 1701859473
transform -1 0 6010 0 1 9630
box -12 -8 32 272
use FILL  FILL_3__3414_
timestamp 1701859473
transform 1 0 8150 0 1 9110
box -12 -8 32 272
use FILL  FILL_3__3415_
timestamp 1701859473
transform 1 0 6430 0 1 9630
box -12 -8 32 272
use FILL  FILL_3__3416_
timestamp 1701859473
transform 1 0 7270 0 1 8590
box -12 -8 32 272
use FILL  FILL_3__3417_
timestamp 1701859473
transform 1 0 7350 0 -1 9110
box -12 -8 32 272
use FILL  FILL_3__3418_
timestamp 1701859473
transform -1 0 7490 0 -1 9630
box -12 -8 32 272
use FILL  FILL_3__3419_
timestamp 1701859473
transform 1 0 7250 0 -1 9630
box -12 -8 32 272
use FILL  FILL_3__3420_
timestamp 1701859473
transform -1 0 6830 0 -1 9630
box -12 -8 32 272
use FILL  FILL_3__3421_
timestamp 1701859473
transform -1 0 7050 0 -1 9630
box -12 -8 32 272
use FILL  FILL_3__3422_
timestamp 1701859473
transform -1 0 7150 0 1 9630
box -12 -8 32 272
use FILL  FILL_3__3423_
timestamp 1701859473
transform -1 0 8210 0 -1 9630
box -12 -8 32 272
use FILL  FILL_3__3424_
timestamp 1701859473
transform -1 0 7730 0 -1 9630
box -12 -8 32 272
use FILL  FILL_3__3425_
timestamp 1701859473
transform -1 0 7390 0 1 9630
box -12 -8 32 272
use FILL  FILL_3__3426_
timestamp 1701859473
transform -1 0 9030 0 -1 10150
box -12 -8 32 272
use FILL  FILL_3__3427_
timestamp 1701859473
transform 1 0 8790 0 -1 10150
box -12 -8 32 272
use FILL  FILL_3__3428_
timestamp 1701859473
transform 1 0 7470 0 1 8590
box -12 -8 32 272
use FILL  FILL_3__3429_
timestamp 1701859473
transform 1 0 7550 0 -1 9110
box -12 -8 32 272
use FILL  FILL_3__3430_
timestamp 1701859473
transform -1 0 7770 0 -1 9110
box -12 -8 32 272
use FILL  FILL_3__3431_
timestamp 1701859473
transform 1 0 7690 0 1 9110
box -12 -8 32 272
use FILL  FILL_3__3432_
timestamp 1701859473
transform 1 0 7930 0 1 9110
box -12 -8 32 272
use FILL  FILL_3__3433_
timestamp 1701859473
transform -1 0 7970 0 -1 9630
box -12 -8 32 272
use FILL  FILL_3__3434_
timestamp 1701859473
transform 1 0 7610 0 1 9630
box -12 -8 32 272
use FILL  FILL_3__3435_
timestamp 1701859473
transform 1 0 10230 0 1 10150
box -12 -8 32 272
use FILL  FILL_3__3436_
timestamp 1701859473
transform -1 0 10230 0 -1 10150
box -12 -8 32 272
use FILL  FILL_3__3437_
timestamp 1701859473
transform 1 0 10670 0 1 10150
box -12 -8 32 272
use FILL  FILL_3__3438_
timestamp 1701859473
transform 1 0 10450 0 1 10150
box -12 -8 32 272
use FILL  FILL_3__3439_
timestamp 1701859473
transform 1 0 10890 0 1 10150
box -12 -8 32 272
use FILL  FILL_3__3440_
timestamp 1701859473
transform -1 0 10710 0 -1 10150
box -12 -8 32 272
use FILL  FILL_3__3441_
timestamp 1701859473
transform -1 0 10570 0 1 9630
box -12 -8 32 272
use FILL  FILL_3__3442_
timestamp 1701859473
transform -1 0 10450 0 -1 10150
box -12 -8 32 272
use FILL  FILL_3__3443_
timestamp 1701859473
transform -1 0 11010 0 1 9630
box -12 -8 32 272
use FILL  FILL_3__3444_
timestamp 1701859473
transform -1 0 8410 0 -1 9630
box -12 -8 32 272
use FILL  FILL_3__3445_
timestamp 1701859473
transform -1 0 8110 0 1 9630
box -12 -8 32 272
use FILL  FILL_3__3446_
timestamp 1701859473
transform 1 0 8550 0 1 9630
box -12 -8 32 272
use FILL  FILL_3__3447_
timestamp 1701859473
transform 1 0 8330 0 1 9630
box -12 -8 32 272
use FILL  FILL_3__3448_
timestamp 1701859473
transform -1 0 8770 0 1 9630
box -12 -8 32 272
use FILL  FILL_3__3449_
timestamp 1701859473
transform -1 0 9810 0 1 10150
box -12 -8 32 272
use FILL  FILL_3__3450_
timestamp 1701859473
transform -1 0 9770 0 -1 10150
box -12 -8 32 272
use FILL  FILL_3__3451_
timestamp 1701859473
transform 1 0 9490 0 -1 10150
box -12 -8 32 272
use FILL  FILL_3__3452_
timestamp 1701859473
transform -1 0 9230 0 1 9630
box -12 -8 32 272
use FILL  FILL_3__3453_
timestamp 1701859473
transform -1 0 9990 0 -1 10150
box -12 -8 32 272
use FILL  FILL_3__3454_
timestamp 1701859473
transform 1 0 9430 0 1 9630
box -12 -8 32 272
use FILL  FILL_3__3455_
timestamp 1701859473
transform 1 0 9650 0 1 9630
box -12 -8 32 272
use FILL  FILL_3__3456_
timestamp 1701859473
transform -1 0 10350 0 1 9630
box -12 -8 32 272
use FILL  FILL_3__3457_
timestamp 1701859473
transform -1 0 9890 0 1 9630
box -12 -8 32 272
use FILL  FILL_3__3458_
timestamp 1701859473
transform -1 0 10130 0 1 9630
box -12 -8 32 272
use FILL  FILL_3__3459_
timestamp 1701859473
transform -1 0 10270 0 -1 9630
box -12 -8 32 272
use FILL  FILL_3__3460_
timestamp 1701859473
transform 1 0 10930 0 -1 10150
box -12 -8 32 272
use FILL  FILL_3__3461_
timestamp 1701859473
transform -1 0 11170 0 -1 9630
box -12 -8 32 272
use FILL  FILL_3__3462_
timestamp 1701859473
transform -1 0 10710 0 -1 9630
box -12 -8 32 272
use FILL  FILL_3__3463_
timestamp 1701859473
transform 1 0 10390 0 -1 11190
box -12 -8 32 272
use FILL  FILL_3__3464_
timestamp 1701859473
transform 1 0 9730 0 -1 11190
box -12 -8 32 272
use FILL  FILL_3__3465_
timestamp 1701859473
transform 1 0 9970 0 -1 11190
box -12 -8 32 272
use FILL  FILL_3__3466_
timestamp 1701859473
transform 1 0 10150 0 -1 11190
box -12 -8 32 272
use FILL  FILL_3__3467_
timestamp 1701859473
transform -1 0 11130 0 1 10670
box -12 -8 32 272
use FILL  FILL_3__3468_
timestamp 1701859473
transform 1 0 10630 0 1 10670
box -12 -8 32 272
use FILL  FILL_3__3469_
timestamp 1701859473
transform 1 0 9350 0 -1 10670
box -12 -8 32 272
use FILL  FILL_3__3470_
timestamp 1701859473
transform 1 0 9590 0 -1 10670
box -12 -8 32 272
use FILL  FILL_3__3471_
timestamp 1701859473
transform 1 0 9730 0 1 10670
box -12 -8 32 272
use FILL  FILL_3__3472_
timestamp 1701859473
transform -1 0 9990 0 1 10670
box -12 -8 32 272
use FILL  FILL_3__3473_
timestamp 1701859473
transform 1 0 8610 0 -1 11190
box -12 -8 32 272
use FILL  FILL_3__3474_
timestamp 1701859473
transform 1 0 8170 0 -1 11190
box -12 -8 32 272
use FILL  FILL_3__3475_
timestamp 1701859473
transform 1 0 8410 0 -1 11190
box -12 -8 32 272
use FILL  FILL_3__3476_
timestamp 1701859473
transform -1 0 8850 0 -1 11190
box -12 -8 32 272
use FILL  FILL_3__3477_
timestamp 1701859473
transform 1 0 9070 0 -1 11190
box -12 -8 32 272
use FILL  FILL_3__3478_
timestamp 1701859473
transform 1 0 9050 0 1 10670
box -12 -8 32 272
use FILL  FILL_3__3479_
timestamp 1701859473
transform 1 0 8330 0 -1 10150
box -12 -8 32 272
use FILL  FILL_3__3480_
timestamp 1701859473
transform -1 0 8590 0 -1 10150
box -12 -8 32 272
use FILL  FILL_3__3481_
timestamp 1701859473
transform -1 0 8370 0 1 9110
box -12 -8 32 272
use FILL  FILL_3__3482_
timestamp 1701859473
transform -1 0 8590 0 1 9110
box -12 -8 32 272
use FILL  FILL_3__3483_
timestamp 1701859473
transform 1 0 8770 0 1 10150
box -12 -8 32 272
use FILL  FILL_3__3484_
timestamp 1701859473
transform -1 0 10070 0 -1 9630
box -12 -8 32 272
use FILL  FILL_3__3485_
timestamp 1701859473
transform 1 0 11090 0 1 10150
box -12 -8 32 272
use FILL  FILL_3__3486_
timestamp 1701859473
transform 1 0 10430 0 1 9110
box -12 -8 32 272
use FILL  FILL_3__3487_
timestamp 1701859473
transform 1 0 10470 0 -1 9630
box -12 -8 32 272
use FILL  FILL_3__3488_
timestamp 1701859473
transform -1 0 10770 0 1 9630
box -12 -8 32 272
use FILL  FILL_3__3489_
timestamp 1701859473
transform 1 0 10610 0 -1 11190
box -12 -8 32 272
use FILL  FILL_3__3490_
timestamp 1701859473
transform 1 0 11070 0 -1 11190
box -12 -8 32 272
use FILL  FILL_3__3491_
timestamp 1701859473
transform -1 0 10870 0 -1 11190
box -12 -8 32 272
use FILL  FILL_3__3492_
timestamp 1701859473
transform -1 0 10430 0 1 10670
box -12 -8 32 272
use FILL  FILL_3__3493_
timestamp 1701859473
transform -1 0 10210 0 1 10670
box -12 -8 32 272
use FILL  FILL_3__3494_
timestamp 1701859473
transform 1 0 9310 0 1 10670
box -12 -8 32 272
use FILL  FILL_3__3495_
timestamp 1701859473
transform -1 0 9510 0 -1 11190
box -12 -8 32 272
use FILL  FILL_3__3496_
timestamp 1701859473
transform 1 0 9270 0 -1 11190
box -12 -8 32 272
use FILL  FILL_3__3497_
timestamp 1701859473
transform -1 0 9370 0 -1 9630
box -12 -8 32 272
use FILL  FILL_3__3498_
timestamp 1701859473
transform -1 0 8870 0 1 9110
box -12 -8 32 272
use FILL  FILL_3__3499_
timestamp 1701859473
transform 1 0 8390 0 -1 9110
box -12 -8 32 272
use FILL  FILL_3__3500_
timestamp 1701859473
transform 1 0 9770 0 1 9110
box -12 -8 32 272
use FILL  FILL_3__3501_
timestamp 1701859473
transform -1 0 10010 0 1 9110
box -12 -8 32 272
use FILL  FILL_3__3502_
timestamp 1701859473
transform -1 0 8270 0 -1 8590
box -12 -8 32 272
use FILL  FILL_3__3503_
timestamp 1701859473
transform -1 0 8650 0 -1 9630
box -12 -8 32 272
use FILL  FILL_3__3504_
timestamp 1701859473
transform 1 0 8870 0 -1 9630
box -12 -8 32 272
use FILL  FILL_3__3505_
timestamp 1701859473
transform -1 0 9130 0 -1 9630
box -12 -8 32 272
use FILL  FILL_3__3506_
timestamp 1701859473
transform -1 0 8650 0 1 8590
box -12 -8 32 272
use FILL  FILL_3__3507_
timestamp 1701859473
transform 1 0 10730 0 -1 9110
box -12 -8 32 272
use FILL  FILL_3__3508_
timestamp 1701859473
transform 1 0 10490 0 -1 9110
box -12 -8 32 272
use FILL  FILL_3__3509_
timestamp 1701859473
transform 1 0 8430 0 1 8590
box -12 -8 32 272
use FILL  FILL_3__3510_
timestamp 1701859473
transform -1 0 8890 0 1 8590
box -12 -8 32 272
use FILL  FILL_3__3511_
timestamp 1701859473
transform 1 0 9950 0 -1 270
box -12 -8 32 272
use FILL  FILL_3__3512_
timestamp 1701859473
transform 1 0 10950 0 -1 9110
box -12 -8 32 272
use FILL  FILL_3__3513_
timestamp 1701859473
transform 1 0 10930 0 -1 9630
box -12 -8 32 272
use FILL  FILL_3__3514_
timestamp 1701859473
transform 1 0 10890 0 1 10670
box -12 -8 32 272
use FILL  FILL_3__3515_
timestamp 1701859473
transform -1 0 10690 0 -1 10670
box -12 -8 32 272
use FILL  FILL_3__3516_
timestamp 1701859473
transform 1 0 10910 0 -1 10670
box -12 -8 32 272
use FILL  FILL_3__3517_
timestamp 1701859473
transform 1 0 9590 0 -1 9630
box -12 -8 32 272
use FILL  FILL_3__3518_
timestamp 1701859473
transform 1 0 9810 0 -1 9630
box -12 -8 32 272
use FILL  FILL_3__3519_
timestamp 1701859473
transform 1 0 9090 0 1 9110
box -12 -8 32 272
use FILL  FILL_3__3520_
timestamp 1701859473
transform -1 0 9330 0 1 9110
box -12 -8 32 272
use FILL  FILL_3__3521_
timestamp 1701859473
transform 1 0 6570 0 1 8590
box -12 -8 32 272
use FILL  FILL_3__3522_
timestamp 1701859473
transform 1 0 7970 0 -1 9110
box -12 -8 32 272
use FILL  FILL_3__3523_
timestamp 1701859473
transform 1 0 6770 0 1 8590
box -12 -8 32 272
use FILL  FILL_3__3524_
timestamp 1701859473
transform 1 0 7490 0 1 9110
box -12 -8 32 272
use FILL  FILL_3__3525_
timestamp 1701859473
transform 1 0 7030 0 1 9110
box -12 -8 32 272
use FILL  FILL_3__3526_
timestamp 1701859473
transform -1 0 7270 0 1 9110
box -12 -8 32 272
use FILL  FILL_3__3539_
timestamp 1701859473
transform 1 0 11130 0 -1 7030
box -12 -8 32 272
use FILL  FILL_3__3540_
timestamp 1701859473
transform 1 0 4630 0 1 10670
box -12 -8 32 272
use FILL  FILL_3__3541_
timestamp 1701859473
transform -1 0 90 0 1 5990
box -12 -8 32 272
use FILL  FILL_3__3542_
timestamp 1701859473
transform -1 0 90 0 -1 8070
box -12 -8 32 272
use FILL  FILL_3__3543_
timestamp 1701859473
transform -1 0 90 0 1 8590
box -12 -8 32 272
use FILL  FILL_3__3544_
timestamp 1701859473
transform -1 0 90 0 1 9110
box -12 -8 32 272
use FILL  FILL_3__3545_
timestamp 1701859473
transform -1 0 1930 0 -1 11190
box -12 -8 32 272
use FILL  FILL_3__3546_
timestamp 1701859473
transform -1 0 550 0 1 9110
box -12 -8 32 272
use FILL  FILL_3__3547_
timestamp 1701859473
transform 1 0 4670 0 -1 11190
box -12 -8 32 272
use FILL  FILL_3__3548_
timestamp 1701859473
transform 1 0 5270 0 1 10670
box -12 -8 32 272
use FILL  FILL_3__3549_
timestamp 1701859473
transform -1 0 4270 0 -1 11190
box -12 -8 32 272
use FILL  FILL_3__3550_
timestamp 1701859473
transform -1 0 5110 0 -1 11190
box -12 -8 32 272
use FILL  FILL_3__3551_
timestamp 1701859473
transform 1 0 5510 0 -1 11190
box -12 -8 32 272
use FILL  FILL_3__3552_
timestamp 1701859473
transform 1 0 5290 0 -1 11190
box -12 -8 32 272
use FILL  FILL_3__3553_
timestamp 1701859473
transform -1 0 90 0 -1 5990
box -12 -8 32 272
use FILL  FILL_3__3554_
timestamp 1701859473
transform -1 0 290 0 1 7030
box -12 -8 32 272
use FILL  FILL_3__3555_
timestamp 1701859473
transform -1 0 5070 0 1 10670
box -12 -8 32 272
use FILL  FILL_3__3556_
timestamp 1701859473
transform 1 0 6210 0 1 10150
box -12 -8 32 272
use FILL  FILL_3__3557_
timestamp 1701859473
transform -1 0 5750 0 -1 11190
box -12 -8 32 272
use FILL  FILL_3__3558_
timestamp 1701859473
transform 1 0 6150 0 -1 11190
box -12 -8 32 272
use FILL  FILL_3__3559_
timestamp 1701859473
transform -1 0 4810 0 -1 10670
box -12 -8 32 272
use FILL  FILL_3__3560_
timestamp 1701859473
transform 1 0 5490 0 1 10670
box -12 -8 32 272
use FILL  FILL_3__3561_
timestamp 1701859473
transform 1 0 5930 0 -1 11190
box -12 -8 32 272
use FILL  FILL_3__3562_
timestamp 1701859473
transform 1 0 5730 0 1 10150
box -12 -8 32 272
use FILL  FILL_3__3563_
timestamp 1701859473
transform 1 0 5190 0 1 3390
box -12 -8 32 272
use FILL  FILL_3_BUFX2_insert0
timestamp 1701859473
transform 1 0 5810 0 -1 10150
box -12 -8 32 272
use FILL  FILL_3_BUFX2_insert1
timestamp 1701859473
transform 1 0 6570 0 1 2350
box -12 -8 32 272
use FILL  FILL_3_BUFX2_insert2
timestamp 1701859473
transform 1 0 5410 0 -1 1830
box -12 -8 32 272
use FILL  FILL_3_BUFX2_insert3
timestamp 1701859473
transform -1 0 550 0 -1 5470
box -12 -8 32 272
use FILL  FILL_3_BUFX2_insert4
timestamp 1701859473
transform 1 0 3290 0 1 4950
box -12 -8 32 272
use FILL  FILL_3_BUFX2_insert5
timestamp 1701859473
transform 1 0 1350 0 -1 1830
box -12 -8 32 272
use FILL  FILL_3_BUFX2_insert6
timestamp 1701859473
transform -1 0 90 0 -1 11190
box -12 -8 32 272
use FILL  FILL_3_BUFX2_insert7
timestamp 1701859473
transform 1 0 1650 0 1 10670
box -12 -8 32 272
use FILL  FILL_3_BUFX2_insert8
timestamp 1701859473
transform 1 0 1610 0 1 1830
box -12 -8 32 272
use FILL  FILL_3_BUFX2_insert9
timestamp 1701859473
transform 1 0 1910 0 -1 3910
box -12 -8 32 272
use FILL  FILL_3_BUFX2_insert10
timestamp 1701859473
transform 1 0 1730 0 -1 4430
box -12 -8 32 272
use FILL  FILL_3_BUFX2_insert11
timestamp 1701859473
transform -1 0 1710 0 -1 3910
box -12 -8 32 272
use FILL  FILL_3_BUFX2_insert12
timestamp 1701859473
transform -1 0 1490 0 -1 3910
box -12 -8 32 272
use FILL  FILL_3_BUFX2_insert13
timestamp 1701859473
transform -1 0 1390 0 -1 1310
box -12 -8 32 272
use FILL  FILL_3_BUFX2_insert14
timestamp 1701859473
transform -1 0 3630 0 1 3390
box -12 -8 32 272
use FILL  FILL_3_BUFX2_insert15
timestamp 1701859473
transform 1 0 4510 0 -1 5470
box -12 -8 32 272
use FILL  FILL_3_BUFX2_insert16
timestamp 1701859473
transform 1 0 1310 0 -1 4950
box -12 -8 32 272
use FILL  FILL_3_BUFX2_insert17
timestamp 1701859473
transform 1 0 3590 0 1 1310
box -12 -8 32 272
use FILL  FILL_3_BUFX2_insert18
timestamp 1701859473
transform -1 0 9730 0 1 2350
box -12 -8 32 272
use FILL  FILL_3_BUFX2_insert19
timestamp 1701859473
transform -1 0 8470 0 -1 790
box -12 -8 32 272
use FILL  FILL_3_BUFX2_insert20
timestamp 1701859473
transform 1 0 9930 0 1 2350
box -12 -8 32 272
use FILL  FILL_3_BUFX2_insert21
timestamp 1701859473
transform -1 0 7770 0 -1 1310
box -12 -8 32 272
use FILL  FILL_3_BUFX2_insert22
timestamp 1701859473
transform -1 0 3170 0 -1 2870
box -12 -8 32 272
use FILL  FILL_3_BUFX2_insert23
timestamp 1701859473
transform -1 0 2710 0 -1 4950
box -12 -8 32 272
use FILL  FILL_3_BUFX2_insert24
timestamp 1701859473
transform -1 0 3610 0 -1 4430
box -12 -8 32 272
use FILL  FILL_3_BUFX2_insert25
timestamp 1701859473
transform 1 0 4350 0 1 4430
box -12 -8 32 272
use FILL  FILL_3_BUFX2_insert26
timestamp 1701859473
transform 1 0 4170 0 1 2870
box -12 -8 32 272
use FILL  FILL_3_BUFX2_insert27
timestamp 1701859473
transform 1 0 9570 0 1 4950
box -12 -8 32 272
use FILL  FILL_3_BUFX2_insert28
timestamp 1701859473
transform -1 0 7450 0 -1 5990
box -12 -8 32 272
use FILL  FILL_3_BUFX2_insert29
timestamp 1701859473
transform -1 0 1250 0 1 6510
box -12 -8 32 272
use FILL  FILL_3_BUFX2_insert30
timestamp 1701859473
transform -1 0 8750 0 -1 3910
box -12 -8 32 272
use FILL  FILL_3_BUFX2_insert31
timestamp 1701859473
transform -1 0 9530 0 1 3910
box -12 -8 32 272
use FILL  FILL_3_BUFX2_insert32
timestamp 1701859473
transform 1 0 5830 0 -1 3910
box -12 -8 32 272
use FILL  FILL_3_BUFX2_insert33
timestamp 1701859473
transform -1 0 9510 0 -1 4950
box -12 -8 32 272
use FILL  FILL_3_BUFX2_insert34
timestamp 1701859473
transform 1 0 5170 0 1 8590
box -12 -8 32 272
use FILL  FILL_3_BUFX2_insert35
timestamp 1701859473
transform -1 0 5930 0 1 7550
box -12 -8 32 272
use FILL  FILL_3_BUFX2_insert36
timestamp 1701859473
transform -1 0 1170 0 1 8590
box -12 -8 32 272
use FILL  FILL_3_BUFX2_insert37
timestamp 1701859473
transform -1 0 9550 0 1 8590
box -12 -8 32 272
use FILL  FILL_3_BUFX2_insert49
timestamp 1701859473
transform -1 0 3010 0 1 6510
box -12 -8 32 272
use FILL  FILL_3_BUFX2_insert50
timestamp 1701859473
transform 1 0 2310 0 -1 8590
box -12 -8 32 272
use FILL  FILL_3_BUFX2_insert51
timestamp 1701859473
transform 1 0 3170 0 -1 8590
box -12 -8 32 272
use FILL  FILL_3_BUFX2_insert52
timestamp 1701859473
transform 1 0 3350 0 1 5470
box -12 -8 32 272
use FILL  FILL_3_BUFX2_insert53
timestamp 1701859473
transform -1 0 11190 0 1 9110
box -12 -8 32 272
use FILL  FILL_3_BUFX2_insert54
timestamp 1701859473
transform -1 0 9130 0 1 8590
box -12 -8 32 272
use FILL  FILL_3_BUFX2_insert55
timestamp 1701859473
transform -1 0 9570 0 1 9110
box -12 -8 32 272
use FILL  FILL_3_BUFX2_insert56
timestamp 1701859473
transform -1 0 10230 0 1 9110
box -12 -8 32 272
use FILL  FILL_3_BUFX2_insert57
timestamp 1701859473
transform -1 0 11190 0 -1 2350
box -12 -8 32 272
use FILL  FILL_3_BUFX2_insert58
timestamp 1701859473
transform -1 0 8930 0 1 2870
box -12 -8 32 272
use FILL  FILL_3_BUFX2_insert59
timestamp 1701859473
transform -1 0 7510 0 1 1830
box -12 -8 32 272
use FILL  FILL_3_BUFX2_insert60
timestamp 1701859473
transform 1 0 10850 0 1 1830
box -12 -8 32 272
use FILL  FILL_3_BUFX2_insert61
timestamp 1701859473
transform -1 0 11130 0 1 2870
box -12 -8 32 272
use FILL  FILL_3_BUFX2_insert62
timestamp 1701859473
transform 1 0 2170 0 1 3910
box -12 -8 32 272
use FILL  FILL_3_BUFX2_insert63
timestamp 1701859473
transform 1 0 2090 0 1 3390
box -12 -8 32 272
use FILL  FILL_3_BUFX2_insert64
timestamp 1701859473
transform -1 0 1750 0 1 3910
box -12 -8 32 272
use FILL  FILL_3_BUFX2_insert65
timestamp 1701859473
transform -1 0 1690 0 1 3390
box -12 -8 32 272
use FILL  FILL_3_BUFX2_insert66
timestamp 1701859473
transform -1 0 4270 0 1 1310
box -12 -8 32 272
use FILL  FILL_3_BUFX2_insert67
timestamp 1701859473
transform -1 0 3570 0 -1 10150
box -12 -8 32 272
use FILL  FILL_3_BUFX2_insert68
timestamp 1701859473
transform -1 0 7130 0 1 2870
box -12 -8 32 272
use FILL  FILL_3_BUFX2_insert69
timestamp 1701859473
transform -1 0 5610 0 -1 3390
box -12 -8 32 272
use FILL  FILL_3_BUFX2_insert70
timestamp 1701859473
transform -1 0 3630 0 -1 1830
box -12 -8 32 272
use FILL  FILL_3_BUFX2_insert71
timestamp 1701859473
transform -1 0 7270 0 1 2350
box -12 -8 32 272
use FILL  FILL_3_BUFX2_insert72
timestamp 1701859473
transform -1 0 6450 0 1 1310
box -12 -8 32 272
use FILL  FILL_3_BUFX2_insert73
timestamp 1701859473
transform 1 0 3570 0 1 5470
box -12 -8 32 272
use FILL  FILL_3_BUFX2_insert74
timestamp 1701859473
transform 1 0 7530 0 -1 2350
box -12 -8 32 272
use FILL  FILL_3_BUFX2_insert75
timestamp 1701859473
transform 1 0 7550 0 1 2870
box -12 -8 32 272
use FILL  FILL_3_BUFX2_insert76
timestamp 1701859473
transform 1 0 7330 0 1 2870
box -12 -8 32 272
use FILL  FILL_3_BUFX2_insert77
timestamp 1701859473
transform -1 0 3390 0 -1 2870
box -12 -8 32 272
use FILL  FILL_3_BUFX2_insert78
timestamp 1701859473
transform 1 0 1890 0 -1 2870
box -12 -8 32 272
use FILL  FILL_3_BUFX2_insert79
timestamp 1701859473
transform -1 0 2130 0 -1 2870
box -12 -8 32 272
use FILL  FILL_3_BUFX2_insert80
timestamp 1701859473
transform 1 0 2370 0 1 4430
box -12 -8 32 272
use FILL  FILL_3_BUFX2_insert81
timestamp 1701859473
transform -1 0 1970 0 1 3910
box -12 -8 32 272
use FILL  FILL_3_BUFX2_insert82
timestamp 1701859473
transform -1 0 290 0 1 8590
box -12 -8 32 272
use FILL  FILL_3_BUFX2_insert83
timestamp 1701859473
transform 1 0 4170 0 -1 10150
box -12 -8 32 272
use FILL  FILL_3_BUFX2_insert84
timestamp 1701859473
transform 1 0 4130 0 -1 7550
box -12 -8 32 272
use FILL  FILL_3_BUFX2_insert85
timestamp 1701859473
transform -1 0 90 0 -1 6510
box -12 -8 32 272
use FILL  FILL_3_BUFX2_insert86
timestamp 1701859473
transform 1 0 1890 0 -1 10150
box -12 -8 32 272
use FILL  FILL_3_CLKBUF1_insert38
timestamp 1701859473
transform 1 0 2890 0 -1 7550
box -12 -8 32 272
use FILL  FILL_3_CLKBUF1_insert39
timestamp 1701859473
transform -1 0 4690 0 -1 6510
box -12 -8 32 272
use FILL  FILL_3_CLKBUF1_insert40
timestamp 1701859473
transform -1 0 990 0 -1 4950
box -12 -8 32 272
use FILL  FILL_3_CLKBUF1_insert41
timestamp 1701859473
transform -1 0 10650 0 -1 270
box -12 -8 32 272
use FILL  FILL_3_CLKBUF1_insert42
timestamp 1701859473
transform 1 0 9710 0 -1 4950
box -12 -8 32 272
use FILL  FILL_3_CLKBUF1_insert43
timestamp 1701859473
transform -1 0 11030 0 1 7030
box -12 -8 32 272
use FILL  FILL_3_CLKBUF1_insert44
timestamp 1701859473
transform -1 0 10770 0 1 4430
box -12 -8 32 272
use FILL  FILL_3_CLKBUF1_insert45
timestamp 1701859473
transform 1 0 5690 0 -1 6510
box -12 -8 32 272
use FILL  FILL_3_CLKBUF1_insert46
timestamp 1701859473
transform 1 0 4010 0 1 5990
box -12 -8 32 272
use FILL  FILL_3_CLKBUF1_insert47
timestamp 1701859473
transform -1 0 2130 0 1 7550
box -12 -8 32 272
use FILL  FILL_3_CLKBUF1_insert48
timestamp 1701859473
transform -1 0 10810 0 -1 7030
box -12 -8 32 272
use FILL  FILL_4__1668_
timestamp 1701859473
transform 1 0 6770 0 -1 3390
box -12 -8 32 272
use FILL  FILL_4__1669_
timestamp 1701859473
transform -1 0 6810 0 -1 790
box -12 -8 32 272
use FILL  FILL_4__1670_
timestamp 1701859473
transform 1 0 6590 0 -1 2870
box -12 -8 32 272
use FILL  FILL_4__1671_
timestamp 1701859473
transform -1 0 6390 0 -1 8590
box -12 -8 32 272
use FILL  FILL_4__1672_
timestamp 1701859473
transform 1 0 5950 0 -1 10670
box -12 -8 32 272
use FILL  FILL_4__1673_
timestamp 1701859473
transform 1 0 6350 0 1 8590
box -12 -8 32 272
use FILL  FILL_4__1674_
timestamp 1701859473
transform -1 0 6430 0 -1 9110
box -12 -8 32 272
use FILL  FILL_4__1675_
timestamp 1701859473
transform 1 0 90 0 -1 5470
box -12 -8 32 272
use FILL  FILL_4__1676_
timestamp 1701859473
transform -1 0 330 0 -1 5470
box -12 -8 32 272
use FILL  FILL_4__1677_
timestamp 1701859473
transform -1 0 570 0 1 5470
box -12 -8 32 272
use FILL  FILL_4__1678_
timestamp 1701859473
transform 1 0 90 0 -1 10670
box -12 -8 32 272
use FILL  FILL_4__1679_
timestamp 1701859473
transform -1 0 310 0 -1 11190
box -12 -8 32 272
use FILL  FILL_4__1680_
timestamp 1701859473
transform 1 0 290 0 -1 10670
box -12 -8 32 272
use FILL  FILL_4__1681_
timestamp 1701859473
transform -1 0 110 0 -1 7030
box -12 -8 32 272
use FILL  FILL_4__1682_
timestamp 1701859473
transform -1 0 110 0 1 7030
box -12 -8 32 272
use FILL  FILL_4__1683_
timestamp 1701859473
transform 1 0 90 0 1 6510
box -12 -8 32 272
use FILL  FILL_4__1684_
timestamp 1701859473
transform 1 0 970 0 -1 11190
box -12 -8 32 272
use FILL  FILL_4__1685_
timestamp 1701859473
transform -1 0 1230 0 -1 11190
box -12 -8 32 272
use FILL  FILL_4__1686_
timestamp 1701859473
transform -1 0 1030 0 1 10670
box -12 -8 32 272
use FILL  FILL_4__1687_
timestamp 1701859473
transform 1 0 1450 0 -1 11190
box -12 -8 32 272
use FILL  FILL_4__1688_
timestamp 1701859473
transform -1 0 1710 0 -1 11190
box -12 -8 32 272
use FILL  FILL_4__1689_
timestamp 1701859473
transform -1 0 1970 0 1 10150
box -12 -8 32 272
use FILL  FILL_4__1690_
timestamp 1701859473
transform 1 0 2130 0 1 9110
box -12 -8 32 272
use FILL  FILL_4__1691_
timestamp 1701859473
transform -1 0 2150 0 -1 9110
box -12 -8 32 272
use FILL  FILL_4__1692_
timestamp 1701859473
transform 1 0 90 0 1 790
box -12 -8 32 272
use FILL  FILL_4__1693_
timestamp 1701859473
transform 1 0 90 0 -1 1310
box -12 -8 32 272
use FILL  FILL_4__1694_
timestamp 1701859473
transform 1 0 510 0 -1 270
box -12 -8 32 272
use FILL  FILL_4__1695_
timestamp 1701859473
transform -1 0 730 0 -1 270
box -12 -8 32 272
use FILL  FILL_4__1696_
timestamp 1701859473
transform 1 0 1150 0 1 2870
box -12 -8 32 272
use FILL  FILL_4__1697_
timestamp 1701859473
transform -1 0 2810 0 -1 2870
box -12 -8 32 272
use FILL  FILL_4__1698_
timestamp 1701859473
transform -1 0 1910 0 1 3390
box -12 -8 32 272
use FILL  FILL_4__1699_
timestamp 1701859473
transform 1 0 3830 0 1 3390
box -12 -8 32 272
use FILL  FILL_4__1700_
timestamp 1701859473
transform -1 0 2630 0 -1 3910
box -12 -8 32 272
use FILL  FILL_4__1701_
timestamp 1701859473
transform -1 0 1170 0 1 270
box -12 -8 32 272
use FILL  FILL_4__1702_
timestamp 1701859473
transform 1 0 930 0 1 270
box -12 -8 32 272
use FILL  FILL_4__1703_
timestamp 1701859473
transform -1 0 1410 0 1 1830
box -12 -8 32 272
use FILL  FILL_4__1704_
timestamp 1701859473
transform -1 0 9170 0 1 2870
box -12 -8 32 272
use FILL  FILL_4__1705_
timestamp 1701859473
transform 1 0 9790 0 -1 790
box -12 -8 32 272
use FILL  FILL_4__1706_
timestamp 1701859473
transform -1 0 8010 0 -1 4950
box -12 -8 32 272
use FILL  FILL_4__1707_
timestamp 1701859473
transform 1 0 8450 0 -1 4950
box -12 -8 32 272
use FILL  FILL_4__1708_
timestamp 1701859473
transform 1 0 5070 0 -1 5990
box -12 -8 32 272
use FILL  FILL_4__1709_
timestamp 1701859473
transform -1 0 11170 0 1 5990
box -12 -8 32 272
use FILL  FILL_4__1710_
timestamp 1701859473
transform 1 0 5450 0 -1 5470
box -12 -8 32 272
use FILL  FILL_4__1711_
timestamp 1701859473
transform -1 0 5290 0 -1 5990
box -12 -8 32 272
use FILL  FILL_4__1712_
timestamp 1701859473
transform -1 0 5110 0 1 5470
box -12 -8 32 272
use FILL  FILL_4__1713_
timestamp 1701859473
transform 1 0 7970 0 1 4430
box -12 -8 32 272
use FILL  FILL_4__1714_
timestamp 1701859473
transform 1 0 7770 0 1 4950
box -12 -8 32 272
use FILL  FILL_4__1715_
timestamp 1701859473
transform -1 0 8010 0 1 4950
box -12 -8 32 272
use FILL  FILL_4__1716_
timestamp 1701859473
transform -1 0 8230 0 1 4430
box -12 -8 32 272
use FILL  FILL_4__1717_
timestamp 1701859473
transform -1 0 8010 0 1 1310
box -12 -8 32 272
use FILL  FILL_4__1718_
timestamp 1701859473
transform -1 0 5950 0 1 5990
box -12 -8 32 272
use FILL  FILL_4__1719_
timestamp 1701859473
transform -1 0 6810 0 -1 5990
box -12 -8 32 272
use FILL  FILL_4__1720_
timestamp 1701859473
transform -1 0 6790 0 1 5470
box -12 -8 32 272
use FILL  FILL_4__1721_
timestamp 1701859473
transform -1 0 7030 0 1 5470
box -12 -8 32 272
use FILL  FILL_4__1722_
timestamp 1701859473
transform -1 0 7730 0 1 4430
box -12 -8 32 272
use FILL  FILL_4__1723_
timestamp 1701859473
transform 1 0 7950 0 1 1830
box -12 -8 32 272
use FILL  FILL_4__1724_
timestamp 1701859473
transform -1 0 7990 0 -1 1310
box -12 -8 32 272
use FILL  FILL_4__1725_
timestamp 1701859473
transform 1 0 6590 0 1 5990
box -12 -8 32 272
use FILL  FILL_4__1726_
timestamp 1701859473
transform 1 0 6790 0 1 5990
box -12 -8 32 272
use FILL  FILL_4__1727_
timestamp 1701859473
transform -1 0 7030 0 1 5990
box -12 -8 32 272
use FILL  FILL_4__1728_
timestamp 1701859473
transform 1 0 7730 0 1 5990
box -12 -8 32 272
use FILL  FILL_4__1729_
timestamp 1701859473
transform -1 0 7670 0 -1 5990
box -12 -8 32 272
use FILL  FILL_4__1730_
timestamp 1701859473
transform -1 0 8150 0 1 3390
box -12 -8 32 272
use FILL  FILL_4__1731_
timestamp 1701859473
transform -1 0 8010 0 -1 270
box -12 -8 32 272
use FILL  FILL_4__1732_
timestamp 1701859473
transform -1 0 7970 0 1 5470
box -12 -8 32 272
use FILL  FILL_4__1733_
timestamp 1701859473
transform -1 0 8190 0 1 5470
box -12 -8 32 272
use FILL  FILL_4__1734_
timestamp 1701859473
transform 1 0 8150 0 -1 5470
box -12 -8 32 272
use FILL  FILL_4__1735_
timestamp 1701859473
transform 1 0 8610 0 -1 5470
box -12 -8 32 272
use FILL  FILL_4__1736_
timestamp 1701859473
transform 1 0 8450 0 1 4950
box -12 -8 32 272
use FILL  FILL_4__1737_
timestamp 1701859473
transform -1 0 8530 0 -1 3910
box -12 -8 32 272
use FILL  FILL_4__1738_
timestamp 1701859473
transform 1 0 8930 0 1 790
box -12 -8 32 272
use FILL  FILL_4__1739_
timestamp 1701859473
transform -1 0 9150 0 -1 790
box -12 -8 32 272
use FILL  FILL_4__1740_
timestamp 1701859473
transform 1 0 6510 0 1 270
box -12 -8 32 272
use FILL  FILL_4__1741_
timestamp 1701859473
transform 1 0 6410 0 1 790
box -12 -8 32 272
use FILL  FILL_4__1742_
timestamp 1701859473
transform -1 0 6350 0 -1 790
box -12 -8 32 272
use FILL  FILL_4__1743_
timestamp 1701859473
transform -1 0 2350 0 -1 3390
box -12 -8 32 272
use FILL  FILL_4__1744_
timestamp 1701859473
transform 1 0 330 0 -1 4950
box -12 -8 32 272
use FILL  FILL_4__1745_
timestamp 1701859473
transform 1 0 2150 0 -1 3910
box -12 -8 32 272
use FILL  FILL_4__1746_
timestamp 1701859473
transform -1 0 5170 0 -1 3390
box -12 -8 32 272
use FILL  FILL_4__1747_
timestamp 1701859473
transform -1 0 330 0 -1 270
box -12 -8 32 272
use FILL  FILL_4__1748_
timestamp 1701859473
transform -1 0 530 0 1 270
box -12 -8 32 272
use FILL  FILL_4__1749_
timestamp 1701859473
transform -1 0 970 0 1 1310
box -12 -8 32 272
use FILL  FILL_4__1750_
timestamp 1701859473
transform -1 0 1190 0 1 1310
box -12 -8 32 272
use FILL  FILL_4__1751_
timestamp 1701859473
transform -1 0 4550 0 -1 2870
box -12 -8 32 272
use FILL  FILL_4__1752_
timestamp 1701859473
transform 1 0 4750 0 -1 2870
box -12 -8 32 272
use FILL  FILL_4__1753_
timestamp 1701859473
transform -1 0 4370 0 1 790
box -12 -8 32 272
use FILL  FILL_4__1754_
timestamp 1701859473
transform 1 0 310 0 -1 790
box -12 -8 32 272
use FILL  FILL_4__1755_
timestamp 1701859473
transform -1 0 530 0 -1 790
box -12 -8 32 272
use FILL  FILL_4__1756_
timestamp 1701859473
transform -1 0 110 0 -1 270
box -12 -8 32 272
use FILL  FILL_4__1757_
timestamp 1701859473
transform 1 0 710 0 -1 790
box -12 -8 32 272
use FILL  FILL_4__1758_
timestamp 1701859473
transform 1 0 90 0 1 2350
box -12 -8 32 272
use FILL  FILL_4__1759_
timestamp 1701859473
transform -1 0 2590 0 -1 2870
box -12 -8 32 272
use FILL  FILL_4__1760_
timestamp 1701859473
transform 1 0 2970 0 -1 2870
box -12 -8 32 272
use FILL  FILL_4__1761_
timestamp 1701859473
transform -1 0 3290 0 -1 3390
box -12 -8 32 272
use FILL  FILL_4__1762_
timestamp 1701859473
transform -1 0 110 0 1 270
box -12 -8 32 272
use FILL  FILL_4__1763_
timestamp 1701859473
transform 1 0 90 0 -1 790
box -12 -8 32 272
use FILL  FILL_4__1764_
timestamp 1701859473
transform 1 0 530 0 1 1310
box -12 -8 32 272
use FILL  FILL_4__1765_
timestamp 1701859473
transform 1 0 1390 0 1 1310
box -12 -8 32 272
use FILL  FILL_4__1766_
timestamp 1701859473
transform -1 0 3190 0 -1 1830
box -12 -8 32 272
use FILL  FILL_4__1767_
timestamp 1701859473
transform 1 0 1490 0 -1 4430
box -12 -8 32 272
use FILL  FILL_4__1768_
timestamp 1701859473
transform 1 0 310 0 -1 1310
box -12 -8 32 272
use FILL  FILL_4__1769_
timestamp 1701859473
transform -1 0 530 0 1 1830
box -12 -8 32 272
use FILL  FILL_4__1770_
timestamp 1701859473
transform 1 0 2130 0 -1 3390
box -12 -8 32 272
use FILL  FILL_4__1771_
timestamp 1701859473
transform -1 0 2390 0 -1 3910
box -12 -8 32 272
use FILL  FILL_4__1772_
timestamp 1701859473
transform -1 0 3050 0 -1 3910
box -12 -8 32 272
use FILL  FILL_4__1773_
timestamp 1701859473
transform 1 0 3950 0 1 2870
box -12 -8 32 272
use FILL  FILL_4__1774_
timestamp 1701859473
transform -1 0 5330 0 -1 2350
box -12 -8 32 272
use FILL  FILL_4__1775_
timestamp 1701859473
transform 1 0 290 0 1 790
box -12 -8 32 272
use FILL  FILL_4__1776_
timestamp 1701859473
transform -1 0 330 0 1 1310
box -12 -8 32 272
use FILL  FILL_4__1777_
timestamp 1701859473
transform 1 0 750 0 -1 1830
box -12 -8 32 272
use FILL  FILL_4__1778_
timestamp 1701859473
transform -1 0 4470 0 1 5470
box -12 -8 32 272
use FILL  FILL_4__1779_
timestamp 1701859473
transform -1 0 6110 0 -1 5470
box -12 -8 32 272
use FILL  FILL_4__1780_
timestamp 1701859473
transform 1 0 4830 0 1 2870
box -12 -8 32 272
use FILL  FILL_4__1781_
timestamp 1701859473
transform 1 0 4410 0 1 2870
box -12 -8 32 272
use FILL  FILL_4__1782_
timestamp 1701859473
transform -1 0 110 0 1 1310
box -12 -8 32 272
use FILL  FILL_4__1783_
timestamp 1701859473
transform -1 0 1390 0 1 2870
box -12 -8 32 272
use FILL  FILL_4__1784_
timestamp 1701859473
transform -1 0 5090 0 1 2870
box -12 -8 32 272
use FILL  FILL_4__1785_
timestamp 1701859473
transform 1 0 5010 0 -1 2870
box -12 -8 32 272
use FILL  FILL_4__1786_
timestamp 1701859473
transform -1 0 5090 0 -1 2350
box -12 -8 32 272
use FILL  FILL_4__1787_
timestamp 1701859473
transform 1 0 5070 0 1 2350
box -12 -8 32 272
use FILL  FILL_4__1788_
timestamp 1701859473
transform -1 0 4870 0 -1 2350
box -12 -8 32 272
use FILL  FILL_4__1789_
timestamp 1701859473
transform 1 0 90 0 1 1830
box -12 -8 32 272
use FILL  FILL_4__1790_
timestamp 1701859473
transform -1 0 330 0 -1 2350
box -12 -8 32 272
use FILL  FILL_4__1791_
timestamp 1701859473
transform -1 0 2130 0 -1 2350
box -12 -8 32 272
use FILL  FILL_4__1792_
timestamp 1701859473
transform -1 0 3510 0 -1 2350
box -12 -8 32 272
use FILL  FILL_4__1793_
timestamp 1701859473
transform -1 0 4610 0 1 1830
box -12 -8 32 272
use FILL  FILL_4__1794_
timestamp 1701859473
transform 1 0 930 0 1 1830
box -12 -8 32 272
use FILL  FILL_4__1795_
timestamp 1701859473
transform -1 0 2190 0 1 2350
box -12 -8 32 272
use FILL  FILL_4__1796_
timestamp 1701859473
transform -1 0 1810 0 -1 1830
box -12 -8 32 272
use FILL  FILL_4__1797_
timestamp 1701859473
transform 1 0 2030 0 -1 1830
box -12 -8 32 272
use FILL  FILL_4__1798_
timestamp 1701859473
transform 1 0 950 0 -1 1310
box -12 -8 32 272
use FILL  FILL_4__1799_
timestamp 1701859473
transform 1 0 3770 0 1 3910
box -12 -8 32 272
use FILL  FILL_4__1800_
timestamp 1701859473
transform 1 0 3450 0 1 1830
box -12 -8 32 272
use FILL  FILL_4__1801_
timestamp 1701859473
transform -1 0 1190 0 1 1830
box -12 -8 32 272
use FILL  FILL_4__1802_
timestamp 1701859473
transform -1 0 3730 0 1 2350
box -12 -8 32 272
use FILL  FILL_4__1803_
timestamp 1701859473
transform -1 0 3950 0 1 2350
box -12 -8 32 272
use FILL  FILL_4__1804_
timestamp 1701859473
transform -1 0 4190 0 1 2350
box -12 -8 32 272
use FILL  FILL_4__1805_
timestamp 1701859473
transform 1 0 5490 0 1 2350
box -12 -8 32 272
use FILL  FILL_4__1806_
timestamp 1701859473
transform -1 0 4890 0 1 2350
box -12 -8 32 272
use FILL  FILL_4__1807_
timestamp 1701859473
transform -1 0 5290 0 1 2350
box -12 -8 32 272
use FILL  FILL_4__1808_
timestamp 1701859473
transform 1 0 4810 0 1 1830
box -12 -8 32 272
use FILL  FILL_4__1809_
timestamp 1701859473
transform -1 0 7170 0 -1 270
box -12 -8 32 272
use FILL  FILL_4__1810_
timestamp 1701859473
transform -1 0 7150 0 1 1310
box -12 -8 32 272
use FILL  FILL_4__1811_
timestamp 1701859473
transform 1 0 7490 0 -1 1830
box -12 -8 32 272
use FILL  FILL_4__1812_
timestamp 1701859473
transform -1 0 7570 0 -1 1310
box -12 -8 32 272
use FILL  FILL_4__1813_
timestamp 1701859473
transform 1 0 9150 0 1 790
box -12 -8 32 272
use FILL  FILL_4__1814_
timestamp 1701859473
transform -1 0 8190 0 -1 1830
box -12 -8 32 272
use FILL  FILL_4__1815_
timestamp 1701859473
transform 1 0 8390 0 1 2350
box -12 -8 32 272
use FILL  FILL_4__1816_
timestamp 1701859473
transform -1 0 9670 0 -1 2350
box -12 -8 32 272
use FILL  FILL_4__1817_
timestamp 1701859473
transform -1 0 9390 0 1 1310
box -12 -8 32 272
use FILL  FILL_4__1818_
timestamp 1701859473
transform -1 0 9590 0 1 270
box -12 -8 32 272
use FILL  FILL_4__1819_
timestamp 1701859473
transform -1 0 8410 0 -1 1830
box -12 -8 32 272
use FILL  FILL_4__1820_
timestamp 1701859473
transform -1 0 8490 0 1 1310
box -12 -8 32 272
use FILL  FILL_4__1821_
timestamp 1701859473
transform -1 0 4930 0 1 1310
box -12 -8 32 272
use FILL  FILL_4__1822_
timestamp 1701859473
transform -1 0 4730 0 -1 790
box -12 -8 32 272
use FILL  FILL_4__1823_
timestamp 1701859473
transform -1 0 4270 0 -1 790
box -12 -8 32 272
use FILL  FILL_4__1824_
timestamp 1701859473
transform 1 0 4650 0 1 2350
box -12 -8 32 272
use FILL  FILL_4__1825_
timestamp 1701859473
transform 1 0 5710 0 1 1830
box -12 -8 32 272
use FILL  FILL_4__1826_
timestamp 1701859473
transform 1 0 8210 0 -1 270
box -12 -8 32 272
use FILL  FILL_4__1827_
timestamp 1701859473
transform 1 0 9350 0 -1 790
box -12 -8 32 272
use FILL  FILL_4__1828_
timestamp 1701859473
transform 1 0 8510 0 1 270
box -12 -8 32 272
use FILL  FILL_4__1829_
timestamp 1701859473
transform 1 0 5810 0 1 270
box -12 -8 32 272
use FILL  FILL_4__1830_
timestamp 1701859473
transform 1 0 3250 0 1 4430
box -12 -8 32 272
use FILL  FILL_4__1831_
timestamp 1701859473
transform -1 0 8030 0 -1 790
box -12 -8 32 272
use FILL  FILL_4__1832_
timestamp 1701859473
transform 1 0 6530 0 -1 790
box -12 -8 32 272
use FILL  FILL_4__1833_
timestamp 1701859473
transform -1 0 730 0 1 270
box -12 -8 32 272
use FILL  FILL_4__1834_
timestamp 1701859473
transform 1 0 1170 0 -1 1310
box -12 -8 32 272
use FILL  FILL_4__1835_
timestamp 1701859473
transform -1 0 2550 0 -1 1310
box -12 -8 32 272
use FILL  FILL_4__1836_
timestamp 1701859473
transform 1 0 1110 0 1 790
box -12 -8 32 272
use FILL  FILL_4__1837_
timestamp 1701859473
transform -1 0 2510 0 1 790
box -12 -8 32 272
use FILL  FILL_4__1838_
timestamp 1701859473
transform 1 0 2250 0 1 790
box -12 -8 32 272
use FILL  FILL_4__1839_
timestamp 1701859473
transform -1 0 310 0 1 270
box -12 -8 32 272
use FILL  FILL_4__1840_
timestamp 1701859473
transform -1 0 950 0 1 2870
box -12 -8 32 272
use FILL  FILL_4__1841_
timestamp 1701859473
transform 1 0 3730 0 1 2870
box -12 -8 32 272
use FILL  FILL_4__1842_
timestamp 1701859473
transform -1 0 2990 0 -1 1830
box -12 -8 32 272
use FILL  FILL_4__1843_
timestamp 1701859473
transform -1 0 3950 0 -1 2350
box -12 -8 32 272
use FILL  FILL_4__1844_
timestamp 1701859473
transform 1 0 3850 0 -1 2870
box -12 -8 32 272
use FILL  FILL_4__1845_
timestamp 1701859473
transform -1 0 1790 0 -1 4950
box -12 -8 32 272
use FILL  FILL_4__1846_
timestamp 1701859473
transform 1 0 4150 0 1 4430
box -12 -8 32 272
use FILL  FILL_4__1847_
timestamp 1701859473
transform 1 0 3470 0 1 4430
box -12 -8 32 272
use FILL  FILL_4__1848_
timestamp 1701859473
transform 1 0 3910 0 1 4430
box -12 -8 32 272
use FILL  FILL_4__1849_
timestamp 1701859473
transform -1 0 4110 0 -1 2870
box -12 -8 32 272
use FILL  FILL_4__1850_
timestamp 1701859473
transform -1 0 930 0 1 790
box -12 -8 32 272
use FILL  FILL_4__1851_
timestamp 1701859473
transform 1 0 1590 0 -1 1830
box -12 -8 32 272
use FILL  FILL_4__1852_
timestamp 1701859473
transform -1 0 2410 0 1 2350
box -12 -8 32 272
use FILL  FILL_4__1853_
timestamp 1701859473
transform 1 0 90 0 -1 2350
box -12 -8 32 272
use FILL  FILL_4__1854_
timestamp 1701859473
transform 1 0 2330 0 -1 2350
box -12 -8 32 272
use FILL  FILL_4__1855_
timestamp 1701859473
transform -1 0 2590 0 -1 2350
box -12 -8 32 272
use FILL  FILL_4__1856_
timestamp 1701859473
transform 1 0 1490 0 -1 790
box -12 -8 32 272
use FILL  FILL_4__1857_
timestamp 1701859473
transform -1 0 2690 0 -1 790
box -12 -8 32 272
use FILL  FILL_4__1858_
timestamp 1701859473
transform 1 0 2430 0 -1 790
box -12 -8 32 272
use FILL  FILL_4__1859_
timestamp 1701859473
transform 1 0 2210 0 -1 790
box -12 -8 32 272
use FILL  FILL_4__1860_
timestamp 1701859473
transform -1 0 1750 0 -1 790
box -12 -8 32 272
use FILL  FILL_4__1861_
timestamp 1701859473
transform -1 0 1990 0 -1 790
box -12 -8 32 272
use FILL  FILL_4__1862_
timestamp 1701859473
transform -1 0 2070 0 1 270
box -12 -8 32 272
use FILL  FILL_4__1863_
timestamp 1701859473
transform 1 0 2290 0 1 270
box -12 -8 32 272
use FILL  FILL_4__1864_
timestamp 1701859473
transform 1 0 3530 0 1 270
box -12 -8 32 272
use FILL  FILL_4__1865_
timestamp 1701859473
transform 1 0 7330 0 -1 1310
box -12 -8 32 272
use FILL  FILL_4__1866_
timestamp 1701859473
transform 1 0 3690 0 -1 1310
box -12 -8 32 272
use FILL  FILL_4__1867_
timestamp 1701859473
transform 1 0 1150 0 -1 1830
box -12 -8 32 272
use FILL  FILL_4__1868_
timestamp 1701859473
transform 1 0 1590 0 1 1310
box -12 -8 32 272
use FILL  FILL_4__1869_
timestamp 1701859473
transform 1 0 2010 0 1 1310
box -12 -8 32 272
use FILL  FILL_4__1870_
timestamp 1701859473
transform -1 0 1630 0 -1 1310
box -12 -8 32 272
use FILL  FILL_4__1871_
timestamp 1701859473
transform -1 0 2750 0 -1 1310
box -12 -8 32 272
use FILL  FILL_4__1872_
timestamp 1701859473
transform -1 0 530 0 1 790
box -12 -8 32 272
use FILL  FILL_4__1873_
timestamp 1701859473
transform 1 0 710 0 1 790
box -12 -8 32 272
use FILL  FILL_4__1874_
timestamp 1701859473
transform -1 0 1350 0 1 790
box -12 -8 32 272
use FILL  FILL_4__1875_
timestamp 1701859473
transform 1 0 930 0 -1 790
box -12 -8 32 272
use FILL  FILL_4__1876_
timestamp 1701859473
transform 1 0 1250 0 -1 790
box -12 -8 32 272
use FILL  FILL_4__1877_
timestamp 1701859473
transform 1 0 2190 0 1 4950
box -12 -8 32 272
use FILL  FILL_4__1878_
timestamp 1701859473
transform 1 0 530 0 -1 1310
box -12 -8 32 272
use FILL  FILL_4__1879_
timestamp 1701859473
transform 1 0 750 0 1 1310
box -12 -8 32 272
use FILL  FILL_4__1880_
timestamp 1701859473
transform -1 0 2010 0 -1 4950
box -12 -8 32 272
use FILL  FILL_4__1881_
timestamp 1701859473
transform -1 0 2250 0 -1 4950
box -12 -8 32 272
use FILL  FILL_4__1882_
timestamp 1701859473
transform 1 0 1570 0 -1 3390
box -12 -8 32 272
use FILL  FILL_4__1883_
timestamp 1701859473
transform 1 0 1050 0 -1 3390
box -12 -8 32 272
use FILL  FILL_4__1884_
timestamp 1701859473
transform -1 0 4070 0 1 3390
box -12 -8 32 272
use FILL  FILL_4__1885_
timestamp 1701859473
transform -1 0 3790 0 -1 3390
box -12 -8 32 272
use FILL  FILL_4__1886_
timestamp 1701859473
transform 1 0 3530 0 -1 3390
box -12 -8 32 272
use FILL  FILL_4__1887_
timestamp 1701859473
transform -1 0 3510 0 1 2870
box -12 -8 32 272
use FILL  FILL_4__1888_
timestamp 1701859473
transform -1 0 2550 0 1 270
box -12 -8 32 272
use FILL  FILL_4__1889_
timestamp 1701859473
transform 1 0 1690 0 -1 2870
box -12 -8 32 272
use FILL  FILL_4__1890_
timestamp 1701859473
transform -1 0 330 0 -1 1830
box -12 -8 32 272
use FILL  FILL_4__1891_
timestamp 1701859473
transform 1 0 90 0 -1 1830
box -12 -8 32 272
use FILL  FILL_4__1892_
timestamp 1701859473
transform 1 0 4930 0 -1 3390
box -12 -8 32 272
use FILL  FILL_4__1893_
timestamp 1701859473
transform 1 0 3930 0 1 1830
box -12 -8 32 272
use FILL  FILL_4__1894_
timestamp 1701859473
transform 1 0 4130 0 1 1830
box -12 -8 32 272
use FILL  FILL_4__1895_
timestamp 1701859473
transform -1 0 1870 0 1 1830
box -12 -8 32 272
use FILL  FILL_4__1896_
timestamp 1701859473
transform 1 0 1890 0 -1 2350
box -12 -8 32 272
use FILL  FILL_4__1897_
timestamp 1701859473
transform 1 0 3510 0 1 2350
box -12 -8 32 272
use FILL  FILL_4__1898_
timestamp 1701859473
transform 1 0 3290 0 1 2350
box -12 -8 32 272
use FILL  FILL_4__1899_
timestamp 1701859473
transform -1 0 3270 0 -1 2350
box -12 -8 32 272
use FILL  FILL_4__1900_
timestamp 1701859473
transform -1 0 4110 0 -1 1830
box -12 -8 32 272
use FILL  FILL_4__1901_
timestamp 1701859473
transform -1 0 750 0 1 1830
box -12 -8 32 272
use FILL  FILL_4__1902_
timestamp 1701859473
transform 1 0 5050 0 1 1830
box -12 -8 32 272
use FILL  FILL_4__1903_
timestamp 1701859473
transform 1 0 3370 0 1 1310
box -12 -8 32 272
use FILL  FILL_4__1904_
timestamp 1701859473
transform -1 0 3470 0 -1 1310
box -12 -8 32 272
use FILL  FILL_4__1905_
timestamp 1701859473
transform 1 0 3010 0 1 270
box -12 -8 32 272
use FILL  FILL_4__1906_
timestamp 1701859473
transform 1 0 290 0 1 2350
box -12 -8 32 272
use FILL  FILL_4__1907_
timestamp 1701859473
transform -1 0 3050 0 -1 2350
box -12 -8 32 272
use FILL  FILL_4__1908_
timestamp 1701859473
transform 1 0 6470 0 -1 2350
box -12 -8 32 272
use FILL  FILL_4__1909_
timestamp 1701859473
transform -1 0 6070 0 -1 2350
box -12 -8 32 272
use FILL  FILL_4__1910_
timestamp 1701859473
transform -1 0 5570 0 -1 2350
box -12 -8 32 272
use FILL  FILL_4__1911_
timestamp 1701859473
transform -1 0 730 0 1 2870
box -12 -8 32 272
use FILL  FILL_4__1912_
timestamp 1701859473
transform -1 0 3330 0 1 3910
box -12 -8 32 272
use FILL  FILL_4__1913_
timestamp 1701859473
transform -1 0 1050 0 -1 2870
box -12 -8 32 272
use FILL  FILL_4__1914_
timestamp 1701859473
transform -1 0 1490 0 1 3390
box -12 -8 32 272
use FILL  FILL_4__1915_
timestamp 1701859473
transform 1 0 2570 0 1 3390
box -12 -8 32 272
use FILL  FILL_4__1916_
timestamp 1701859473
transform -1 0 3430 0 1 3390
box -12 -8 32 272
use FILL  FILL_4__1917_
timestamp 1701859473
transform -1 0 4710 0 -1 3390
box -12 -8 32 272
use FILL  FILL_4__1918_
timestamp 1701859473
transform 1 0 1750 0 1 4950
box -12 -8 32 272
use FILL  FILL_4__1919_
timestamp 1701859473
transform -1 0 1270 0 -1 2870
box -12 -8 32 272
use FILL  FILL_4__1920_
timestamp 1701859473
transform -1 0 5050 0 1 4430
box -12 -8 32 272
use FILL  FILL_4__1921_
timestamp 1701859473
transform 1 0 4810 0 1 4430
box -12 -8 32 272
use FILL  FILL_4__1922_
timestamp 1701859473
transform -1 0 4610 0 1 4430
box -12 -8 32 272
use FILL  FILL_4__1923_
timestamp 1701859473
transform 1 0 4470 0 -1 3390
box -12 -8 32 272
use FILL  FILL_4__1924_
timestamp 1701859473
transform 1 0 1970 0 1 4950
box -12 -8 32 272
use FILL  FILL_4__1925_
timestamp 1701859473
transform 1 0 6110 0 -1 4430
box -12 -8 32 272
use FILL  FILL_4__1926_
timestamp 1701859473
transform 1 0 730 0 -1 1310
box -12 -8 32 272
use FILL  FILL_4__1927_
timestamp 1701859473
transform 1 0 2970 0 -1 1310
box -12 -8 32 272
use FILL  FILL_4__1928_
timestamp 1701859473
transform -1 0 3230 0 -1 1310
box -12 -8 32 272
use FILL  FILL_4__1929_
timestamp 1701859473
transform 1 0 3410 0 1 790
box -12 -8 32 272
use FILL  FILL_4__1930_
timestamp 1701859473
transform 1 0 3230 0 1 270
box -12 -8 32 272
use FILL  FILL_4__1931_
timestamp 1701859473
transform 1 0 3830 0 1 270
box -12 -8 32 272
use FILL  FILL_4__1932_
timestamp 1701859473
transform -1 0 4070 0 1 270
box -12 -8 32 272
use FILL  FILL_4__1933_
timestamp 1701859473
transform -1 0 1870 0 1 270
box -12 -8 32 272
use FILL  FILL_4__1934_
timestamp 1701859473
transform -1 0 5490 0 1 790
box -12 -8 32 272
use FILL  FILL_4__1935_
timestamp 1701859473
transform 1 0 5610 0 -1 270
box -12 -8 32 272
use FILL  FILL_4__1936_
timestamp 1701859473
transform -1 0 8370 0 1 3390
box -12 -8 32 272
use FILL  FILL_4__1937_
timestamp 1701859473
transform -1 0 7590 0 -1 270
box -12 -8 32 272
use FILL  FILL_4__1938_
timestamp 1701859473
transform -1 0 7790 0 -1 270
box -12 -8 32 272
use FILL  FILL_4__1939_
timestamp 1701859473
transform -1 0 6710 0 -1 270
box -12 -8 32 272
use FILL  FILL_4__1940_
timestamp 1701859473
transform -1 0 5830 0 -1 270
box -12 -8 32 272
use FILL  FILL_4__1941_
timestamp 1701859473
transform 1 0 5850 0 -1 790
box -12 -8 32 272
use FILL  FILL_4__1942_
timestamp 1701859473
transform 1 0 4830 0 -1 1310
box -12 -8 32 272
use FILL  FILL_4__1943_
timestamp 1701859473
transform 1 0 8090 0 1 270
box -12 -8 32 272
use FILL  FILL_4__1944_
timestamp 1701859473
transform -1 0 8330 0 1 270
box -12 -8 32 272
use FILL  FILL_4__1945_
timestamp 1701859473
transform 1 0 7870 0 1 270
box -12 -8 32 272
use FILL  FILL_4__1946_
timestamp 1701859473
transform -1 0 6070 0 1 270
box -12 -8 32 272
use FILL  FILL_4__1947_
timestamp 1701859473
transform -1 0 6090 0 -1 790
box -12 -8 32 272
use FILL  FILL_4__1948_
timestamp 1701859473
transform 1 0 5370 0 -1 790
box -12 -8 32 272
use FILL  FILL_4__1949_
timestamp 1701859473
transform 1 0 4610 0 -1 1310
box -12 -8 32 272
use FILL  FILL_4__1950_
timestamp 1701859473
transform -1 0 8250 0 -1 790
box -12 -8 32 272
use FILL  FILL_4__1951_
timestamp 1701859473
transform 1 0 530 0 -1 2350
box -12 -8 32 272
use FILL  FILL_4__1952_
timestamp 1701859473
transform -1 0 5710 0 1 2350
box -12 -8 32 272
use FILL  FILL_4__1953_
timestamp 1701859473
transform 1 0 5810 0 -1 2350
box -12 -8 32 272
use FILL  FILL_4__1954_
timestamp 1701859473
transform 1 0 8190 0 -1 1310
box -12 -8 32 272
use FILL  FILL_4__1955_
timestamp 1701859473
transform -1 0 8730 0 1 1310
box -12 -8 32 272
use FILL  FILL_4__1956_
timestamp 1701859473
transform -1 0 6270 0 -1 1310
box -12 -8 32 272
use FILL  FILL_4__1957_
timestamp 1701859473
transform -1 0 6030 0 -1 1310
box -12 -8 32 272
use FILL  FILL_4__1958_
timestamp 1701859473
transform 1 0 5290 0 -1 1310
box -12 -8 32 272
use FILL  FILL_4__1959_
timestamp 1701859473
transform 1 0 5730 0 -1 2870
box -12 -8 32 272
use FILL  FILL_4__1960_
timestamp 1701859473
transform -1 0 6170 0 -1 2870
box -12 -8 32 272
use FILL  FILL_4__1961_
timestamp 1701859473
transform -1 0 4430 0 1 2350
box -12 -8 32 272
use FILL  FILL_4__1962_
timestamp 1701859473
transform 1 0 5890 0 1 2350
box -12 -8 32 272
use FILL  FILL_4__1963_
timestamp 1701859473
transform 1 0 5350 0 1 1310
box -12 -8 32 272
use FILL  FILL_4__1964_
timestamp 1701859473
transform 1 0 9170 0 1 1310
box -12 -8 32 272
use FILL  FILL_4__1965_
timestamp 1701859473
transform 1 0 7570 0 1 790
box -12 -8 32 272
use FILL  FILL_4__1966_
timestamp 1701859473
transform -1 0 7690 0 1 270
box -12 -8 32 272
use FILL  FILL_4__1967_
timestamp 1701859473
transform -1 0 6750 0 1 270
box -12 -8 32 272
use FILL  FILL_4__1968_
timestamp 1701859473
transform 1 0 5530 0 -1 1310
box -12 -8 32 272
use FILL  FILL_4__1969_
timestamp 1701859473
transform 1 0 5730 0 1 2870
box -12 -8 32 272
use FILL  FILL_4__1970_
timestamp 1701859473
transform 1 0 5370 0 -1 3390
box -12 -8 32 272
use FILL  FILL_4__1971_
timestamp 1701859473
transform 1 0 5810 0 1 3910
box -12 -8 32 272
use FILL  FILL_4__1972_
timestamp 1701859473
transform 1 0 5750 0 1 4950
box -12 -8 32 272
use FILL  FILL_4__1973_
timestamp 1701859473
transform -1 0 6090 0 -1 3910
box -12 -8 32 272
use FILL  FILL_4__1974_
timestamp 1701859473
transform 1 0 6270 0 -1 3910
box -12 -8 32 272
use FILL  FILL_4__1975_
timestamp 1701859473
transform -1 0 6070 0 1 3910
box -12 -8 32 272
use FILL  FILL_4__1976_
timestamp 1701859473
transform -1 0 6530 0 -1 3910
box -12 -8 32 272
use FILL  FILL_4__1977_
timestamp 1701859473
transform 1 0 6850 0 1 2870
box -12 -8 32 272
use FILL  FILL_4__1978_
timestamp 1701859473
transform -1 0 6390 0 -1 2870
box -12 -8 32 272
use FILL  FILL_4__1979_
timestamp 1701859473
transform 1 0 6430 0 1 2870
box -12 -8 32 272
use FILL  FILL_4__1980_
timestamp 1701859473
transform 1 0 6630 0 1 2870
box -12 -8 32 272
use FILL  FILL_4__1981_
timestamp 1701859473
transform 1 0 6210 0 1 2870
box -12 -8 32 272
use FILL  FILL_4__1982_
timestamp 1701859473
transform -1 0 5670 0 -1 1830
box -12 -8 32 272
use FILL  FILL_4__1983_
timestamp 1701859473
transform -1 0 4770 0 -1 270
box -12 -8 32 272
use FILL  FILL_4__1984_
timestamp 1701859473
transform -1 0 6470 0 -1 1310
box -12 -8 32 272
use FILL  FILL_4__1985_
timestamp 1701859473
transform 1 0 5030 0 -1 1310
box -12 -8 32 272
use FILL  FILL_4__1986_
timestamp 1701859473
transform 1 0 8230 0 1 790
box -12 -8 32 272
use FILL  FILL_4__1987_
timestamp 1701859473
transform 1 0 6910 0 1 1310
box -12 -8 32 272
use FILL  FILL_4__1988_
timestamp 1701859473
transform -1 0 7370 0 1 1310
box -12 -8 32 272
use FILL  FILL_4__1989_
timestamp 1701859473
transform 1 0 2730 0 -1 5470
box -12 -8 32 272
use FILL  FILL_4__1990_
timestamp 1701859473
transform 1 0 2050 0 1 1830
box -12 -8 32 272
use FILL  FILL_4__1991_
timestamp 1701859473
transform -1 0 2770 0 1 1830
box -12 -8 32 272
use FILL  FILL_4__1992_
timestamp 1701859473
transform -1 0 4170 0 -1 2350
box -12 -8 32 272
use FILL  FILL_4__1993_
timestamp 1701859473
transform -1 0 4410 0 -1 2350
box -12 -8 32 272
use FILL  FILL_4__1994_
timestamp 1701859473
transform 1 0 2510 0 1 1830
box -12 -8 32 272
use FILL  FILL_4__1995_
timestamp 1701859473
transform 1 0 2990 0 1 1830
box -12 -8 32 272
use FILL  FILL_4__1996_
timestamp 1701859473
transform -1 0 6670 0 1 790
box -12 -8 32 272
use FILL  FILL_4__1997_
timestamp 1701859473
transform -1 0 5010 0 1 790
box -12 -8 32 272
use FILL  FILL_4__1998_
timestamp 1701859473
transform 1 0 4270 0 1 270
box -12 -8 32 272
use FILL  FILL_4__1999_
timestamp 1701859473
transform -1 0 3870 0 -1 270
box -12 -8 32 272
use FILL  FILL_4__2000_
timestamp 1701859473
transform -1 0 4550 0 -1 270
box -12 -8 32 272
use FILL  FILL_4__2001_
timestamp 1701859473
transform -1 0 5930 0 -1 2870
box -12 -8 32 272
use FILL  FILL_4__2002_
timestamp 1701859473
transform -1 0 1870 0 1 2870
box -12 -8 32 272
use FILL  FILL_4__2003_
timestamp 1701859473
transform 1 0 1370 0 -1 3390
box -12 -8 32 272
use FILL  FILL_4__2004_
timestamp 1701859473
transform 1 0 2790 0 -1 3390
box -12 -8 32 272
use FILL  FILL_4__2005_
timestamp 1701859473
transform -1 0 3070 0 1 2870
box -12 -8 32 272
use FILL  FILL_4__2006_
timestamp 1701859473
transform 1 0 2810 0 1 2870
box -12 -8 32 272
use FILL  FILL_4__2007_
timestamp 1701859473
transform 1 0 6830 0 -1 2870
box -12 -8 32 272
use FILL  FILL_4__2008_
timestamp 1701859473
transform 1 0 510 0 -1 1830
box -12 -8 32 272
use FILL  FILL_4__2009_
timestamp 1701859473
transform -1 0 4030 0 -1 3390
box -12 -8 32 272
use FILL  FILL_4__2010_
timestamp 1701859473
transform -1 0 4330 0 -1 2870
box -12 -8 32 272
use FILL  FILL_4__2011_
timestamp 1701859473
transform -1 0 2070 0 1 790
box -12 -8 32 272
use FILL  FILL_4__2012_
timestamp 1701859473
transform 1 0 1570 0 1 790
box -12 -8 32 272
use FILL  FILL_4__2013_
timestamp 1701859473
transform -1 0 1830 0 1 790
box -12 -8 32 272
use FILL  FILL_4__2014_
timestamp 1701859473
transform 1 0 4490 0 1 1310
box -12 -8 32 272
use FILL  FILL_4__2015_
timestamp 1701859473
transform 1 0 3210 0 1 1830
box -12 -8 32 272
use FILL  FILL_4__2016_
timestamp 1701859473
transform -1 0 3710 0 1 1830
box -12 -8 32 272
use FILL  FILL_4__2017_
timestamp 1701859473
transform -1 0 5230 0 -1 1830
box -12 -8 32 272
use FILL  FILL_4__2018_
timestamp 1701859473
transform 1 0 4990 0 -1 1830
box -12 -8 32 272
use FILL  FILL_4__2019_
timestamp 1701859473
transform -1 0 5510 0 -1 2870
box -12 -8 32 272
use FILL  FILL_4__2020_
timestamp 1701859473
transform -1 0 5270 0 -1 2870
box -12 -8 32 272
use FILL  FILL_4__2021_
timestamp 1701859473
transform -1 0 6910 0 -1 1310
box -12 -8 32 272
use FILL  FILL_4__2022_
timestamp 1701859473
transform -1 0 7150 0 1 790
box -12 -8 32 272
use FILL  FILL_4__2023_
timestamp 1701859473
transform 1 0 8190 0 1 1830
box -12 -8 32 272
use FILL  FILL_4__2024_
timestamp 1701859473
transform -1 0 8410 0 1 1830
box -12 -8 32 272
use FILL  FILL_4__2025_
timestamp 1701859473
transform 1 0 9570 0 -1 790
box -12 -8 32 272
use FILL  FILL_4__2026_
timestamp 1701859473
transform -1 0 8710 0 1 790
box -12 -8 32 272
use FILL  FILL_4__2027_
timestamp 1701859473
transform -1 0 6910 0 1 790
box -12 -8 32 272
use FILL  FILL_4__2028_
timestamp 1701859473
transform 1 0 7010 0 -1 790
box -12 -8 32 272
use FILL  FILL_4__2029_
timestamp 1701859473
transform 1 0 7450 0 1 270
box -12 -8 32 272
use FILL  FILL_4__2030_
timestamp 1701859473
transform -1 0 7130 0 -1 1310
box -12 -8 32 272
use FILL  FILL_4__2031_
timestamp 1701859473
transform 1 0 7450 0 -1 790
box -12 -8 32 272
use FILL  FILL_4__2032_
timestamp 1701859473
transform -1 0 8750 0 1 270
box -12 -8 32 272
use FILL  FILL_4__2033_
timestamp 1701859473
transform 1 0 8230 0 1 1310
box -12 -8 32 272
use FILL  FILL_4__2034_
timestamp 1701859473
transform -1 0 8910 0 -1 1310
box -12 -8 32 272
use FILL  FILL_4__2035_
timestamp 1701859473
transform -1 0 8490 0 1 790
box -12 -8 32 272
use FILL  FILL_4__2036_
timestamp 1701859473
transform -1 0 8650 0 -1 1830
box -12 -8 32 272
use FILL  FILL_4__2037_
timestamp 1701859473
transform -1 0 8710 0 -1 790
box -12 -8 32 272
use FILL  FILL_4__2038_
timestamp 1701859473
transform 1 0 8010 0 1 790
box -12 -8 32 272
use FILL  FILL_4__2039_
timestamp 1701859473
transform 1 0 7790 0 1 790
box -12 -8 32 272
use FILL  FILL_4__2040_
timestamp 1701859473
transform -1 0 7710 0 -1 790
box -12 -8 32 272
use FILL  FILL_4__2041_
timestamp 1701859473
transform -1 0 6930 0 -1 270
box -12 -8 32 272
use FILL  FILL_4__2042_
timestamp 1701859473
transform 1 0 8910 0 -1 790
box -12 -8 32 272
use FILL  FILL_4__2043_
timestamp 1701859473
transform 1 0 7230 0 1 270
box -12 -8 32 272
use FILL  FILL_4__2044_
timestamp 1701859473
transform 1 0 6970 0 1 270
box -12 -8 32 272
use FILL  FILL_4__2045_
timestamp 1701859473
transform -1 0 6290 0 1 270
box -12 -8 32 272
use FILL  FILL_4__2046_
timestamp 1701859473
transform 1 0 6470 0 -1 270
box -12 -8 32 272
use FILL  FILL_4__2047_
timestamp 1701859473
transform -1 0 6250 0 -1 270
box -12 -8 32 272
use FILL  FILL_4__2048_
timestamp 1701859473
transform -1 0 6050 0 -1 270
box -12 -8 32 272
use FILL  FILL_4__2049_
timestamp 1701859473
transform -1 0 7230 0 -1 790
box -12 -8 32 272
use FILL  FILL_4__2050_
timestamp 1701859473
transform 1 0 1470 0 -1 2870
box -12 -8 32 272
use FILL  FILL_4__2051_
timestamp 1701859473
transform 1 0 6270 0 -1 2350
box -12 -8 32 272
use FILL  FILL_4__2052_
timestamp 1701859473
transform -1 0 6170 0 1 790
box -12 -8 32 272
use FILL  FILL_4__2053_
timestamp 1701859473
transform -1 0 4390 0 1 1830
box -12 -8 32 272
use FILL  FILL_4__2054_
timestamp 1701859473
transform 1 0 2890 0 1 1310
box -12 -8 32 272
use FILL  FILL_4__2055_
timestamp 1701859473
transform -1 0 3150 0 1 1310
box -12 -8 32 272
use FILL  FILL_4__2056_
timestamp 1701859473
transform -1 0 1870 0 -1 1310
box -12 -8 32 272
use FILL  FILL_4__2057_
timestamp 1701859473
transform 1 0 2730 0 1 790
box -12 -8 32 272
use FILL  FILL_4__2058_
timestamp 1701859473
transform 1 0 3650 0 1 790
box -12 -8 32 272
use FILL  FILL_4__2059_
timestamp 1701859473
transform 1 0 3890 0 1 790
box -12 -8 32 272
use FILL  FILL_4__2060_
timestamp 1701859473
transform -1 0 4130 0 1 790
box -12 -8 32 272
use FILL  FILL_4__2061_
timestamp 1701859473
transform -1 0 2990 0 -1 270
box -12 -8 32 272
use FILL  FILL_4__2062_
timestamp 1701859473
transform 1 0 2770 0 1 270
box -12 -8 32 272
use FILL  FILL_4__2063_
timestamp 1701859473
transform 1 0 3150 0 -1 270
box -12 -8 32 272
use FILL  FILL_4__2064_
timestamp 1701859473
transform 1 0 3390 0 -1 270
box -12 -8 32 272
use FILL  FILL_4__2065_
timestamp 1701859473
transform -1 0 3630 0 -1 270
box -12 -8 32 272
use FILL  FILL_4__2066_
timestamp 1701859473
transform -1 0 5410 0 -1 270
box -12 -8 32 272
use FILL  FILL_4__2067_
timestamp 1701859473
transform 1 0 7350 0 1 790
box -12 -8 32 272
use FILL  FILL_4__2068_
timestamp 1701859473
transform 1 0 5910 0 1 790
box -12 -8 32 272
use FILL  FILL_4__2069_
timestamp 1701859473
transform 1 0 3390 0 -1 1830
box -12 -8 32 272
use FILL  FILL_4__2070_
timestamp 1701859473
transform -1 0 3870 0 -1 1830
box -12 -8 32 272
use FILL  FILL_4__2071_
timestamp 1701859473
transform -1 0 5710 0 1 790
box -12 -8 32 272
use FILL  FILL_4__2072_
timestamp 1701859473
transform -1 0 7770 0 1 1310
box -12 -8 32 272
use FILL  FILL_4__2073_
timestamp 1701859473
transform 1 0 6650 0 1 1310
box -12 -8 32 272
use FILL  FILL_4__2074_
timestamp 1701859473
transform 1 0 1790 0 1 1310
box -12 -8 32 272
use FILL  FILL_4__2075_
timestamp 1701859473
transform -1 0 2270 0 1 1310
box -12 -8 32 272
use FILL  FILL_4__2076_
timestamp 1701859473
transform -1 0 2310 0 -1 1310
box -12 -8 32 272
use FILL  FILL_4__2077_
timestamp 1701859473
transform 1 0 4170 0 -1 1310
box -12 -8 32 272
use FILL  FILL_4__2078_
timestamp 1701859473
transform -1 0 2310 0 1 1830
box -12 -8 32 272
use FILL  FILL_4__2079_
timestamp 1701859473
transform -1 0 950 0 -1 1830
box -12 -8 32 272
use FILL  FILL_4__2080_
timestamp 1701859473
transform 1 0 2270 0 -1 1830
box -12 -8 32 272
use FILL  FILL_4__2081_
timestamp 1701859473
transform 1 0 2510 0 -1 1830
box -12 -8 32 272
use FILL  FILL_4__2082_
timestamp 1701859473
transform -1 0 2730 0 -1 1830
box -12 -8 32 272
use FILL  FILL_4__2083_
timestamp 1701859473
transform 1 0 4410 0 -1 1310
box -12 -8 32 272
use FILL  FILL_4__2084_
timestamp 1701859473
transform -1 0 5250 0 1 790
box -12 -8 32 272
use FILL  FILL_4__2085_
timestamp 1701859473
transform -1 0 5090 0 -1 270
box -12 -8 32 272
use FILL  FILL_4__2086_
timestamp 1701859473
transform -1 0 4310 0 -1 270
box -12 -8 32 272
use FILL  FILL_4__2087_
timestamp 1701859473
transform -1 0 4790 0 1 790
box -12 -8 32 272
use FILL  FILL_4__2088_
timestamp 1701859473
transform -1 0 5630 0 1 270
box -12 -8 32 272
use FILL  FILL_4__2089_
timestamp 1701859473
transform 1 0 5390 0 1 270
box -12 -8 32 272
use FILL  FILL_4__2090_
timestamp 1701859473
transform -1 0 4970 0 -1 790
box -12 -8 32 272
use FILL  FILL_4__2091_
timestamp 1701859473
transform 1 0 3190 0 1 790
box -12 -8 32 272
use FILL  FILL_4__2092_
timestamp 1701859473
transform 1 0 2750 0 -1 270
box -12 -8 32 272
use FILL  FILL_4__2093_
timestamp 1701859473
transform -1 0 2910 0 -1 790
box -12 -8 32 272
use FILL  FILL_4__2094_
timestamp 1701859473
transform 1 0 2310 0 -1 270
box -12 -8 32 272
use FILL  FILL_4__2095_
timestamp 1701859473
transform 1 0 2510 0 -1 270
box -12 -8 32 272
use FILL  FILL_4__2096_
timestamp 1701859473
transform -1 0 4970 0 1 270
box -12 -8 32 272
use FILL  FILL_4__2097_
timestamp 1701859473
transform -1 0 5190 0 1 270
box -12 -8 32 272
use FILL  FILL_4__2098_
timestamp 1701859473
transform 1 0 4730 0 1 270
box -12 -8 32 272
use FILL  FILL_4__2099_
timestamp 1701859473
transform 1 0 4050 0 -1 270
box -12 -8 32 272
use FILL  FILL_4__2100_
timestamp 1701859473
transform -1 0 5910 0 -1 1830
box -12 -8 32 272
use FILL  FILL_4__2101_
timestamp 1701859473
transform -1 0 5830 0 1 1310
box -12 -8 32 272
use FILL  FILL_4__2102_
timestamp 1701859473
transform -1 0 6230 0 1 1310
box -12 -8 32 272
use FILL  FILL_4__2103_
timestamp 1701859473
transform 1 0 5790 0 -1 1310
box -12 -8 32 272
use FILL  FILL_4__2104_
timestamp 1701859473
transform -1 0 6030 0 1 1310
box -12 -8 32 272
use FILL  FILL_4__2105_
timestamp 1701859473
transform -1 0 4330 0 -1 1830
box -12 -8 32 272
use FILL  FILL_4__2106_
timestamp 1701859473
transform 1 0 4010 0 -1 790
box -12 -8 32 272
use FILL  FILL_4__2107_
timestamp 1701859473
transform -1 0 3590 0 -1 790
box -12 -8 32 272
use FILL  FILL_4__2108_
timestamp 1701859473
transform 1 0 2950 0 1 790
box -12 -8 32 272
use FILL  FILL_4__2109_
timestamp 1701859473
transform -1 0 3370 0 -1 790
box -12 -8 32 272
use FILL  FILL_4__2110_
timestamp 1701859473
transform 1 0 3130 0 -1 790
box -12 -8 32 272
use FILL  FILL_4__2111_
timestamp 1701859473
transform -1 0 3810 0 -1 790
box -12 -8 32 272
use FILL  FILL_4__2112_
timestamp 1701859473
transform -1 0 5170 0 -1 790
box -12 -8 32 272
use FILL  FILL_4__2113_
timestamp 1701859473
transform -1 0 5150 0 1 1310
box -12 -8 32 272
use FILL  FILL_4__2114_
timestamp 1701859473
transform -1 0 5590 0 1 1310
box -12 -8 32 272
use FILL  FILL_4__2115_
timestamp 1701859473
transform -1 0 5630 0 -1 790
box -12 -8 32 272
use FILL  FILL_4__2116_
timestamp 1701859473
transform 1 0 2450 0 1 1310
box -12 -8 32 272
use FILL  FILL_4__2117_
timestamp 1701859473
transform 1 0 2650 0 1 1310
box -12 -8 32 272
use FILL  FILL_4__2118_
timestamp 1701859473
transform 1 0 3830 0 1 1310
box -12 -8 32 272
use FILL  FILL_4__2119_
timestamp 1701859473
transform -1 0 4090 0 1 1310
box -12 -8 32 272
use FILL  FILL_4__2120_
timestamp 1701859473
transform 1 0 3950 0 -1 1310
box -12 -8 32 272
use FILL  FILL_4__2121_
timestamp 1701859473
transform -1 0 4530 0 1 270
box -12 -8 32 272
use FILL  FILL_4__2122_
timestamp 1701859473
transform -1 0 2870 0 1 2350
box -12 -8 32 272
use FILL  FILL_4__2123_
timestamp 1701859473
transform 1 0 2810 0 -1 2350
box -12 -8 32 272
use FILL  FILL_4__2124_
timestamp 1701859473
transform -1 0 3710 0 -1 2350
box -12 -8 32 272
use FILL  FILL_4__2125_
timestamp 1701859473
transform 1 0 5830 0 -1 3390
box -12 -8 32 272
use FILL  FILL_4__2126_
timestamp 1701859473
transform 1 0 5510 0 1 2870
box -12 -8 32 272
use FILL  FILL_4__2127_
timestamp 1701859473
transform -1 0 5990 0 1 2870
box -12 -8 32 272
use FILL  FILL_4__2128_
timestamp 1701859473
transform 1 0 4610 0 1 2870
box -12 -8 32 272
use FILL  FILL_4__2129_
timestamp 1701859473
transform 1 0 5290 0 1 2870
box -12 -8 32 272
use FILL  FILL_4__2130_
timestamp 1701859473
transform -1 0 4650 0 -1 2350
box -12 -8 32 272
use FILL  FILL_4__2131_
timestamp 1701859473
transform 1 0 4690 0 1 1310
box -12 -8 32 272
use FILL  FILL_4__2132_
timestamp 1701859473
transform -1 0 4570 0 1 790
box -12 -8 32 272
use FILL  FILL_4__2133_
timestamp 1701859473
transform 1 0 4490 0 -1 790
box -12 -8 32 272
use FILL  FILL_4__2134_
timestamp 1701859473
transform 1 0 3610 0 -1 2870
box -12 -8 32 272
use FILL  FILL_4__2135_
timestamp 1701859473
transform 1 0 4230 0 -1 3390
box -12 -8 32 272
use FILL  FILL_4__2136_
timestamp 1701859473
transform -1 0 2770 0 1 3390
box -12 -8 32 272
use FILL  FILL_4__2137_
timestamp 1701859473
transform 1 0 2330 0 1 3390
box -12 -8 32 272
use FILL  FILL_4__2138_
timestamp 1701859473
transform 1 0 3130 0 -1 4430
box -12 -8 32 272
use FILL  FILL_4__2139_
timestamp 1701859473
transform -1 0 2910 0 -1 4430
box -12 -8 32 272
use FILL  FILL_4__2140_
timestamp 1701859473
transform 1 0 2830 0 1 4430
box -12 -8 32 272
use FILL  FILL_4__2141_
timestamp 1701859473
transform -1 0 3070 0 1 4430
box -12 -8 32 272
use FILL  FILL_4__2142_
timestamp 1701859473
transform 1 0 2950 0 1 3390
box -12 -8 32 272
use FILL  FILL_4__2143_
timestamp 1701859473
transform -1 0 7450 0 -1 3390
box -12 -8 32 272
use FILL  FILL_4__2144_
timestamp 1701859473
transform 1 0 2090 0 1 2870
box -12 -8 32 272
use FILL  FILL_4__2145_
timestamp 1701859473
transform -1 0 10070 0 -1 2870
box -12 -8 32 272
use FILL  FILL_4__2146_
timestamp 1701859473
transform -1 0 7650 0 -1 3390
box -12 -8 32 272
use FILL  FILL_4__2147_
timestamp 1701859473
transform 1 0 7610 0 -1 3910
box -12 -8 32 272
use FILL  FILL_4__2148_
timestamp 1701859473
transform 1 0 7450 0 1 3390
box -12 -8 32 272
use FILL  FILL_4__2149_
timestamp 1701859473
transform 1 0 7650 0 1 3390
box -12 -8 32 272
use FILL  FILL_4__2150_
timestamp 1701859473
transform -1 0 7910 0 1 3390
box -12 -8 32 272
use FILL  FILL_4__2151_
timestamp 1701859473
transform 1 0 7190 0 -1 3390
box -12 -8 32 272
use FILL  FILL_4__2152_
timestamp 1701859473
transform 1 0 6950 0 -1 3390
box -12 -8 32 272
use FILL  FILL_4__2153_
timestamp 1701859473
transform -1 0 6090 0 -1 3390
box -12 -8 32 272
use FILL  FILL_4__2154_
timestamp 1701859473
transform 1 0 2850 0 -1 7030
box -12 -8 32 272
use FILL  FILL_4__2155_
timestamp 1701859473
transform 1 0 6410 0 1 5990
box -12 -8 32 272
use FILL  FILL_4__2156_
timestamp 1701859473
transform -1 0 4630 0 1 3910
box -12 -8 32 272
use FILL  FILL_4__2157_
timestamp 1701859473
transform -1 0 4770 0 -1 4430
box -12 -8 32 272
use FILL  FILL_4__2158_
timestamp 1701859473
transform -1 0 2630 0 1 2350
box -12 -8 32 272
use FILL  FILL_4__2159_
timestamp 1701859473
transform 1 0 3530 0 1 3910
box -12 -8 32 272
use FILL  FILL_4__2160_
timestamp 1701859473
transform -1 0 3850 0 -1 4430
box -12 -8 32 272
use FILL  FILL_4__2161_
timestamp 1701859473
transform -1 0 3990 0 1 3910
box -12 -8 32 272
use FILL  FILL_4__2162_
timestamp 1701859473
transform -1 0 4430 0 1 3910
box -12 -8 32 272
use FILL  FILL_4__2163_
timestamp 1701859473
transform 1 0 3750 0 -1 3910
box -12 -8 32 272
use FILL  FILL_4__2164_
timestamp 1701859473
transform -1 0 570 0 -1 4950
box -12 -8 32 272
use FILL  FILL_4__2165_
timestamp 1701859473
transform -1 0 3270 0 -1 3910
box -12 -8 32 272
use FILL  FILL_4__2166_
timestamp 1701859473
transform 1 0 3970 0 -1 3910
box -12 -8 32 272
use FILL  FILL_4__2167_
timestamp 1701859473
transform 1 0 4170 0 1 3910
box -12 -8 32 272
use FILL  FILL_4__2168_
timestamp 1701859473
transform 1 0 3090 0 1 3910
box -12 -8 32 272
use FILL  FILL_4__2169_
timestamp 1701859473
transform 1 0 2450 0 -1 4430
box -12 -8 32 272
use FILL  FILL_4__2170_
timestamp 1701859473
transform -1 0 2710 0 -1 4430
box -12 -8 32 272
use FILL  FILL_4__2171_
timestamp 1701859473
transform 1 0 4050 0 -1 4430
box -12 -8 32 272
use FILL  FILL_4__2172_
timestamp 1701859473
transform 1 0 4290 0 -1 4430
box -12 -8 32 272
use FILL  FILL_4__2173_
timestamp 1701859473
transform -1 0 4530 0 -1 4430
box -12 -8 32 272
use FILL  FILL_4__2174_
timestamp 1701859473
transform 1 0 6030 0 1 7030
box -12 -8 32 272
use FILL  FILL_4__2175_
timestamp 1701859473
transform -1 0 2530 0 1 8070
box -12 -8 32 272
use FILL  FILL_4__2176_
timestamp 1701859473
transform -1 0 6450 0 -1 8070
box -12 -8 32 272
use FILL  FILL_4__2177_
timestamp 1701859473
transform 1 0 4970 0 1 8070
box -12 -8 32 272
use FILL  FILL_4__2178_
timestamp 1701859473
transform -1 0 4150 0 -1 8590
box -12 -8 32 272
use FILL  FILL_4__2179_
timestamp 1701859473
transform -1 0 5970 0 -1 8070
box -12 -8 32 272
use FILL  FILL_4__2180_
timestamp 1701859473
transform -1 0 2990 0 -1 9630
box -12 -8 32 272
use FILL  FILL_4__2181_
timestamp 1701859473
transform 1 0 5050 0 1 7550
box -12 -8 32 272
use FILL  FILL_4__2182_
timestamp 1701859473
transform 1 0 5570 0 -1 10150
box -12 -8 32 272
use FILL  FILL_4__2183_
timestamp 1701859473
transform -1 0 3550 0 1 10150
box -12 -8 32 272
use FILL  FILL_4__2184_
timestamp 1701859473
transform 1 0 4370 0 1 8070
box -12 -8 32 272
use FILL  FILL_4__2185_
timestamp 1701859473
transform 1 0 5970 0 1 10150
box -12 -8 32 272
use FILL  FILL_4__2186_
timestamp 1701859473
transform 1 0 3530 0 1 10670
box -12 -8 32 272
use FILL  FILL_4__2187_
timestamp 1701859473
transform -1 0 5450 0 -1 10670
box -12 -8 32 272
use FILL  FILL_4__2188_
timestamp 1701859473
transform 1 0 2130 0 -1 10670
box -12 -8 32 272
use FILL  FILL_4__2189_
timestamp 1701859473
transform 1 0 5690 0 -1 10670
box -12 -8 32 272
use FILL  FILL_4__2190_
timestamp 1701859473
transform -1 0 2850 0 1 10150
box -12 -8 32 272
use FILL  FILL_4__2191_
timestamp 1701859473
transform -1 0 5330 0 -1 10150
box -12 -8 32 272
use FILL  FILL_4__2192_
timestamp 1701859473
transform -1 0 11130 0 1 3910
box -12 -8 32 272
use FILL  FILL_4__2193_
timestamp 1701859473
transform 1 0 1250 0 -1 3910
box -12 -8 32 272
use FILL  FILL_4__2194_
timestamp 1701859473
transform 1 0 1050 0 -1 3910
box -12 -8 32 272
use FILL  FILL_4__2195_
timestamp 1701859473
transform 1 0 2630 0 1 3910
box -12 -8 32 272
use FILL  FILL_4__2196_
timestamp 1701859473
transform 1 0 2870 0 1 3910
box -12 -8 32 272
use FILL  FILL_4__2197_
timestamp 1701859473
transform 1 0 5350 0 1 3910
box -12 -8 32 272
use FILL  FILL_4__2198_
timestamp 1701859473
transform 1 0 290 0 1 1830
box -12 -8 32 272
use FILL  FILL_4__2199_
timestamp 1701859473
transform -1 0 2850 0 -1 3910
box -12 -8 32 272
use FILL  FILL_4__2200_
timestamp 1701859473
transform 1 0 5370 0 -1 3910
box -12 -8 32 272
use FILL  FILL_4__2201_
timestamp 1701859473
transform -1 0 5610 0 1 3910
box -12 -8 32 272
use FILL  FILL_4__2202_
timestamp 1701859473
transform -1 0 8190 0 -1 4430
box -12 -8 32 272
use FILL  FILL_4__2203_
timestamp 1701859473
transform -1 0 4910 0 -1 3910
box -12 -8 32 272
use FILL  FILL_4__2204_
timestamp 1701859473
transform 1 0 5130 0 -1 3910
box -12 -8 32 272
use FILL  FILL_4__2205_
timestamp 1701859473
transform -1 0 8990 0 -1 3910
box -12 -8 32 272
use FILL  FILL_4__2206_
timestamp 1701859473
transform 1 0 9070 0 1 3910
box -12 -8 32 272
use FILL  FILL_4__2207_
timestamp 1701859473
transform 1 0 9530 0 -1 3910
box -12 -8 32 272
use FILL  FILL_4__2208_
timestamp 1701859473
transform -1 0 9790 0 -1 3910
box -12 -8 32 272
use FILL  FILL_4__2209_
timestamp 1701859473
transform -1 0 9590 0 1 4430
box -12 -8 32 272
use FILL  FILL_4__2210_
timestamp 1701859473
transform -1 0 10590 0 -1 4950
box -12 -8 32 272
use FILL  FILL_4__2211_
timestamp 1701859473
transform 1 0 9290 0 -1 3910
box -12 -8 32 272
use FILL  FILL_4__2212_
timestamp 1701859473
transform -1 0 8870 0 1 3910
box -12 -8 32 272
use FILL  FILL_4__2213_
timestamp 1701859473
transform -1 0 9310 0 1 3910
box -12 -8 32 272
use FILL  FILL_4__2214_
timestamp 1701859473
transform -1 0 9510 0 -1 4430
box -12 -8 32 272
use FILL  FILL_4__2215_
timestamp 1701859473
transform 1 0 9710 0 -1 4430
box -12 -8 32 272
use FILL  FILL_4__2216_
timestamp 1701859473
transform -1 0 9470 0 -1 7030
box -12 -8 32 272
use FILL  FILL_4__2217_
timestamp 1701859473
transform 1 0 9250 0 -1 4430
box -12 -8 32 272
use FILL  FILL_4__2218_
timestamp 1701859473
transform -1 0 9770 0 1 3910
box -12 -8 32 272
use FILL  FILL_4__2219_
timestamp 1701859473
transform 1 0 9950 0 1 3910
box -12 -8 32 272
use FILL  FILL_4__2220_
timestamp 1701859473
transform 1 0 10330 0 -1 4950
box -12 -8 32 272
use FILL  FILL_4__2221_
timestamp 1701859473
transform -1 0 9710 0 -1 7030
box -12 -8 32 272
use FILL  FILL_4__2222_
timestamp 1701859473
transform 1 0 10070 0 1 4430
box -12 -8 32 272
use FILL  FILL_4__2223_
timestamp 1701859473
transform -1 0 9970 0 -1 4430
box -12 -8 32 272
use FILL  FILL_4__2224_
timestamp 1701859473
transform -1 0 9830 0 1 4430
box -12 -8 32 272
use FILL  FILL_4__2225_
timestamp 1701859473
transform 1 0 10070 0 -1 4950
box -12 -8 32 272
use FILL  FILL_4__2226_
timestamp 1701859473
transform 1 0 8950 0 -1 7030
box -12 -8 32 272
use FILL  FILL_4__2227_
timestamp 1701859473
transform -1 0 9230 0 -1 7030
box -12 -8 32 272
use FILL  FILL_4__2228_
timestamp 1701859473
transform -1 0 5770 0 -1 7030
box -12 -8 32 272
use FILL  FILL_4__2229_
timestamp 1701859473
transform 1 0 4330 0 1 3390
box -12 -8 32 272
use FILL  FILL_4__2230_
timestamp 1701859473
transform -1 0 4430 0 -1 3910
box -12 -8 32 272
use FILL  FILL_4__2231_
timestamp 1701859473
transform -1 0 4210 0 -1 3910
box -12 -8 32 272
use FILL  FILL_4__2232_
timestamp 1701859473
transform 1 0 1610 0 1 2870
box -12 -8 32 272
use FILL  FILL_4__2233_
timestamp 1701859473
transform 1 0 2330 0 1 2870
box -12 -8 32 272
use FILL  FILL_4__2234_
timestamp 1701859473
transform -1 0 2590 0 1 2870
box -12 -8 32 272
use FILL  FILL_4__2235_
timestamp 1701859473
transform 1 0 6350 0 1 3390
box -12 -8 32 272
use FILL  FILL_4__2236_
timestamp 1701859473
transform -1 0 5630 0 -1 3910
box -12 -8 32 272
use FILL  FILL_4__2237_
timestamp 1701859473
transform -1 0 4670 0 -1 3910
box -12 -8 32 272
use FILL  FILL_4__2238_
timestamp 1701859473
transform 1 0 4730 0 -1 4950
box -12 -8 32 272
use FILL  FILL_4__2239_
timestamp 1701859473
transform 1 0 2850 0 1 4950
box -12 -8 32 272
use FILL  FILL_4__2240_
timestamp 1701859473
transform 1 0 2410 0 1 3910
box -12 -8 32 272
use FILL  FILL_4__2241_
timestamp 1701859473
transform -1 0 2430 0 1 4950
box -12 -8 32 272
use FILL  FILL_4__2242_
timestamp 1701859473
transform 1 0 2470 0 -1 4950
box -12 -8 32 272
use FILL  FILL_4__2243_
timestamp 1701859473
transform 1 0 2650 0 1 4950
box -12 -8 32 272
use FILL  FILL_4__2244_
timestamp 1701859473
transform 1 0 3070 0 1 4950
box -12 -8 32 272
use FILL  FILL_4__2245_
timestamp 1701859473
transform 1 0 2910 0 1 5990
box -12 -8 32 272
use FILL  FILL_4__2246_
timestamp 1701859473
transform 1 0 2930 0 -1 4950
box -12 -8 32 272
use FILL  FILL_4__2247_
timestamp 1701859473
transform -1 0 3050 0 -1 6510
box -12 -8 32 272
use FILL  FILL_4__2248_
timestamp 1701859473
transform 1 0 3510 0 -1 7030
box -12 -8 32 272
use FILL  FILL_4__2249_
timestamp 1701859473
transform 1 0 6290 0 1 7030
box -12 -8 32 272
use FILL  FILL_4__2250_
timestamp 1701859473
transform -1 0 10590 0 -1 7550
box -12 -8 32 272
use FILL  FILL_4__2251_
timestamp 1701859473
transform -1 0 10650 0 1 8070
box -12 -8 32 272
use FILL  FILL_4__2252_
timestamp 1701859473
transform -1 0 10950 0 -1 8070
box -12 -8 32 272
use FILL  FILL_4__2253_
timestamp 1701859473
transform -1 0 10710 0 -1 8070
box -12 -8 32 272
use FILL  FILL_4__2254_
timestamp 1701859473
transform 1 0 5410 0 1 8070
box -12 -8 32 272
use FILL  FILL_4__2255_
timestamp 1701859473
transform 1 0 3030 0 1 7030
box -12 -8 32 272
use FILL  FILL_4__2256_
timestamp 1701859473
transform -1 0 5150 0 1 7030
box -12 -8 32 272
use FILL  FILL_4__2257_
timestamp 1701859473
transform 1 0 5090 0 -1 7550
box -12 -8 32 272
use FILL  FILL_4__2258_
timestamp 1701859473
transform 1 0 5730 0 -1 8590
box -12 -8 32 272
use FILL  FILL_4__2259_
timestamp 1701859473
transform 1 0 10350 0 -1 7550
box -12 -8 32 272
use FILL  FILL_4__2260_
timestamp 1701859473
transform 1 0 9930 0 1 8070
box -12 -8 32 272
use FILL  FILL_4__2261_
timestamp 1701859473
transform -1 0 10230 0 1 7550
box -12 -8 32 272
use FILL  FILL_4__2262_
timestamp 1701859473
transform -1 0 9990 0 1 7550
box -12 -8 32 272
use FILL  FILL_4__2263_
timestamp 1701859473
transform 1 0 5490 0 1 7550
box -12 -8 32 272
use FILL  FILL_4__2264_
timestamp 1701859473
transform 1 0 1650 0 -1 6510
box -12 -8 32 272
use FILL  FILL_4__2265_
timestamp 1701859473
transform 1 0 1830 0 -1 6510
box -12 -8 32 272
use FILL  FILL_4__2266_
timestamp 1701859473
transform 1 0 3930 0 1 6510
box -12 -8 32 272
use FILL  FILL_4__2267_
timestamp 1701859473
transform -1 0 3690 0 -1 7550
box -12 -8 32 272
use FILL  FILL_4__2268_
timestamp 1701859473
transform 1 0 4370 0 -1 7550
box -12 -8 32 272
use FILL  FILL_4__2269_
timestamp 1701859473
transform 1 0 5690 0 1 7550
box -12 -8 32 272
use FILL  FILL_4__2270_
timestamp 1701859473
transform 1 0 8610 0 1 7550
box -12 -8 32 272
use FILL  FILL_4__2271_
timestamp 1701859473
transform -1 0 8890 0 -1 8070
box -12 -8 32 272
use FILL  FILL_4__2272_
timestamp 1701859473
transform -1 0 9150 0 -1 8070
box -12 -8 32 272
use FILL  FILL_4__2273_
timestamp 1701859473
transform -1 0 8650 0 -1 8070
box -12 -8 32 272
use FILL  FILL_4__2274_
timestamp 1701859473
transform -1 0 6010 0 -1 9630
box -12 -8 32 272
use FILL  FILL_4__2275_
timestamp 1701859473
transform -1 0 2310 0 1 8070
box -12 -8 32 272
use FILL  FILL_4__2276_
timestamp 1701859473
transform -1 0 3190 0 1 8070
box -12 -8 32 272
use FILL  FILL_4__2277_
timestamp 1701859473
transform -1 0 3670 0 -1 8590
box -12 -8 32 272
use FILL  FILL_4__2278_
timestamp 1701859473
transform 1 0 6570 0 1 9110
box -12 -8 32 272
use FILL  FILL_4__2279_
timestamp 1701859473
transform -1 0 10270 0 1 5990
box -12 -8 32 272
use FILL  FILL_4__2280_
timestamp 1701859473
transform 1 0 10450 0 1 5990
box -12 -8 32 272
use FILL  FILL_4__2281_
timestamp 1701859473
transform -1 0 10730 0 -1 5990
box -12 -8 32 272
use FILL  FILL_4__2282_
timestamp 1701859473
transform -1 0 10510 0 -1 6510
box -12 -8 32 272
use FILL  FILL_4__2283_
timestamp 1701859473
transform 1 0 5970 0 -1 8590
box -12 -8 32 272
use FILL  FILL_4__2284_
timestamp 1701859473
transform -1 0 2090 0 1 8070
box -12 -8 32 272
use FILL  FILL_4__2285_
timestamp 1701859473
transform -1 0 4150 0 1 8070
box -12 -8 32 272
use FILL  FILL_4__2286_
timestamp 1701859473
transform 1 0 5050 0 -1 8590
box -12 -8 32 272
use FILL  FILL_4__2287_
timestamp 1701859473
transform -1 0 6130 0 1 8590
box -12 -8 32 272
use FILL  FILL_4__2288_
timestamp 1701859473
transform -1 0 8850 0 1 7550
box -12 -8 32 272
use FILL  FILL_4__2289_
timestamp 1701859473
transform 1 0 8510 0 1 8070
box -12 -8 32 272
use FILL  FILL_4__2290_
timestamp 1701859473
transform -1 0 10010 0 -1 8070
box -12 -8 32 272
use FILL  FILL_4__2291_
timestamp 1701859473
transform -1 0 8790 0 1 8070
box -12 -8 32 272
use FILL  FILL_4__2292_
timestamp 1701859473
transform -1 0 6230 0 -1 9110
box -12 -8 32 272
use FILL  FILL_4__2293_
timestamp 1701859473
transform -1 0 2550 0 -1 8590
box -12 -8 32 272
use FILL  FILL_4__2294_
timestamp 1701859473
transform -1 0 4030 0 1 8590
box -12 -8 32 272
use FILL  FILL_4__2295_
timestamp 1701859473
transform 1 0 4950 0 1 8590
box -12 -8 32 272
use FILL  FILL_4__2296_
timestamp 1701859473
transform 1 0 6670 0 -1 9110
box -12 -8 32 272
use FILL  FILL_4__2297_
timestamp 1701859473
transform -1 0 9570 0 -1 5990
box -12 -8 32 272
use FILL  FILL_4__2298_
timestamp 1701859473
transform -1 0 10010 0 -1 5470
box -12 -8 32 272
use FILL  FILL_4__2299_
timestamp 1701859473
transform -1 0 9350 0 -1 6510
box -12 -8 32 272
use FILL  FILL_4__2300_
timestamp 1701859473
transform 1 0 9550 0 1 5990
box -12 -8 32 272
use FILL  FILL_4__2301_
timestamp 1701859473
transform 1 0 5590 0 1 9630
box -12 -8 32 272
use FILL  FILL_4__2302_
timestamp 1701859473
transform -1 0 3490 0 -1 9110
box -12 -8 32 272
use FILL  FILL_4__2303_
timestamp 1701859473
transform 1 0 2610 0 1 9110
box -12 -8 32 272
use FILL  FILL_4__2304_
timestamp 1701859473
transform 1 0 2810 0 -1 9110
box -12 -8 32 272
use FILL  FILL_4__2305_
timestamp 1701859473
transform -1 0 3790 0 1 8590
box -12 -8 32 272
use FILL  FILL_4__2306_
timestamp 1701859473
transform 1 0 4470 0 1 8590
box -12 -8 32 272
use FILL  FILL_4__2307_
timestamp 1701859473
transform 1 0 6330 0 1 9110
box -12 -8 32 272
use FILL  FILL_4__2308_
timestamp 1701859473
transform -1 0 8910 0 -1 6510
box -12 -8 32 272
use FILL  FILL_4__2309_
timestamp 1701859473
transform -1 0 8610 0 1 5990
box -12 -8 32 272
use FILL  FILL_4__2310_
timestamp 1701859473
transform -1 0 9110 0 -1 6510
box -12 -8 32 272
use FILL  FILL_4__2311_
timestamp 1701859473
transform -1 0 8670 0 -1 6510
box -12 -8 32 272
use FILL  FILL_4__2312_
timestamp 1701859473
transform -1 0 5570 0 -1 9630
box -12 -8 32 272
use FILL  FILL_4__2313_
timestamp 1701859473
transform -1 0 1850 0 1 8590
box -12 -8 32 272
use FILL  FILL_4__2314_
timestamp 1701859473
transform 1 0 1450 0 -1 8590
box -12 -8 32 272
use FILL  FILL_4__2315_
timestamp 1701859473
transform 1 0 1890 0 -1 8590
box -12 -8 32 272
use FILL  FILL_4__2316_
timestamp 1701859473
transform -1 0 4250 0 1 8590
box -12 -8 32 272
use FILL  FILL_4__2317_
timestamp 1701859473
transform 1 0 4710 0 1 8590
box -12 -8 32 272
use FILL  FILL_4__2318_
timestamp 1701859473
transform 1 0 6810 0 1 9110
box -12 -8 32 272
use FILL  FILL_4__2319_
timestamp 1701859473
transform -1 0 11130 0 1 4430
box -12 -8 32 272
use FILL  FILL_4__2320_
timestamp 1701859473
transform 1 0 5110 0 1 3910
box -12 -8 32 272
use FILL  FILL_4__2321_
timestamp 1701859473
transform 1 0 6530 0 1 3910
box -12 -8 32 272
use FILL  FILL_4__2322_
timestamp 1701859473
transform -1 0 7910 0 1 3910
box -12 -8 32 272
use FILL  FILL_4__2323_
timestamp 1701859473
transform 1 0 7950 0 -1 4430
box -12 -8 32 272
use FILL  FILL_4__2324_
timestamp 1701859473
transform -1 0 11170 0 -1 2870
box -12 -8 32 272
use FILL  FILL_4__2325_
timestamp 1701859473
transform -1 0 8150 0 1 3910
box -12 -8 32 272
use FILL  FILL_4__2326_
timestamp 1701859473
transform -1 0 3190 0 -1 4950
box -12 -8 32 272
use FILL  FILL_4__2327_
timestamp 1701859473
transform -1 0 3390 0 -1 4950
box -12 -8 32 272
use FILL  FILL_4__2328_
timestamp 1701859473
transform 1 0 3870 0 -1 5470
box -12 -8 32 272
use FILL  FILL_4__2329_
timestamp 1701859473
transform 1 0 3630 0 -1 5470
box -12 -8 32 272
use FILL  FILL_4__2330_
timestamp 1701859473
transform 1 0 3770 0 1 4950
box -12 -8 32 272
use FILL  FILL_4__2331_
timestamp 1701859473
transform 1 0 4850 0 1 3910
box -12 -8 32 272
use FILL  FILL_4__2332_
timestamp 1701859473
transform -1 0 4190 0 1 4950
box -12 -8 32 272
use FILL  FILL_4__2333_
timestamp 1701859473
transform -1 0 11150 0 -1 4430
box -12 -8 32 272
use FILL  FILL_4__2334_
timestamp 1701859473
transform 1 0 9030 0 -1 4430
box -12 -8 32 272
use FILL  FILL_4__2335_
timestamp 1701859473
transform 1 0 5210 0 -1 5470
box -12 -8 32 272
use FILL  FILL_4__2336_
timestamp 1701859473
transform -1 0 5070 0 1 5990
box -12 -8 32 272
use FILL  FILL_4__2337_
timestamp 1701859473
transform 1 0 4570 0 1 3390
box -12 -8 32 272
use FILL  FILL_4__2338_
timestamp 1701859473
transform 1 0 3170 0 1 3390
box -12 -8 32 272
use FILL  FILL_4__2339_
timestamp 1701859473
transform 1 0 4750 0 1 3390
box -12 -8 32 272
use FILL  FILL_4__2340_
timestamp 1701859473
transform 1 0 4990 0 1 3390
box -12 -8 32 272
use FILL  FILL_4__2341_
timestamp 1701859473
transform -1 0 570 0 1 5990
box -12 -8 32 272
use FILL  FILL_4__2342_
timestamp 1701859473
transform 1 0 2670 0 1 5470
box -12 -8 32 272
use FILL  FILL_4__2343_
timestamp 1701859473
transform -1 0 4610 0 1 6510
box -12 -8 32 272
use FILL  FILL_4__2344_
timestamp 1701859473
transform -1 0 4890 0 1 5470
box -12 -8 32 272
use FILL  FILL_4__2345_
timestamp 1701859473
transform -1 0 4690 0 1 5470
box -12 -8 32 272
use FILL  FILL_4__2346_
timestamp 1701859473
transform -1 0 4850 0 -1 5990
box -12 -8 32 272
use FILL  FILL_4__2347_
timestamp 1701859473
transform -1 0 5710 0 -1 5990
box -12 -8 32 272
use FILL  FILL_4__2348_
timestamp 1701859473
transform 1 0 5270 0 -1 6510
box -12 -8 32 272
use FILL  FILL_4__2349_
timestamp 1701859473
transform -1 0 5050 0 -1 6510
box -12 -8 32 272
use FILL  FILL_4__2350_
timestamp 1701859473
transform -1 0 4470 0 -1 6510
box -12 -8 32 272
use FILL  FILL_4__2351_
timestamp 1701859473
transform 1 0 5610 0 1 7030
box -12 -8 32 272
use FILL  FILL_4__2352_
timestamp 1701859473
transform -1 0 5830 0 1 7030
box -12 -8 32 272
use FILL  FILL_4__2353_
timestamp 1701859473
transform -1 0 770 0 1 7030
box -12 -8 32 272
use FILL  FILL_4__2354_
timestamp 1701859473
transform 1 0 5470 0 -1 5990
box -12 -8 32 272
use FILL  FILL_4__2355_
timestamp 1701859473
transform 1 0 5370 0 1 7030
box -12 -8 32 272
use FILL  FILL_4__2356_
timestamp 1701859473
transform -1 0 4870 0 -1 7550
box -12 -8 32 272
use FILL  FILL_4__2357_
timestamp 1701859473
transform 1 0 4730 0 1 8070
box -12 -8 32 272
use FILL  FILL_4__2358_
timestamp 1701859473
transform 1 0 5210 0 1 8070
box -12 -8 32 272
use FILL  FILL_4__2359_
timestamp 1701859473
transform -1 0 5530 0 -1 8590
box -12 -8 32 272
use FILL  FILL_4__2360_
timestamp 1701859473
transform -1 0 770 0 -1 6510
box -12 -8 32 272
use FILL  FILL_4__2361_
timestamp 1701859473
transform -1 0 5270 0 1 5990
box -12 -8 32 272
use FILL  FILL_4__2362_
timestamp 1701859473
transform 1 0 5270 0 1 6510
box -12 -8 32 272
use FILL  FILL_4__2363_
timestamp 1701859473
transform 1 0 5290 0 -1 7030
box -12 -8 32 272
use FILL  FILL_4__2364_
timestamp 1701859473
transform 1 0 5290 0 -1 8070
box -12 -8 32 272
use FILL  FILL_4__2365_
timestamp 1701859473
transform 1 0 5530 0 -1 8070
box -12 -8 32 272
use FILL  FILL_4__2366_
timestamp 1701859473
transform -1 0 5750 0 -1 8070
box -12 -8 32 272
use FILL  FILL_4__2367_
timestamp 1701859473
transform 1 0 2710 0 -1 7550
box -12 -8 32 272
use FILL  FILL_4__2368_
timestamp 1701859473
transform -1 0 5550 0 -1 7030
box -12 -8 32 272
use FILL  FILL_4__2369_
timestamp 1701859473
transform 1 0 5250 0 1 7550
box -12 -8 32 272
use FILL  FILL_4__2370_
timestamp 1701859473
transform -1 0 5290 0 -1 8590
box -12 -8 32 272
use FILL  FILL_4__2371_
timestamp 1701859473
transform 1 0 5970 0 -1 9110
box -12 -8 32 272
use FILL  FILL_4__2372_
timestamp 1701859473
transform 1 0 6130 0 1 9110
box -12 -8 32 272
use FILL  FILL_4__2373_
timestamp 1701859473
transform -1 0 6210 0 -1 9630
box -12 -8 32 272
use FILL  FILL_4__2374_
timestamp 1701859473
transform 1 0 90 0 -1 9110
box -12 -8 32 272
use FILL  FILL_4__2375_
timestamp 1701859473
transform -1 0 4230 0 1 5470
box -12 -8 32 272
use FILL  FILL_4__2376_
timestamp 1701859473
transform 1 0 4570 0 -1 5990
box -12 -8 32 272
use FILL  FILL_4__2377_
timestamp 1701859473
transform -1 0 3990 0 -1 6510
box -12 -8 32 272
use FILL  FILL_4__2378_
timestamp 1701859473
transform 1 0 3730 0 -1 6510
box -12 -8 32 272
use FILL  FILL_4__2379_
timestamp 1701859473
transform -1 0 5050 0 1 6510
box -12 -8 32 272
use FILL  FILL_4__2380_
timestamp 1701859473
transform -1 0 4830 0 -1 8590
box -12 -8 32 272
use FILL  FILL_4__2381_
timestamp 1701859473
transform 1 0 3890 0 -1 8590
box -12 -8 32 272
use FILL  FILL_4__2382_
timestamp 1701859473
transform -1 0 4590 0 -1 8590
box -12 -8 32 272
use FILL  FILL_4__2383_
timestamp 1701859473
transform -1 0 5670 0 1 8590
box -12 -8 32 272
use FILL  FILL_4__2384_
timestamp 1701859473
transform -1 0 5890 0 1 8590
box -12 -8 32 272
use FILL  FILL_4__2385_
timestamp 1701859473
transform 1 0 1270 0 -1 10150
box -12 -8 32 272
use FILL  FILL_4__2386_
timestamp 1701859473
transform 1 0 5530 0 -1 7550
box -12 -8 32 272
use FILL  FILL_4__2387_
timestamp 1701859473
transform 1 0 5510 0 -1 9110
box -12 -8 32 272
use FILL  FILL_4__2388_
timestamp 1701859473
transform -1 0 5310 0 -1 9110
box -12 -8 32 272
use FILL  FILL_4__2389_
timestamp 1701859473
transform -1 0 5090 0 -1 9630
box -12 -8 32 272
use FILL  FILL_4__2390_
timestamp 1701859473
transform 1 0 5150 0 1 9630
box -12 -8 32 272
use FILL  FILL_4__2391_
timestamp 1701859473
transform -1 0 5370 0 1 9630
box -12 -8 32 272
use FILL  FILL_4__2392_
timestamp 1701859473
transform 1 0 1470 0 -1 10150
box -12 -8 32 272
use FILL  FILL_4__2393_
timestamp 1701859473
transform -1 0 5330 0 -1 7550
box -12 -8 32 272
use FILL  FILL_4__2394_
timestamp 1701859473
transform 1 0 5410 0 1 8590
box -12 -8 32 272
use FILL  FILL_4__2395_
timestamp 1701859473
transform -1 0 5770 0 -1 9110
box -12 -8 32 272
use FILL  FILL_4__2396_
timestamp 1701859473
transform 1 0 5690 0 1 9110
box -12 -8 32 272
use FILL  FILL_4__2397_
timestamp 1701859473
transform 1 0 5930 0 1 9110
box -12 -8 32 272
use FILL  FILL_4__2398_
timestamp 1701859473
transform 1 0 5750 0 -1 9630
box -12 -8 32 272
use FILL  FILL_4__2399_
timestamp 1701859473
transform -1 0 3190 0 -1 5470
box -12 -8 32 272
use FILL  FILL_4__2400_
timestamp 1701859473
transform -1 0 3370 0 1 5990
box -12 -8 32 272
use FILL  FILL_4__2401_
timestamp 1701859473
transform 1 0 3290 0 -1 6510
box -12 -8 32 272
use FILL  FILL_4__2402_
timestamp 1701859473
transform -1 0 2230 0 -1 4430
box -12 -8 32 272
use FILL  FILL_4__2403_
timestamp 1701859473
transform -1 0 2630 0 1 4430
box -12 -8 32 272
use FILL  FILL_4__2404_
timestamp 1701859473
transform -1 0 2950 0 -1 5470
box -12 -8 32 272
use FILL  FILL_4__2405_
timestamp 1701859473
transform 1 0 2330 0 -1 2870
box -12 -8 32 272
use FILL  FILL_4__2406_
timestamp 1701859473
transform 1 0 3030 0 -1 3390
box -12 -8 32 272
use FILL  FILL_4__2407_
timestamp 1701859473
transform -1 0 3170 0 1 5470
box -12 -8 32 272
use FILL  FILL_4__2408_
timestamp 1701859473
transform 1 0 790 0 -1 2870
box -12 -8 32 272
use FILL  FILL_4__2409_
timestamp 1701859473
transform 1 0 810 0 -1 3910
box -12 -8 32 272
use FILL  FILL_4__2410_
timestamp 1701859473
transform 1 0 1210 0 1 4430
box -12 -8 32 272
use FILL  FILL_4__2411_
timestamp 1701859473
transform -1 0 770 0 -1 4950
box -12 -8 32 272
use FILL  FILL_4__2412_
timestamp 1701859473
transform 1 0 2450 0 -1 5990
box -12 -8 32 272
use FILL  FILL_4__2413_
timestamp 1701859473
transform 1 0 2910 0 1 5470
box -12 -8 32 272
use FILL  FILL_4__2414_
timestamp 1701859473
transform 1 0 4070 0 -1 5470
box -12 -8 32 272
use FILL  FILL_4__2415_
timestamp 1701859473
transform -1 0 4010 0 1 7030
box -12 -8 32 272
use FILL  FILL_4__2416_
timestamp 1701859473
transform 1 0 3970 0 1 4950
box -12 -8 32 272
use FILL  FILL_4__2417_
timestamp 1701859473
transform 1 0 4310 0 -1 5470
box -12 -8 32 272
use FILL  FILL_4__2418_
timestamp 1701859473
transform -1 0 1570 0 -1 4950
box -12 -8 32 272
use FILL  FILL_4__2419_
timestamp 1701859473
transform 1 0 2150 0 1 4430
box -12 -8 32 272
use FILL  FILL_4__2420_
timestamp 1701859473
transform 1 0 3810 0 1 5990
box -12 -8 32 272
use FILL  FILL_4__2421_
timestamp 1701859473
transform -1 0 3590 0 1 5990
box -12 -8 32 272
use FILL  FILL_4__2422_
timestamp 1701859473
transform -1 0 3470 0 -1 5990
box -12 -8 32 272
use FILL  FILL_4__2423_
timestamp 1701859473
transform -1 0 3690 0 -1 5990
box -12 -8 32 272
use FILL  FILL_4__2424_
timestamp 1701859473
transform 1 0 3230 0 -1 5990
box -12 -8 32 272
use FILL  FILL_4__2425_
timestamp 1701859473
transform 1 0 4370 0 1 5990
box -12 -8 32 272
use FILL  FILL_4__2426_
timestamp 1701859473
transform 1 0 3970 0 -1 7030
box -12 -8 32 272
use FILL  FILL_4__2427_
timestamp 1701859473
transform 1 0 4790 0 1 5990
box -12 -8 32 272
use FILL  FILL_4__2428_
timestamp 1701859473
transform 1 0 4550 0 1 5990
box -12 -8 32 272
use FILL  FILL_4__2429_
timestamp 1701859473
transform -1 0 4230 0 -1 6510
box -12 -8 32 272
use FILL  FILL_4__2430_
timestamp 1701859473
transform 1 0 4790 0 1 6510
box -12 -8 32 272
use FILL  FILL_4__2431_
timestamp 1701859473
transform -1 0 4890 0 -1 7030
box -12 -8 32 272
use FILL  FILL_4__2432_
timestamp 1701859473
transform 1 0 5110 0 -1 7030
box -12 -8 32 272
use FILL  FILL_4__2433_
timestamp 1701859473
transform -1 0 4370 0 -1 8070
box -12 -8 32 272
use FILL  FILL_4__2434_
timestamp 1701859473
transform 1 0 4850 0 1 7550
box -12 -8 32 272
use FILL  FILL_4__2435_
timestamp 1701859473
transform 1 0 4190 0 1 7030
box -12 -8 32 272
use FILL  FILL_4__2436_
timestamp 1701859473
transform -1 0 4630 0 -1 7550
box -12 -8 32 272
use FILL  FILL_4__2437_
timestamp 1701859473
transform -1 0 4610 0 -1 8070
box -12 -8 32 272
use FILL  FILL_4__2438_
timestamp 1701859473
transform -1 0 4850 0 -1 8070
box -12 -8 32 272
use FILL  FILL_4__2439_
timestamp 1701859473
transform -1 0 5090 0 -1 8070
box -12 -8 32 272
use FILL  FILL_4__2440_
timestamp 1701859473
transform 1 0 4630 0 1 10150
box -12 -8 32 272
use FILL  FILL_4__2441_
timestamp 1701859473
transform 1 0 3910 0 -1 7550
box -12 -8 32 272
use FILL  FILL_4__2442_
timestamp 1701859473
transform -1 0 4130 0 -1 8070
box -12 -8 32 272
use FILL  FILL_4__2443_
timestamp 1701859473
transform -1 0 3910 0 1 8070
box -12 -8 32 272
use FILL  FILL_4__2444_
timestamp 1701859473
transform 1 0 3650 0 1 8070
box -12 -8 32 272
use FILL  FILL_4__2445_
timestamp 1701859473
transform -1 0 4630 0 1 7550
box -12 -8 32 272
use FILL  FILL_4__2446_
timestamp 1701859473
transform 1 0 4550 0 1 8070
box -12 -8 32 272
use FILL  FILL_4__2447_
timestamp 1701859473
transform 1 0 4290 0 1 9110
box -12 -8 32 272
use FILL  FILL_4__2448_
timestamp 1701859473
transform 1 0 4950 0 1 9110
box -12 -8 32 272
use FILL  FILL_4__2449_
timestamp 1701859473
transform 1 0 5210 0 1 9110
box -12 -8 32 272
use FILL  FILL_4__2450_
timestamp 1701859473
transform 1 0 5450 0 1 9110
box -12 -8 32 272
use FILL  FILL_4__2451_
timestamp 1701859473
transform -1 0 5330 0 -1 9630
box -12 -8 32 272
use FILL  FILL_4__2452_
timestamp 1701859473
transform -1 0 5250 0 -1 10670
box -12 -8 32 272
use FILL  FILL_4__2453_
timestamp 1701859473
transform 1 0 3790 0 -1 10150
box -12 -8 32 272
use FILL  FILL_4__2454_
timestamp 1701859473
transform 1 0 3910 0 1 7550
box -12 -8 32 272
use FILL  FILL_4__2455_
timestamp 1701859473
transform 1 0 3870 0 -1 8070
box -12 -8 32 272
use FILL  FILL_4__2456_
timestamp 1701859473
transform -1 0 3650 0 -1 8070
box -12 -8 32 272
use FILL  FILL_4__2457_
timestamp 1701859473
transform 1 0 3410 0 1 8070
box -12 -8 32 272
use FILL  FILL_4__2458_
timestamp 1701859473
transform -1 0 4350 0 -1 8590
box -12 -8 32 272
use FILL  FILL_4__2459_
timestamp 1701859473
transform -1 0 4510 0 -1 11190
box -12 -8 32 272
use FILL  FILL_4__2460_
timestamp 1701859473
transform 1 0 4150 0 -1 10670
box -12 -8 32 272
use FILL  FILL_4__2461_
timestamp 1701859473
transform 1 0 4330 0 -1 9110
box -12 -8 32 272
use FILL  FILL_4__2462_
timestamp 1701859473
transform -1 0 4590 0 -1 9110
box -12 -8 32 272
use FILL  FILL_4__2463_
timestamp 1701859473
transform -1 0 4830 0 -1 9110
box -12 -8 32 272
use FILL  FILL_4__2464_
timestamp 1701859473
transform -1 0 5070 0 -1 9110
box -12 -8 32 272
use FILL  FILL_4__2465_
timestamp 1701859473
transform -1 0 4930 0 -1 11190
box -12 -8 32 272
use FILL  FILL_4__2466_
timestamp 1701859473
transform -1 0 4010 0 -1 10150
box -12 -8 32 272
use FILL  FILL_4__2467_
timestamp 1701859473
transform -1 0 4110 0 -1 9630
box -12 -8 32 272
use FILL  FILL_4__2468_
timestamp 1701859473
transform -1 0 4370 0 -1 9630
box -12 -8 32 272
use FILL  FILL_4__2469_
timestamp 1701859473
transform -1 0 4230 0 1 9630
box -12 -8 32 272
use FILL  FILL_4__2470_
timestamp 1701859473
transform -1 0 4470 0 1 9630
box -12 -8 32 272
use FILL  FILL_4__2471_
timestamp 1701859473
transform -1 0 5050 0 -1 10670
box -12 -8 32 272
use FILL  FILL_4__2472_
timestamp 1701859473
transform 1 0 4010 0 1 9630
box -12 -8 32 272
use FILL  FILL_4__2473_
timestamp 1701859473
transform 1 0 4570 0 -1 9630
box -12 -8 32 272
use FILL  FILL_4__2474_
timestamp 1701859473
transform -1 0 4850 0 -1 9630
box -12 -8 32 272
use FILL  FILL_4__2475_
timestamp 1701859473
transform 1 0 4690 0 1 9630
box -12 -8 32 272
use FILL  FILL_4__2476_
timestamp 1701859473
transform -1 0 4930 0 1 9630
box -12 -8 32 272
use FILL  FILL_4__2477_
timestamp 1701859473
transform 1 0 4870 0 1 10670
box -12 -8 32 272
use FILL  FILL_4__2478_
timestamp 1701859473
transform 1 0 3110 0 1 5990
box -12 -8 32 272
use FILL  FILL_4__2479_
timestamp 1701859473
transform -1 0 2670 0 1 5990
box -12 -8 32 272
use FILL  FILL_4__2480_
timestamp 1701859473
transform -1 0 2690 0 -1 5990
box -12 -8 32 272
use FILL  FILL_4__2481_
timestamp 1701859473
transform -1 0 2930 0 -1 5990
box -12 -8 32 272
use FILL  FILL_4__2482_
timestamp 1701859473
transform 1 0 1510 0 -1 5990
box -12 -8 32 272
use FILL  FILL_4__2483_
timestamp 1701859473
transform 1 0 2330 0 1 6510
box -12 -8 32 272
use FILL  FILL_4__2484_
timestamp 1701859473
transform -1 0 1950 0 1 6510
box -12 -8 32 272
use FILL  FILL_4__2485_
timestamp 1701859473
transform -1 0 2150 0 1 6510
box -12 -8 32 272
use FILL  FILL_4__2486_
timestamp 1701859473
transform 1 0 2350 0 -1 7030
box -12 -8 32 272
use FILL  FILL_4__2487_
timestamp 1701859473
transform 1 0 2110 0 -1 7030
box -12 -8 32 272
use FILL  FILL_4__2488_
timestamp 1701859473
transform -1 0 1910 0 -1 7030
box -12 -8 32 272
use FILL  FILL_4__2489_
timestamp 1701859473
transform 1 0 1410 0 -1 7030
box -12 -8 32 272
use FILL  FILL_4__2490_
timestamp 1701859473
transform -1 0 1010 0 1 5470
box -12 -8 32 272
use FILL  FILL_4__2491_
timestamp 1701859473
transform 1 0 1210 0 1 5470
box -12 -8 32 272
use FILL  FILL_4__2492_
timestamp 1701859473
transform -1 0 2070 0 -1 6510
box -12 -8 32 272
use FILL  FILL_4__2493_
timestamp 1701859473
transform 1 0 1950 0 1 5990
box -12 -8 32 272
use FILL  FILL_4__2494_
timestamp 1701859473
transform -1 0 1510 0 1 5990
box -12 -8 32 272
use FILL  FILL_4__2495_
timestamp 1701859473
transform 1 0 1250 0 1 5990
box -12 -8 32 272
use FILL  FILL_4__2496_
timestamp 1701859473
transform 1 0 1650 0 -1 7030
box -12 -8 32 272
use FILL  FILL_4__2497_
timestamp 1701859473
transform -1 0 1850 0 -1 7550
box -12 -8 32 272
use FILL  FILL_4__2498_
timestamp 1701859473
transform 1 0 790 0 1 8070
box -12 -8 32 272
use FILL  FILL_4__2499_
timestamp 1701859473
transform 1 0 2470 0 1 7550
box -12 -8 32 272
use FILL  FILL_4__2500_
timestamp 1701859473
transform 1 0 1890 0 1 7550
box -12 -8 32 272
use FILL  FILL_4__2501_
timestamp 1701859473
transform 1 0 1670 0 1 7550
box -12 -8 32 272
use FILL  FILL_4__2502_
timestamp 1701859473
transform -1 0 1210 0 1 7550
box -12 -8 32 272
use FILL  FILL_4__2503_
timestamp 1701859473
transform -1 0 1450 0 1 8070
box -12 -8 32 272
use FILL  FILL_4__2504_
timestamp 1701859473
transform -1 0 1870 0 1 8070
box -12 -8 32 272
use FILL  FILL_4__2505_
timestamp 1701859473
transform 1 0 1210 0 1 8070
box -12 -8 32 272
use FILL  FILL_4__2506_
timestamp 1701859473
transform -1 0 1730 0 -1 8070
box -12 -8 32 272
use FILL  FILL_4__2507_
timestamp 1701859473
transform 1 0 1470 0 -1 8070
box -12 -8 32 272
use FILL  FILL_4__2508_
timestamp 1701859473
transform 1 0 990 0 1 8070
box -12 -8 32 272
use FILL  FILL_4__2509_
timestamp 1701859473
transform 1 0 550 0 -1 8590
box -12 -8 32 272
use FILL  FILL_4__2510_
timestamp 1701859473
transform -1 0 1490 0 1 9110
box -12 -8 32 272
use FILL  FILL_4__2511_
timestamp 1701859473
transform -1 0 1430 0 -1 9630
box -12 -8 32 272
use FILL  FILL_4__2512_
timestamp 1701859473
transform 1 0 990 0 -1 9630
box -12 -8 32 272
use FILL  FILL_4__2513_
timestamp 1701859473
transform -1 0 990 0 1 8590
box -12 -8 32 272
use FILL  FILL_4__2514_
timestamp 1701859473
transform 1 0 2070 0 -1 8590
box -12 -8 32 272
use FILL  FILL_4__2515_
timestamp 1701859473
transform 1 0 1190 0 -1 9110
box -12 -8 32 272
use FILL  FILL_4__2516_
timestamp 1701859473
transform -1 0 1030 0 1 9110
box -12 -8 32 272
use FILL  FILL_4__2517_
timestamp 1701859473
transform -1 0 790 0 1 9110
box -12 -8 32 272
use FILL  FILL_4__2518_
timestamp 1701859473
transform 1 0 1650 0 -1 9630
box -12 -8 32 272
use FILL  FILL_4__2519_
timestamp 1701859473
transform 1 0 1750 0 1 9630
box -12 -8 32 272
use FILL  FILL_4__2520_
timestamp 1701859473
transform -1 0 2590 0 -1 9110
box -12 -8 32 272
use FILL  FILL_4__2521_
timestamp 1701859473
transform 1 0 2330 0 -1 9110
box -12 -8 32 272
use FILL  FILL_4__2522_
timestamp 1701859473
transform -1 0 1950 0 1 9630
box -12 -8 32 272
use FILL  FILL_4__2523_
timestamp 1701859473
transform -1 0 2170 0 1 9630
box -12 -8 32 272
use FILL  FILL_4__2524_
timestamp 1701859473
transform -1 0 1910 0 -1 9110
box -12 -8 32 272
use FILL  FILL_4__2525_
timestamp 1701859473
transform 1 0 790 0 -1 8590
box -12 -8 32 272
use FILL  FILL_4__2526_
timestamp 1701859473
transform -1 0 1690 0 -1 8590
box -12 -8 32 272
use FILL  FILL_4__2527_
timestamp 1701859473
transform -1 0 1230 0 -1 8590
box -12 -8 32 272
use FILL  FILL_4__2528_
timestamp 1701859473
transform -1 0 1010 0 -1 8590
box -12 -8 32 272
use FILL  FILL_4__2529_
timestamp 1701859473
transform -1 0 1250 0 1 9110
box -12 -8 32 272
use FILL  FILL_4__2530_
timestamp 1701859473
transform -1 0 7510 0 -1 6510
box -12 -8 32 272
use FILL  FILL_4__2531_
timestamp 1701859473
transform 1 0 7930 0 1 7550
box -12 -8 32 272
use FILL  FILL_4__2532_
timestamp 1701859473
transform -1 0 9830 0 1 2870
box -12 -8 32 272
use FILL  FILL_4__2533_
timestamp 1701859473
transform -1 0 8910 0 1 4430
box -12 -8 32 272
use FILL  FILL_4__2534_
timestamp 1701859473
transform -1 0 9310 0 -1 5470
box -12 -8 32 272
use FILL  FILL_4__2535_
timestamp 1701859473
transform 1 0 90 0 -1 4950
box -12 -8 32 272
use FILL  FILL_4__2536_
timestamp 1701859473
transform 1 0 650 0 1 4950
box -12 -8 32 272
use FILL  FILL_4__2537_
timestamp 1701859473
transform 1 0 790 0 1 3390
box -12 -8 32 272
use FILL  FILL_4__2538_
timestamp 1701859473
transform -1 0 350 0 -1 3910
box -12 -8 32 272
use FILL  FILL_4__2539_
timestamp 1701859473
transform -1 0 110 0 1 4950
box -12 -8 32 272
use FILL  FILL_4__2540_
timestamp 1701859473
transform 1 0 3050 0 1 2350
box -12 -8 32 272
use FILL  FILL_4__2541_
timestamp 1701859473
transform -1 0 3310 0 1 2870
box -12 -8 32 272
use FILL  FILL_4__2542_
timestamp 1701859473
transform -1 0 2310 0 -1 6510
box -12 -8 32 272
use FILL  FILL_4__2543_
timestamp 1701859473
transform 1 0 870 0 1 4950
box -12 -8 32 272
use FILL  FILL_4__2544_
timestamp 1701859473
transform 1 0 1430 0 1 4430
box -12 -8 32 272
use FILL  FILL_4__2545_
timestamp 1701859473
transform 1 0 1290 0 -1 5470
box -12 -8 32 272
use FILL  FILL_4__2546_
timestamp 1701859473
transform -1 0 2030 0 -1 5470
box -12 -8 32 272
use FILL  FILL_4__2547_
timestamp 1701859473
transform 1 0 1970 0 -1 4430
box -12 -8 32 272
use FILL  FILL_4__2548_
timestamp 1701859473
transform 1 0 1090 0 1 4950
box -12 -8 32 272
use FILL  FILL_4__2549_
timestamp 1701859473
transform 1 0 1310 0 1 4950
box -12 -8 32 272
use FILL  FILL_4__2550_
timestamp 1701859473
transform -1 0 1790 0 -1 5470
box -12 -8 32 272
use FILL  FILL_4__2551_
timestamp 1701859473
transform 1 0 2570 0 -1 9630
box -12 -8 32 272
use FILL  FILL_4__2552_
timestamp 1701859473
transform 1 0 3410 0 -1 5470
box -12 -8 32 272
use FILL  FILL_4__2553_
timestamp 1701859473
transform -1 0 2790 0 -1 6510
box -12 -8 32 272
use FILL  FILL_4__2554_
timestamp 1701859473
transform -1 0 3250 0 1 6510
box -12 -8 32 272
use FILL  FILL_4__2555_
timestamp 1701859473
transform -1 0 3490 0 1 6510
box -12 -8 32 272
use FILL  FILL_4__2556_
timestamp 1701859473
transform -1 0 2810 0 1 6510
box -12 -8 32 272
use FILL  FILL_4__2557_
timestamp 1701859473
transform 1 0 2510 0 -1 6510
box -12 -8 32 272
use FILL  FILL_4__2558_
timestamp 1701859473
transform 1 0 3250 0 -1 7550
box -12 -8 32 272
use FILL  FILL_4__2559_
timestamp 1701859473
transform 1 0 3450 0 -1 7550
box -12 -8 32 272
use FILL  FILL_4__2560_
timestamp 1701859473
transform -1 0 3510 0 1 7030
box -12 -8 32 272
use FILL  FILL_4__2561_
timestamp 1701859473
transform -1 0 1530 0 1 4950
box -12 -8 32 272
use FILL  FILL_4__2562_
timestamp 1701859473
transform 1 0 3250 0 1 7030
box -12 -8 32 272
use FILL  FILL_4__2563_
timestamp 1701859473
transform 1 0 3810 0 1 5470
box -12 -8 32 272
use FILL  FILL_4__2564_
timestamp 1701859473
transform -1 0 3690 0 1 6510
box -12 -8 32 272
use FILL  FILL_4__2565_
timestamp 1701859473
transform 1 0 3750 0 1 7030
box -12 -8 32 272
use FILL  FILL_4__2566_
timestamp 1701859473
transform 1 0 3210 0 1 7550
box -12 -8 32 272
use FILL  FILL_4__2567_
timestamp 1701859473
transform 1 0 3170 0 -1 8070
box -12 -8 32 272
use FILL  FILL_4__2568_
timestamp 1701859473
transform -1 0 2990 0 -1 8590
box -12 -8 32 272
use FILL  FILL_4__2569_
timestamp 1701859473
transform 1 0 2750 0 -1 8590
box -12 -8 32 272
use FILL  FILL_4__2570_
timestamp 1701859473
transform 1 0 2930 0 -1 8070
box -12 -8 32 272
use FILL  FILL_4__2571_
timestamp 1701859473
transform -1 0 3890 0 -1 9630
box -12 -8 32 272
use FILL  FILL_4__2572_
timestamp 1701859473
transform -1 0 3910 0 -1 5990
box -12 -8 32 272
use FILL  FILL_4__2573_
timestamp 1701859473
transform -1 0 3770 0 -1 7030
box -12 -8 32 272
use FILL  FILL_4__2574_
timestamp 1701859473
transform 1 0 3490 0 -1 6510
box -12 -8 32 272
use FILL  FILL_4__2575_
timestamp 1701859473
transform 1 0 3390 0 -1 8070
box -12 -8 32 272
use FILL  FILL_4__2576_
timestamp 1701859473
transform -1 0 3430 0 -1 8590
box -12 -8 32 272
use FILL  FILL_4__2577_
timestamp 1701859473
transform 1 0 3310 0 1 9110
box -12 -8 32 272
use FILL  FILL_4__2578_
timestamp 1701859473
transform 1 0 3810 0 1 9110
box -12 -8 32 272
use FILL  FILL_4__2579_
timestamp 1701859473
transform -1 0 2790 0 -1 9630
box -12 -8 32 272
use FILL  FILL_4__2580_
timestamp 1701859473
transform -1 0 4150 0 -1 9110
box -12 -8 32 272
use FILL  FILL_4__2581_
timestamp 1701859473
transform -1 0 4070 0 1 9110
box -12 -8 32 272
use FILL  FILL_4__2582_
timestamp 1701859473
transform 1 0 3570 0 1 9110
box -12 -8 32 272
use FILL  FILL_4__2583_
timestamp 1701859473
transform 1 0 3070 0 1 9110
box -12 -8 32 272
use FILL  FILL_4__2584_
timestamp 1701859473
transform 1 0 2830 0 1 9110
box -12 -8 32 272
use FILL  FILL_4__2585_
timestamp 1701859473
transform 1 0 3930 0 -1 9110
box -12 -8 32 272
use FILL  FILL_4__2586_
timestamp 1701859473
transform 1 0 3090 0 1 9630
box -12 -8 32 272
use FILL  FILL_4__2587_
timestamp 1701859473
transform 1 0 3670 0 -1 9110
box -12 -8 32 272
use FILL  FILL_4__2588_
timestamp 1701859473
transform 1 0 3270 0 1 8590
box -12 -8 32 272
use FILL  FILL_4__2589_
timestamp 1701859473
transform 1 0 3110 0 -1 10150
box -12 -8 32 272
use FILL  FILL_4__2590_
timestamp 1701859473
transform 1 0 2850 0 -1 10150
box -12 -8 32 272
use FILL  FILL_4__2591_
timestamp 1701859473
transform -1 0 3610 0 -1 11190
box -12 -8 32 272
use FILL  FILL_4__2592_
timestamp 1701859473
transform -1 0 3670 0 -1 9630
box -12 -8 32 272
use FILL  FILL_4__2593_
timestamp 1701859473
transform -1 0 3190 0 -1 9630
box -12 -8 32 272
use FILL  FILL_4__2594_
timestamp 1701859473
transform -1 0 3350 0 -1 10150
box -12 -8 32 272
use FILL  FILL_4__2595_
timestamp 1701859473
transform 1 0 3070 0 -1 11190
box -12 -8 32 272
use FILL  FILL_4__2596_
timestamp 1701859473
transform 1 0 3350 0 -1 11190
box -12 -8 32 272
use FILL  FILL_4__2597_
timestamp 1701859473
transform 1 0 2810 0 -1 10670
box -12 -8 32 272
use FILL  FILL_4__2598_
timestamp 1701859473
transform -1 0 3550 0 1 9630
box -12 -8 32 272
use FILL  FILL_4__2599_
timestamp 1701859473
transform -1 0 3330 0 1 9630
box -12 -8 32 272
use FILL  FILL_4__2600_
timestamp 1701859473
transform -1 0 3050 0 1 10150
box -12 -8 32 272
use FILL  FILL_4__2601_
timestamp 1701859473
transform 1 0 3010 0 -1 10670
box -12 -8 32 272
use FILL  FILL_4__2602_
timestamp 1701859473
transform -1 0 3270 0 -1 10670
box -12 -8 32 272
use FILL  FILL_4__2603_
timestamp 1701859473
transform 1 0 3470 0 -1 10670
box -12 -8 32 272
use FILL  FILL_4__2604_
timestamp 1701859473
transform 1 0 3270 0 1 10150
box -12 -8 32 272
use FILL  FILL_4__2605_
timestamp 1701859473
transform 1 0 2390 0 1 10670
box -12 -8 32 272
use FILL  FILL_4__2606_
timestamp 1701859473
transform 1 0 2590 0 1 10670
box -12 -8 32 272
use FILL  FILL_4__2607_
timestamp 1701859473
transform -1 0 2830 0 1 10670
box -12 -8 32 272
use FILL  FILL_4__2608_
timestamp 1701859473
transform -1 0 3790 0 1 9630
box -12 -8 32 272
use FILL  FILL_4__2609_
timestamp 1701859473
transform -1 0 2410 0 1 9630
box -12 -8 32 272
use FILL  FILL_4__2610_
timestamp 1701859473
transform -1 0 2630 0 -1 10150
box -12 -8 32 272
use FILL  FILL_4__2611_
timestamp 1701859473
transform -1 0 2350 0 -1 10670
box -12 -8 32 272
use FILL  FILL_4__2612_
timestamp 1701859473
transform 1 0 2570 0 -1 10670
box -12 -8 32 272
use FILL  FILL_4__2613_
timestamp 1701859473
transform 1 0 1890 0 1 10670
box -12 -8 32 272
use FILL  FILL_4__2614_
timestamp 1701859473
transform 1 0 1890 0 -1 10670
box -12 -8 32 272
use FILL  FILL_4__2615_
timestamp 1701859473
transform -1 0 2410 0 -1 11190
box -12 -8 32 272
use FILL  FILL_4__2616_
timestamp 1701859473
transform -1 0 3430 0 -1 9630
box -12 -8 32 272
use FILL  FILL_4__2617_
timestamp 1701859473
transform 1 0 2330 0 -1 9630
box -12 -8 32 272
use FILL  FILL_4__2618_
timestamp 1701859473
transform -1 0 2610 0 1 10150
box -12 -8 32 272
use FILL  FILL_4__2619_
timestamp 1701859473
transform 1 0 2110 0 1 10670
box -12 -8 32 272
use FILL  FILL_4__2620_
timestamp 1701859473
transform 1 0 2150 0 -1 11190
box -12 -8 32 272
use FILL  FILL_4__2621_
timestamp 1701859473
transform -1 0 1430 0 1 5470
box -12 -8 32 272
use FILL  FILL_4__2622_
timestamp 1701859473
transform -1 0 1270 0 -1 5990
box -12 -8 32 272
use FILL  FILL_4__2623_
timestamp 1701859473
transform 1 0 2490 0 -1 5470
box -12 -8 32 272
use FILL  FILL_4__2624_
timestamp 1701859473
transform -1 0 2450 0 1 5470
box -12 -8 32 272
use FILL  FILL_4__2625_
timestamp 1701859473
transform 1 0 2250 0 -1 5470
box -12 -8 32 272
use FILL  FILL_4__2626_
timestamp 1701859473
transform -1 0 990 0 -1 5470
box -12 -8 32 272
use FILL  FILL_4__2627_
timestamp 1701859473
transform -1 0 1510 0 1 3910
box -12 -8 32 272
use FILL  FILL_4__2628_
timestamp 1701859473
transform 1 0 1190 0 1 3910
box -12 -8 32 272
use FILL  FILL_4__2629_
timestamp 1701859473
transform -1 0 790 0 -1 5470
box -12 -8 32 272
use FILL  FILL_4__2630_
timestamp 1701859473
transform 1 0 770 0 -1 5990
box -12 -8 32 272
use FILL  FILL_4__2631_
timestamp 1701859473
transform -1 0 770 0 1 5990
box -12 -8 32 272
use FILL  FILL_4__2632_
timestamp 1701859473
transform 1 0 2150 0 1 10150
box -12 -8 32 272
use FILL  FILL_4__2633_
timestamp 1701859473
transform -1 0 2390 0 1 10150
box -12 -8 32 272
use FILL  FILL_4__2634_
timestamp 1701859473
transform 1 0 2350 0 -1 10150
box -12 -8 32 272
use FILL  FILL_4__2635_
timestamp 1701859473
transform 1 0 2130 0 -1 10150
box -12 -8 32 272
use FILL  FILL_4__2636_
timestamp 1701859473
transform -1 0 770 0 -1 10150
box -12 -8 32 272
use FILL  FILL_4__2637_
timestamp 1701859473
transform -1 0 570 0 1 6510
box -12 -8 32 272
use FILL  FILL_4__2638_
timestamp 1701859473
transform -1 0 350 0 1 6510
box -12 -8 32 272
use FILL  FILL_4__2639_
timestamp 1701859473
transform -1 0 330 0 -1 6510
box -12 -8 32 272
use FILL  FILL_4__2640_
timestamp 1701859473
transform -1 0 330 0 1 5990
box -12 -8 32 272
use FILL  FILL_4__2641_
timestamp 1701859473
transform 1 0 90 0 -1 7550
box -12 -8 32 272
use FILL  FILL_4__2642_
timestamp 1701859473
transform -1 0 430 0 1 4950
box -12 -8 32 272
use FILL  FILL_4__2643_
timestamp 1701859473
transform -1 0 2570 0 1 6510
box -12 -8 32 272
use FILL  FILL_4__2644_
timestamp 1701859473
transform 1 0 2610 0 -1 7030
box -12 -8 32 272
use FILL  FILL_4__2645_
timestamp 1701859473
transform 1 0 2790 0 1 7030
box -12 -8 32 272
use FILL  FILL_4__2646_
timestamp 1701859473
transform 1 0 2090 0 1 7030
box -12 -8 32 272
use FILL  FILL_4__2647_
timestamp 1701859473
transform 1 0 770 0 1 7550
box -12 -8 32 272
use FILL  FILL_4__2648_
timestamp 1701859473
transform 1 0 310 0 1 7550
box -12 -8 32 272
use FILL  FILL_4__2649_
timestamp 1701859473
transform 1 0 290 0 -1 7550
box -12 -8 32 272
use FILL  FILL_4__2650_
timestamp 1701859473
transform -1 0 770 0 -1 7550
box -12 -8 32 272
use FILL  FILL_4__2651_
timestamp 1701859473
transform 1 0 510 0 -1 7550
box -12 -8 32 272
use FILL  FILL_4__2652_
timestamp 1701859473
transform 1 0 510 0 1 7030
box -12 -8 32 272
use FILL  FILL_4__2653_
timestamp 1701859473
transform 1 0 90 0 1 7550
box -12 -8 32 272
use FILL  FILL_4__2654_
timestamp 1701859473
transform -1 0 570 0 1 7550
box -12 -8 32 272
use FILL  FILL_4__2655_
timestamp 1701859473
transform 1 0 1890 0 1 7030
box -12 -8 32 272
use FILL  FILL_4__2656_
timestamp 1701859473
transform 1 0 1530 0 -1 5470
box -12 -8 32 272
use FILL  FILL_4__2657_
timestamp 1701859473
transform -1 0 1730 0 1 5990
box -12 -8 32 272
use FILL  FILL_4__2658_
timestamp 1701859473
transform -1 0 2210 0 1 5470
box -12 -8 32 272
use FILL  FILL_4__2659_
timestamp 1701859473
transform 1 0 1970 0 -1 5990
box -12 -8 32 272
use FILL  FILL_4__2660_
timestamp 1701859473
transform -1 0 1970 0 1 5470
box -12 -8 32 272
use FILL  FILL_4__2661_
timestamp 1701859473
transform -1 0 1650 0 1 5470
box -12 -8 32 272
use FILL  FILL_4__2662_
timestamp 1701859473
transform 1 0 750 0 1 5470
box -12 -8 32 272
use FILL  FILL_4__2663_
timestamp 1701859473
transform -1 0 1030 0 -1 5990
box -12 -8 32 272
use FILL  FILL_4__2664_
timestamp 1701859473
transform 1 0 750 0 -1 7030
box -12 -8 32 272
use FILL  FILL_4__2665_
timestamp 1701859473
transform 1 0 1210 0 -1 7030
box -12 -8 32 272
use FILL  FILL_4__2666_
timestamp 1701859473
transform 1 0 1410 0 1 7030
box -12 -8 32 272
use FILL  FILL_4__2667_
timestamp 1701859473
transform 1 0 950 0 -1 7030
box -12 -8 32 272
use FILL  FILL_4__2668_
timestamp 1701859473
transform -1 0 2750 0 1 7550
box -12 -8 32 272
use FILL  FILL_4__2669_
timestamp 1701859473
transform 1 0 2690 0 -1 8070
box -12 -8 32 272
use FILL  FILL_4__2670_
timestamp 1701859473
transform 1 0 1950 0 -1 8070
box -12 -8 32 272
use FILL  FILL_4__2671_
timestamp 1701859473
transform -1 0 1450 0 1 7550
box -12 -8 32 272
use FILL  FILL_4__2672_
timestamp 1701859473
transform 1 0 1170 0 -1 7550
box -12 -8 32 272
use FILL  FILL_4__2673_
timestamp 1701859473
transform -1 0 1370 0 -1 7550
box -12 -8 32 272
use FILL  FILL_4__2674_
timestamp 1701859473
transform 1 0 1650 0 1 7030
box -12 -8 32 272
use FILL  FILL_4__2675_
timestamp 1701859473
transform 1 0 1590 0 -1 7550
box -12 -8 32 272
use FILL  FILL_4__2676_
timestamp 1701859473
transform -1 0 2030 0 -1 7550
box -12 -8 32 272
use FILL  FILL_4__2677_
timestamp 1701859473
transform 1 0 2430 0 -1 8070
box -12 -8 32 272
use FILL  FILL_4__2678_
timestamp 1701859473
transform -1 0 2210 0 -1 8070
box -12 -8 32 272
use FILL  FILL_4__2679_
timestamp 1701859473
transform -1 0 1650 0 1 8070
box -12 -8 32 272
use FILL  FILL_4__2680_
timestamp 1701859473
transform -1 0 330 0 -1 8590
box -12 -8 32 272
use FILL  FILL_4__2681_
timestamp 1701859473
transform 1 0 950 0 -1 7550
box -12 -8 32 272
use FILL  FILL_4__2682_
timestamp 1701859473
transform -1 0 330 0 -1 8070
box -12 -8 32 272
use FILL  FILL_4__2683_
timestamp 1701859473
transform -1 0 110 0 -1 9630
box -12 -8 32 272
use FILL  FILL_4__2684_
timestamp 1701859473
transform -1 0 110 0 1 10150
box -12 -8 32 272
use FILL  FILL_4__2685_
timestamp 1701859473
transform 1 0 990 0 1 5990
box -12 -8 32 272
use FILL  FILL_4__2686_
timestamp 1701859473
transform 1 0 970 0 1 7550
box -12 -8 32 272
use FILL  FILL_4__2687_
timestamp 1701859473
transform -1 0 970 0 -1 10150
box -12 -8 32 272
use FILL  FILL_4__2688_
timestamp 1701859473
transform 1 0 90 0 -1 10150
box -12 -8 32 272
use FILL  FILL_4__2689_
timestamp 1701859473
transform 1 0 310 0 -1 9630
box -12 -8 32 272
use FILL  FILL_4__2690_
timestamp 1701859473
transform 1 0 310 0 1 9110
box -12 -8 32 272
use FILL  FILL_4__2691_
timestamp 1701859473
transform 1 0 2770 0 1 8590
box -12 -8 32 272
use FILL  FILL_4__2692_
timestamp 1701859473
transform 1 0 2530 0 1 8590
box -12 -8 32 272
use FILL  FILL_4__2693_
timestamp 1701859473
transform -1 0 1190 0 -1 9630
box -12 -8 32 272
use FILL  FILL_4__2694_
timestamp 1701859473
transform 1 0 770 0 -1 9630
box -12 -8 32 272
use FILL  FILL_4__2695_
timestamp 1701859473
transform 1 0 90 0 1 9630
box -12 -8 32 272
use FILL  FILL_4__2696_
timestamp 1701859473
transform -1 0 570 0 -1 10150
box -12 -8 32 272
use FILL  FILL_4__2697_
timestamp 1701859473
transform 1 0 310 0 -1 10150
box -12 -8 32 272
use FILL  FILL_4__2698_
timestamp 1701859473
transform 1 0 330 0 1 9630
box -12 -8 32 272
use FILL  FILL_4__2699_
timestamp 1701859473
transform 1 0 550 0 -1 9630
box -12 -8 32 272
use FILL  FILL_4__2700_
timestamp 1701859473
transform 1 0 570 0 1 9630
box -12 -8 32 272
use FILL  FILL_4__2701_
timestamp 1701859473
transform -1 0 790 0 -1 10670
box -12 -8 32 272
use FILL  FILL_4__2702_
timestamp 1701859473
transform 1 0 3510 0 1 8590
box -12 -8 32 272
use FILL  FILL_4__2703_
timestamp 1701859473
transform -1 0 3050 0 1 8590
box -12 -8 32 272
use FILL  FILL_4__2704_
timestamp 1701859473
transform -1 0 1530 0 1 9630
box -12 -8 32 272
use FILL  FILL_4__2705_
timestamp 1701859473
transform 1 0 1270 0 1 9630
box -12 -8 32 272
use FILL  FILL_4__2706_
timestamp 1701859473
transform 1 0 290 0 1 10150
box -12 -8 32 272
use FILL  FILL_4__2707_
timestamp 1701859473
transform -1 0 530 0 1 10150
box -12 -8 32 272
use FILL  FILL_4__2708_
timestamp 1701859473
transform 1 0 730 0 1 10150
box -12 -8 32 272
use FILL  FILL_4__2709_
timestamp 1701859473
transform -1 0 550 0 -1 10670
box -12 -8 32 272
use FILL  FILL_4__2710_
timestamp 1701859473
transform 1 0 1730 0 1 10150
box -12 -8 32 272
use FILL  FILL_4__2711_
timestamp 1701859473
transform 1 0 2270 0 1 8590
box -12 -8 32 272
use FILL  FILL_4__2712_
timestamp 1701859473
transform -1 0 2050 0 1 8590
box -12 -8 32 272
use FILL  FILL_4__2713_
timestamp 1701859473
transform -1 0 1910 0 -1 9630
box -12 -8 32 272
use FILL  FILL_4__2714_
timestamp 1701859473
transform 1 0 1670 0 -1 10150
box -12 -8 32 272
use FILL  FILL_4__2715_
timestamp 1701859473
transform 1 0 990 0 1 10150
box -12 -8 32 272
use FILL  FILL_4__2716_
timestamp 1701859473
transform 1 0 1230 0 1 10150
box -12 -8 32 272
use FILL  FILL_4__2717_
timestamp 1701859473
transform 1 0 1490 0 1 10150
box -12 -8 32 272
use FILL  FILL_4__2718_
timestamp 1701859473
transform -1 0 10070 0 1 4950
box -12 -8 32 272
use FILL  FILL_4__2719_
timestamp 1701859473
transform -1 0 9830 0 1 4950
box -12 -8 32 272
use FILL  FILL_4__2720_
timestamp 1701859473
transform -1 0 4610 0 1 4950
box -12 -8 32 272
use FILL  FILL_4__2721_
timestamp 1701859473
transform -1 0 7370 0 -1 2350
box -12 -8 32 272
use FILL  FILL_4__2722_
timestamp 1701859473
transform 1 0 10010 0 -1 790
box -12 -8 32 272
use FILL  FILL_4__2723_
timestamp 1701859473
transform -1 0 7130 0 1 1830
box -12 -8 32 272
use FILL  FILL_4__2724_
timestamp 1701859473
transform -1 0 7130 0 -1 2350
box -12 -8 32 272
use FILL  FILL_4__2725_
timestamp 1701859473
transform 1 0 6990 0 1 3390
box -12 -8 32 272
use FILL  FILL_4__2726_
timestamp 1701859473
transform -1 0 7230 0 1 3390
box -12 -8 32 272
use FILL  FILL_4__2727_
timestamp 1701859473
transform -1 0 5450 0 1 3390
box -12 -8 32 272
use FILL  FILL_4__2728_
timestamp 1701859473
transform -1 0 5670 0 1 3390
box -12 -8 32 272
use FILL  FILL_4__2729_
timestamp 1701859473
transform -1 0 6770 0 -1 3910
box -12 -8 32 272
use FILL  FILL_4__2730_
timestamp 1701859473
transform 1 0 8270 0 -1 3910
box -12 -8 32 272
use FILL  FILL_4__2731_
timestamp 1701859473
transform 1 0 9290 0 1 1830
box -12 -8 32 272
use FILL  FILL_4__2732_
timestamp 1701859473
transform 1 0 7730 0 1 1830
box -12 -8 32 272
use FILL  FILL_4__2733_
timestamp 1701859473
transform 1 0 8610 0 1 2350
box -12 -8 32 272
use FILL  FILL_4__2734_
timestamp 1701859473
transform 1 0 7190 0 -1 5470
box -12 -8 32 272
use FILL  FILL_4__2735_
timestamp 1701859473
transform 1 0 7270 0 -1 2870
box -12 -8 32 272
use FILL  FILL_4__2736_
timestamp 1701859473
transform -1 0 7550 0 1 1310
box -12 -8 32 272
use FILL  FILL_4__2737_
timestamp 1701859473
transform 1 0 8610 0 1 1830
box -12 -8 32 272
use FILL  FILL_4__2738_
timestamp 1701859473
transform -1 0 7990 0 -1 2870
box -12 -8 32 272
use FILL  FILL_4__2739_
timestamp 1701859473
transform -1 0 7810 0 1 2870
box -12 -8 32 272
use FILL  FILL_4__2740_
timestamp 1701859473
transform -1 0 6590 0 -1 1830
box -12 -8 32 272
use FILL  FILL_4__2741_
timestamp 1701859473
transform 1 0 6790 0 -1 1830
box -12 -8 32 272
use FILL  FILL_4__2742_
timestamp 1701859473
transform -1 0 8230 0 -1 2870
box -12 -8 32 272
use FILL  FILL_4__2743_
timestamp 1701859473
transform -1 0 8250 0 1 2870
box -12 -8 32 272
use FILL  FILL_4__2744_
timestamp 1701859473
transform -1 0 7370 0 -1 270
box -12 -8 32 272
use FILL  FILL_4__2745_
timestamp 1701859473
transform -1 0 7330 0 1 1830
box -12 -8 32 272
use FILL  FILL_4__2746_
timestamp 1701859473
transform 1 0 7990 0 1 2870
box -12 -8 32 272
use FILL  FILL_4__2747_
timestamp 1701859473
transform -1 0 7790 0 -1 2350
box -12 -8 32 272
use FILL  FILL_4__2748_
timestamp 1701859473
transform 1 0 7970 0 -1 2350
box -12 -8 32 272
use FILL  FILL_4__2749_
timestamp 1701859473
transform 1 0 5930 0 1 1830
box -12 -8 32 272
use FILL  FILL_4__2750_
timestamp 1701859473
transform -1 0 6690 0 -1 1310
box -12 -8 32 272
use FILL  FILL_4__2751_
timestamp 1701859473
transform -1 0 6410 0 1 1830
box -12 -8 32 272
use FILL  FILL_4__2752_
timestamp 1701859473
transform -1 0 7770 0 1 2350
box -12 -8 32 272
use FILL  FILL_4__2753_
timestamp 1701859473
transform -1 0 7510 0 1 2350
box -12 -8 32 272
use FILL  FILL_4__2754_
timestamp 1701859473
transform 1 0 8850 0 -1 4950
box -12 -8 32 272
use FILL  FILL_4__2755_
timestamp 1701859473
transform 1 0 9750 0 1 790
box -12 -8 32 272
use FILL  FILL_4__2756_
timestamp 1701859473
transform -1 0 9990 0 1 790
box -12 -8 32 272
use FILL  FILL_4__2757_
timestamp 1701859473
transform 1 0 10690 0 -1 2870
box -12 -8 32 272
use FILL  FILL_4__2758_
timestamp 1701859473
transform -1 0 9190 0 -1 2870
box -12 -8 32 272
use FILL  FILL_4__2759_
timestamp 1701859473
transform 1 0 9110 0 1 4430
box -12 -8 32 272
use FILL  FILL_4__2760_
timestamp 1701859473
transform 1 0 10450 0 -1 790
box -12 -8 32 272
use FILL  FILL_4__2761_
timestamp 1701859473
transform 1 0 10210 0 -1 790
box -12 -8 32 272
use FILL  FILL_4__2762_
timestamp 1701859473
transform -1 0 10890 0 -1 1830
box -12 -8 32 272
use FILL  FILL_4__2763_
timestamp 1701859473
transform 1 0 6630 0 1 1830
box -12 -8 32 272
use FILL  FILL_4__2764_
timestamp 1701859473
transform -1 0 6890 0 1 1830
box -12 -8 32 272
use FILL  FILL_4__2765_
timestamp 1701859473
transform -1 0 10190 0 1 1830
box -12 -8 32 272
use FILL  FILL_4__2766_
timestamp 1701859473
transform -1 0 10010 0 -1 1830
box -12 -8 32 272
use FILL  FILL_4__2767_
timestamp 1701859473
transform -1 0 10430 0 -1 1830
box -12 -8 32 272
use FILL  FILL_4__2768_
timestamp 1701859473
transform -1 0 10410 0 1 1830
box -12 -8 32 272
use FILL  FILL_4__2769_
timestamp 1701859473
transform -1 0 10870 0 1 2350
box -12 -8 32 272
use FILL  FILL_4__2770_
timestamp 1701859473
transform -1 0 10650 0 -1 1830
box -12 -8 32 272
use FILL  FILL_4__2771_
timestamp 1701859473
transform 1 0 11070 0 1 2350
box -12 -8 32 272
use FILL  FILL_4__2772_
timestamp 1701859473
transform -1 0 10730 0 1 4950
box -12 -8 32 272
use FILL  FILL_4__2773_
timestamp 1701859473
transform 1 0 10470 0 -1 3910
box -12 -8 32 272
use FILL  FILL_4__2774_
timestamp 1701859473
transform -1 0 10770 0 -1 2350
box -12 -8 32 272
use FILL  FILL_4__2775_
timestamp 1701859473
transform -1 0 9130 0 -1 1310
box -12 -8 32 272
use FILL  FILL_4__2776_
timestamp 1701859473
transform 1 0 10670 0 -1 790
box -12 -8 32 272
use FILL  FILL_4__2777_
timestamp 1701859473
transform -1 0 8430 0 -1 270
box -12 -8 32 272
use FILL  FILL_4__2778_
timestamp 1701859473
transform 1 0 10970 0 1 270
box -12 -8 32 272
use FILL  FILL_4__2779_
timestamp 1701859473
transform 1 0 9050 0 -1 1830
box -12 -8 32 272
use FILL  FILL_4__2780_
timestamp 1701859473
transform -1 0 10070 0 1 1310
box -12 -8 32 272
use FILL  FILL_4__2781_
timestamp 1701859473
transform 1 0 10210 0 -1 1310
box -12 -8 32 272
use FILL  FILL_4__2782_
timestamp 1701859473
transform 1 0 8830 0 1 1830
box -12 -8 32 272
use FILL  FILL_4__2783_
timestamp 1701859473
transform 1 0 8390 0 -1 1310
box -12 -8 32 272
use FILL  FILL_4__2784_
timestamp 1701859473
transform 1 0 8630 0 -1 1310
box -12 -8 32 272
use FILL  FILL_4__2785_
timestamp 1701859473
transform 1 0 8850 0 -1 1830
box -12 -8 32 272
use FILL  FILL_4__2786_
timestamp 1701859473
transform -1 0 9330 0 -1 1310
box -12 -8 32 272
use FILL  FILL_4__2787_
timestamp 1701859473
transform -1 0 9530 0 -1 1830
box -12 -8 32 272
use FILL  FILL_4__2788_
timestamp 1701859473
transform 1 0 10210 0 -1 1830
box -12 -8 32 272
use FILL  FILL_4__2789_
timestamp 1701859473
transform 1 0 10290 0 1 1310
box -12 -8 32 272
use FILL  FILL_4__2790_
timestamp 1701859473
transform -1 0 10090 0 -1 2350
box -12 -8 32 272
use FILL  FILL_4__2791_
timestamp 1701859473
transform 1 0 9850 0 -1 2350
box -12 -8 32 272
use FILL  FILL_4__2792_
timestamp 1701859473
transform -1 0 10310 0 -1 2350
box -12 -8 32 272
use FILL  FILL_4__2793_
timestamp 1701859473
transform -1 0 10550 0 -1 2350
box -12 -8 32 272
use FILL  FILL_4__2794_
timestamp 1701859473
transform -1 0 10970 0 -1 2350
box -12 -8 32 272
use FILL  FILL_4__2795_
timestamp 1701859473
transform -1 0 10930 0 -1 2870
box -12 -8 32 272
use FILL  FILL_4__2796_
timestamp 1701859473
transform -1 0 10270 0 -1 2870
box -12 -8 32 272
use FILL  FILL_4__2797_
timestamp 1701859473
transform -1 0 9770 0 -1 1830
box -12 -8 32 272
use FILL  FILL_4__2798_
timestamp 1701859473
transform -1 0 10650 0 1 2350
box -12 -8 32 272
use FILL  FILL_4__2799_
timestamp 1701859473
transform 1 0 10430 0 -1 2870
box -12 -8 32 272
use FILL  FILL_4__2800_
timestamp 1701859473
transform -1 0 10450 0 -1 4430
box -12 -8 32 272
use FILL  FILL_4__2801_
timestamp 1701859473
transform -1 0 9410 0 -1 2870
box -12 -8 32 272
use FILL  FILL_4__2802_
timestamp 1701859473
transform -1 0 7270 0 -1 1830
box -12 -8 32 272
use FILL  FILL_4__2803_
timestamp 1701859473
transform 1 0 8470 0 -1 2870
box -12 -8 32 272
use FILL  FILL_4__2804_
timestamp 1701859473
transform -1 0 9530 0 -1 3390
box -12 -8 32 272
use FILL  FILL_4__2805_
timestamp 1701859473
transform -1 0 9830 0 -1 2870
box -12 -8 32 272
use FILL  FILL_4__2806_
timestamp 1701859473
transform 1 0 9590 0 -1 2870
box -12 -8 32 272
use FILL  FILL_4__2807_
timestamp 1701859473
transform 1 0 8930 0 -1 2350
box -12 -8 32 272
use FILL  FILL_4__2808_
timestamp 1701859473
transform 1 0 8690 0 -1 2350
box -12 -8 32 272
use FILL  FILL_4__2809_
timestamp 1701859473
transform 1 0 10410 0 1 2350
box -12 -8 32 272
use FILL  FILL_4__2810_
timestamp 1701859473
transform -1 0 10190 0 1 2350
box -12 -8 32 272
use FILL  FILL_4__2811_
timestamp 1701859473
transform 1 0 4970 0 -1 4430
box -12 -8 32 272
use FILL  FILL_4__2812_
timestamp 1701859473
transform -1 0 8930 0 1 4950
box -12 -8 32 272
use FILL  FILL_4__2813_
timestamp 1701859473
transform 1 0 9030 0 1 3390
box -12 -8 32 272
use FILL  FILL_4__2814_
timestamp 1701859473
transform -1 0 8850 0 -1 4430
box -12 -8 32 272
use FILL  FILL_4__2815_
timestamp 1701859473
transform -1 0 8630 0 1 3910
box -12 -8 32 272
use FILL  FILL_4__2816_
timestamp 1701859473
transform -1 0 8250 0 1 4950
box -12 -8 32 272
use FILL  FILL_4__2817_
timestamp 1701859473
transform 1 0 8690 0 1 4950
box -12 -8 32 272
use FILL  FILL_4__2818_
timestamp 1701859473
transform 1 0 8390 0 -1 4430
box -12 -8 32 272
use FILL  FILL_4__2819_
timestamp 1701859473
transform 1 0 8590 0 -1 4430
box -12 -8 32 272
use FILL  FILL_4__2820_
timestamp 1701859473
transform -1 0 9550 0 1 2350
box -12 -8 32 272
use FILL  FILL_4__2821_
timestamp 1701859473
transform 1 0 9070 0 1 2350
box -12 -8 32 272
use FILL  FILL_4__2822_
timestamp 1701859473
transform -1 0 9070 0 1 1830
box -12 -8 32 272
use FILL  FILL_4__2823_
timestamp 1701859473
transform -1 0 8850 0 1 2350
box -12 -8 32 272
use FILL  FILL_4__2824_
timestamp 1701859473
transform 1 0 9970 0 -1 3390
box -12 -8 32 272
use FILL  FILL_4__2825_
timestamp 1701859473
transform -1 0 10690 0 -1 3390
box -12 -8 32 272
use FILL  FILL_4__2826_
timestamp 1701859473
transform 1 0 9550 0 1 790
box -12 -8 32 272
use FILL  FILL_4__2827_
timestamp 1701859473
transform -1 0 9290 0 -1 1830
box -12 -8 32 272
use FILL  FILL_4__2828_
timestamp 1701859473
transform 1 0 7010 0 -1 1830
box -12 -8 32 272
use FILL  FILL_4__2829_
timestamp 1701859473
transform -1 0 10030 0 1 2870
box -12 -8 32 272
use FILL  FILL_4__2830_
timestamp 1701859473
transform 1 0 8330 0 -1 3390
box -12 -8 32 272
use FILL  FILL_4__2831_
timestamp 1701859473
transform 1 0 8370 0 1 3910
box -12 -8 32 272
use FILL  FILL_4__2832_
timestamp 1701859473
transform -1 0 9350 0 1 2350
box -12 -8 32 272
use FILL  FILL_4__2833_
timestamp 1701859473
transform -1 0 9290 0 -1 3390
box -12 -8 32 272
use FILL  FILL_4__2834_
timestamp 1701859473
transform -1 0 9050 0 -1 3390
box -12 -8 32 272
use FILL  FILL_4__2835_
timestamp 1701859473
transform -1 0 9350 0 1 790
box -12 -8 32 272
use FILL  FILL_4__2836_
timestamp 1701859473
transform 1 0 8930 0 1 1310
box -12 -8 32 272
use FILL  FILL_4__2837_
timestamp 1701859473
transform -1 0 9610 0 1 1310
box -12 -8 32 272
use FILL  FILL_4__2838_
timestamp 1701859473
transform -1 0 9730 0 1 3390
box -12 -8 32 272
use FILL  FILL_4__2839_
timestamp 1701859473
transform -1 0 9770 0 -1 3390
box -12 -8 32 272
use FILL  FILL_4__2840_
timestamp 1701859473
transform 1 0 9090 0 -1 270
box -12 -8 32 272
use FILL  FILL_4__2841_
timestamp 1701859473
transform -1 0 8890 0 -1 270
box -12 -8 32 272
use FILL  FILL_4__2842_
timestamp 1701859473
transform 1 0 9310 0 -1 270
box -12 -8 32 272
use FILL  FILL_4__2843_
timestamp 1701859473
transform 1 0 9550 0 -1 270
box -12 -8 32 272
use FILL  FILL_4__2844_
timestamp 1701859473
transform 1 0 9350 0 1 270
box -12 -8 32 272
use FILL  FILL_4__2845_
timestamp 1701859473
transform -1 0 10030 0 1 270
box -12 -8 32 272
use FILL  FILL_4__2846_
timestamp 1701859473
transform 1 0 9770 0 1 270
box -12 -8 32 272
use FILL  FILL_4__2847_
timestamp 1701859473
transform -1 0 11170 0 -1 10670
box -12 -8 32 272
use FILL  FILL_4__2848_
timestamp 1701859473
transform -1 0 10650 0 -1 1310
box -12 -8 32 272
use FILL  FILL_4__2849_
timestamp 1701859473
transform -1 0 10990 0 1 1310
box -12 -8 32 272
use FILL  FILL_4__2850_
timestamp 1701859473
transform -1 0 11130 0 -1 1830
box -12 -8 32 272
use FILL  FILL_4__2851_
timestamp 1701859473
transform 1 0 10730 0 -1 3910
box -12 -8 32 272
use FILL  FILL_4__2852_
timestamp 1701859473
transform -1 0 8930 0 1 270
box -12 -8 32 272
use FILL  FILL_4__2853_
timestamp 1701859473
transform -1 0 9150 0 1 270
box -12 -8 32 272
use FILL  FILL_4__2854_
timestamp 1701859473
transform 1 0 10650 0 1 790
box -12 -8 32 272
use FILL  FILL_4__2855_
timestamp 1701859473
transform -1 0 9850 0 1 1310
box -12 -8 32 272
use FILL  FILL_4__2856_
timestamp 1701859473
transform -1 0 10510 0 1 1310
box -12 -8 32 272
use FILL  FILL_4__2857_
timestamp 1701859473
transform -1 0 10750 0 1 1310
box -12 -8 32 272
use FILL  FILL_4__2858_
timestamp 1701859473
transform -1 0 11110 0 1 1830
box -12 -8 32 272
use FILL  FILL_4__2859_
timestamp 1701859473
transform 1 0 10970 0 -1 3910
box -12 -8 32 272
use FILL  FILL_4__2860_
timestamp 1701859473
transform 1 0 10890 0 -1 3390
box -12 -8 32 272
use FILL  FILL_4__2861_
timestamp 1701859473
transform 1 0 9770 0 -1 270
box -12 -8 32 272
use FILL  FILL_4__2862_
timestamp 1701859473
transform 1 0 8630 0 -1 270
box -12 -8 32 272
use FILL  FILL_4__2863_
timestamp 1701859473
transform -1 0 10270 0 1 270
box -12 -8 32 272
use FILL  FILL_4__2864_
timestamp 1701859473
transform 1 0 10510 0 1 270
box -12 -8 32 272
use FILL  FILL_4__2865_
timestamp 1701859473
transform -1 0 10750 0 1 270
box -12 -8 32 272
use FILL  FILL_4__2866_
timestamp 1701859473
transform -1 0 11130 0 -1 790
box -12 -8 32 272
use FILL  FILL_4__2867_
timestamp 1701859473
transform 1 0 11090 0 -1 3390
box -12 -8 32 272
use FILL  FILL_4__2868_
timestamp 1701859473
transform 1 0 11070 0 1 790
box -12 -8 32 272
use FILL  FILL_4__2869_
timestamp 1701859473
transform 1 0 10190 0 1 790
box -12 -8 32 272
use FILL  FILL_4__2870_
timestamp 1701859473
transform -1 0 10410 0 1 790
box -12 -8 32 272
use FILL  FILL_4__2871_
timestamp 1701859473
transform -1 0 10850 0 1 790
box -12 -8 32 272
use FILL  FILL_4__2872_
timestamp 1701859473
transform -1 0 11190 0 1 1310
box -12 -8 32 272
use FILL  FILL_4__2873_
timestamp 1701859473
transform -1 0 9970 0 1 3390
box -12 -8 32 272
use FILL  FILL_4__2874_
timestamp 1701859473
transform -1 0 10210 0 1 3390
box -12 -8 32 272
use FILL  FILL_4__2875_
timestamp 1701859473
transform -1 0 10790 0 -1 4950
box -12 -8 32 272
use FILL  FILL_4__2876_
timestamp 1701859473
transform -1 0 9750 0 1 1830
box -12 -8 32 272
use FILL  FILL_4__2877_
timestamp 1701859473
transform 1 0 9930 0 1 1830
box -12 -8 32 272
use FILL  FILL_4__2878_
timestamp 1701859473
transform 1 0 9750 0 -1 1310
box -12 -8 32 272
use FILL  FILL_4__2879_
timestamp 1701859473
transform -1 0 9990 0 -1 1310
box -12 -8 32 272
use FILL  FILL_4__2880_
timestamp 1701859473
transform 1 0 9490 0 1 1830
box -12 -8 32 272
use FILL  FILL_4__2881_
timestamp 1701859473
transform 1 0 10870 0 -1 790
box -12 -8 32 272
use FILL  FILL_4__2882_
timestamp 1701859473
transform -1 0 9550 0 -1 1310
box -12 -8 32 272
use FILL  FILL_4__2883_
timestamp 1701859473
transform -1 0 10450 0 -1 1310
box -12 -8 32 272
use FILL  FILL_4__2884_
timestamp 1701859473
transform 1 0 11090 0 -1 1310
box -12 -8 32 272
use FILL  FILL_4__2885_
timestamp 1701859473
transform -1 0 10870 0 -1 1310
box -12 -8 32 272
use FILL  FILL_4__2886_
timestamp 1701859473
transform 1 0 10630 0 1 1830
box -12 -8 32 272
use FILL  FILL_4__2887_
timestamp 1701859473
transform 1 0 10190 0 -1 4430
box -12 -8 32 272
use FILL  FILL_4__2888_
timestamp 1701859473
transform -1 0 4010 0 1 5470
box -12 -8 32 272
use FILL  FILL_4__2889_
timestamp 1701859473
transform 1 0 6130 0 1 2350
box -12 -8 32 272
use FILL  FILL_4__2890_
timestamp 1701859473
transform -1 0 8410 0 1 5990
box -12 -8 32 272
use FILL  FILL_4__2891_
timestamp 1701859473
transform -1 0 8210 0 1 5990
box -12 -8 32 272
use FILL  FILL_4__2892_
timestamp 1701859473
transform 1 0 7430 0 -1 5470
box -12 -8 32 272
use FILL  FILL_4__2893_
timestamp 1701859473
transform 1 0 7250 0 1 5470
box -12 -8 32 272
use FILL  FILL_4__2894_
timestamp 1701859473
transform 1 0 6530 0 -1 6510
box -12 -8 32 272
use FILL  FILL_4__2895_
timestamp 1701859473
transform 1 0 6670 0 1 6510
box -12 -8 32 272
use FILL  FILL_4__2896_
timestamp 1701859473
transform -1 0 7930 0 -1 5470
box -12 -8 32 272
use FILL  FILL_4__2897_
timestamp 1701859473
transform 1 0 7730 0 1 5470
box -12 -8 32 272
use FILL  FILL_4__2898_
timestamp 1701859473
transform 1 0 7250 0 -1 6510
box -12 -8 32 272
use FILL  FILL_4__2899_
timestamp 1701859473
transform 1 0 6770 0 -1 6510
box -12 -8 32 272
use FILL  FILL_4__2900_
timestamp 1701859473
transform -1 0 6310 0 -1 6510
box -12 -8 32 272
use FILL  FILL_4__2901_
timestamp 1701859473
transform 1 0 6050 0 -1 6510
box -12 -8 32 272
use FILL  FILL_4__2902_
timestamp 1701859473
transform -1 0 7970 0 1 5990
box -12 -8 32 272
use FILL  FILL_4__2903_
timestamp 1701859473
transform 1 0 7250 0 1 5990
box -12 -8 32 272
use FILL  FILL_4__2904_
timestamp 1701859473
transform 1 0 8370 0 -1 5470
box -12 -8 32 272
use FILL  FILL_4__2905_
timestamp 1701859473
transform 1 0 8390 0 1 5470
box -12 -8 32 272
use FILL  FILL_4__2906_
timestamp 1701859473
transform 1 0 8130 0 -1 5990
box -12 -8 32 272
use FILL  FILL_4__2907_
timestamp 1701859473
transform -1 0 7910 0 -1 5990
box -12 -8 32 272
use FILL  FILL_4__2908_
timestamp 1701859473
transform -1 0 8230 0 -1 4950
box -12 -8 32 272
use FILL  FILL_4__2909_
timestamp 1701859473
transform 1 0 3370 0 -1 4430
box -12 -8 32 272
use FILL  FILL_4__2910_
timestamp 1701859473
transform -1 0 6530 0 -1 4430
box -12 -8 32 272
use FILL  FILL_4__2911_
timestamp 1701859473
transform -1 0 6870 0 1 4430
box -12 -8 32 272
use FILL  FILL_4__2912_
timestamp 1701859473
transform 1 0 8650 0 -1 4950
box -12 -8 32 272
use FILL  FILL_4__2913_
timestamp 1701859473
transform -1 0 6830 0 -1 4950
box -12 -8 32 272
use FILL  FILL_4__2914_
timestamp 1701859473
transform 1 0 7090 0 -1 8070
box -12 -8 32 272
use FILL  FILL_4__2915_
timestamp 1701859473
transform 1 0 7210 0 -1 5990
box -12 -8 32 272
use FILL  FILL_4__2916_
timestamp 1701859473
transform 1 0 6970 0 -1 5990
box -12 -8 32 272
use FILL  FILL_4__2917_
timestamp 1701859473
transform -1 0 6350 0 -1 5990
box -12 -8 32 272
use FILL  FILL_4__2918_
timestamp 1701859473
transform 1 0 6270 0 1 5470
box -12 -8 32 272
use FILL  FILL_4__2919_
timestamp 1701859473
transform 1 0 6190 0 1 4950
box -12 -8 32 272
use FILL  FILL_4__2920_
timestamp 1701859473
transform 1 0 5950 0 1 4950
box -12 -8 32 272
use FILL  FILL_4__2921_
timestamp 1701859473
transform -1 0 7410 0 -1 3910
box -12 -8 32 272
use FILL  FILL_4__2922_
timestamp 1701859473
transform -1 0 7450 0 1 3910
box -12 -8 32 272
use FILL  FILL_4__2923_
timestamp 1701859473
transform -1 0 6770 0 -1 4430
box -12 -8 32 272
use FILL  FILL_4__2924_
timestamp 1701859473
transform 1 0 6390 0 1 4950
box -12 -8 32 272
use FILL  FILL_4__2925_
timestamp 1701859473
transform 1 0 7290 0 1 7550
box -12 -8 32 272
use FILL  FILL_4__2926_
timestamp 1701859473
transform -1 0 7530 0 1 4430
box -12 -8 32 272
use FILL  FILL_4__2927_
timestamp 1701859473
transform 1 0 7310 0 -1 4950
box -12 -8 32 272
use FILL  FILL_4__2928_
timestamp 1701859473
transform 1 0 7050 0 -1 4950
box -12 -8 32 272
use FILL  FILL_4__2929_
timestamp 1701859473
transform -1 0 6630 0 1 4950
box -12 -8 32 272
use FILL  FILL_4__2930_
timestamp 1701859473
transform 1 0 6170 0 1 1830
box -12 -8 32 272
use FILL  FILL_4__2931_
timestamp 1701859473
transform 1 0 7050 0 -1 2870
box -12 -8 32 272
use FILL  FILL_4__2932_
timestamp 1701859473
transform 1 0 5210 0 -1 4430
box -12 -8 32 272
use FILL  FILL_4__2933_
timestamp 1701859473
transform 1 0 5410 0 -1 4430
box -12 -8 32 272
use FILL  FILL_4__2934_
timestamp 1701859473
transform 1 0 5650 0 -1 4430
box -12 -8 32 272
use FILL  FILL_4__2935_
timestamp 1701859473
transform 1 0 6470 0 1 6510
box -12 -8 32 272
use FILL  FILL_4__2936_
timestamp 1701859473
transform 1 0 6350 0 -1 4950
box -12 -8 32 272
use FILL  FILL_4__2937_
timestamp 1701859473
transform 1 0 6570 0 -1 4950
box -12 -8 32 272
use FILL  FILL_4__2938_
timestamp 1701859473
transform 1 0 5050 0 1 4950
box -12 -8 32 272
use FILL  FILL_4__2939_
timestamp 1701859473
transform 1 0 4830 0 1 4950
box -12 -8 32 272
use FILL  FILL_4__2940_
timestamp 1701859473
transform -1 0 5890 0 -1 5470
box -12 -8 32 272
use FILL  FILL_4__2941_
timestamp 1701859473
transform 1 0 5650 0 -1 5470
box -12 -8 32 272
use FILL  FILL_4__2942_
timestamp 1701859473
transform -1 0 9350 0 1 4430
box -12 -8 32 272
use FILL  FILL_4__2943_
timestamp 1701859473
transform 1 0 6310 0 -1 4430
box -12 -8 32 272
use FILL  FILL_4__2944_
timestamp 1701859473
transform -1 0 6330 0 1 3910
box -12 -8 32 272
use FILL  FILL_4__2945_
timestamp 1701859473
transform -1 0 6410 0 1 4430
box -12 -8 32 272
use FILL  FILL_4__2946_
timestamp 1701859473
transform 1 0 6170 0 1 4430
box -12 -8 32 272
use FILL  FILL_4__2947_
timestamp 1701859473
transform -1 0 6570 0 -1 5990
box -12 -8 32 272
use FILL  FILL_4__2948_
timestamp 1701859473
transform 1 0 6110 0 -1 5990
box -12 -8 32 272
use FILL  FILL_4__2949_
timestamp 1701859473
transform -1 0 5930 0 -1 5990
box -12 -8 32 272
use FILL  FILL_4__2950_
timestamp 1701859473
transform 1 0 5790 0 1 5470
box -12 -8 32 272
use FILL  FILL_4__2951_
timestamp 1701859473
transform -1 0 6050 0 1 5470
box -12 -8 32 272
use FILL  FILL_4__2952_
timestamp 1701859473
transform -1 0 6130 0 -1 4950
box -12 -8 32 272
use FILL  FILL_4__2953_
timestamp 1701859473
transform -1 0 4410 0 1 4950
box -12 -8 32 272
use FILL  FILL_4__2954_
timestamp 1701859473
transform -1 0 6670 0 1 4430
box -12 -8 32 272
use FILL  FILL_4__2955_
timestamp 1701859473
transform -1 0 5950 0 1 4430
box -12 -8 32 272
use FILL  FILL_4__2956_
timestamp 1701859473
transform 1 0 5230 0 1 4430
box -12 -8 32 272
use FILL  FILL_4__2957_
timestamp 1701859473
transform 1 0 5170 0 -1 4950
box -12 -8 32 272
use FILL  FILL_4__2958_
timestamp 1701859473
transform -1 0 5490 0 1 4430
box -12 -8 32 272
use FILL  FILL_4__2959_
timestamp 1701859473
transform 1 0 6990 0 -1 5470
box -12 -8 32 272
use FILL  FILL_4__2960_
timestamp 1701859473
transform -1 0 6530 0 1 5470
box -12 -8 32 272
use FILL  FILL_4__2961_
timestamp 1701859473
transform 1 0 6290 0 -1 5470
box -12 -8 32 272
use FILL  FILL_4__2962_
timestamp 1701859473
transform -1 0 6550 0 -1 5470
box -12 -8 32 272
use FILL  FILL_4__2963_
timestamp 1701859473
transform -1 0 6790 0 -1 5470
box -12 -8 32 272
use FILL  FILL_4__2964_
timestamp 1701859473
transform -1 0 5430 0 -1 4950
box -12 -8 32 272
use FILL  FILL_4__2965_
timestamp 1701859473
transform 1 0 4930 0 -1 4950
box -12 -8 32 272
use FILL  FILL_4__2966_
timestamp 1701859473
transform -1 0 6390 0 1 2350
box -12 -8 32 272
use FILL  FILL_4__2967_
timestamp 1701859473
transform 1 0 7650 0 1 3910
box -12 -8 32 272
use FILL  FILL_4__2968_
timestamp 1701859473
transform -1 0 6970 0 -1 3910
box -12 -8 32 272
use FILL  FILL_4__2969_
timestamp 1701859473
transform -1 0 7190 0 -1 3910
box -12 -8 32 272
use FILL  FILL_4__2970_
timestamp 1701859473
transform -1 0 7230 0 1 3910
box -12 -8 32 272
use FILL  FILL_4__2971_
timestamp 1701859473
transform -1 0 6750 0 1 3910
box -12 -8 32 272
use FILL  FILL_4__2972_
timestamp 1701859473
transform 1 0 6970 0 1 3910
box -12 -8 32 272
use FILL  FILL_4__2973_
timestamp 1701859473
transform -1 0 7090 0 1 4430
box -12 -8 32 272
use FILL  FILL_4__2974_
timestamp 1701859473
transform 1 0 6990 0 -1 4430
box -12 -8 32 272
use FILL  FILL_4__2975_
timestamp 1701859473
transform -1 0 7750 0 -1 4430
box -12 -8 32 272
use FILL  FILL_4__2976_
timestamp 1701859473
transform -1 0 7510 0 -1 4430
box -12 -8 32 272
use FILL  FILL_4__2977_
timestamp 1701859473
transform 1 0 7230 0 -1 4430
box -12 -8 32 272
use FILL  FILL_4__2978_
timestamp 1701859473
transform 1 0 7290 0 1 4430
box -12 -8 32 272
use FILL  FILL_4__2979_
timestamp 1701859473
transform -1 0 3630 0 -1 4950
box -12 -8 32 272
use FILL  FILL_4__2980_
timestamp 1701859473
transform -1 0 3010 0 1 7550
box -12 -8 32 272
use FILL  FILL_4__2981_
timestamp 1701859473
transform 1 0 3530 0 1 4950
box -12 -8 32 272
use FILL  FILL_4__2982_
timestamp 1701859473
transform 1 0 9590 0 1 6510
box -12 -8 32 272
use FILL  FILL_4__2983_
timestamp 1701859473
transform 1 0 1910 0 1 4430
box -12 -8 32 272
use FILL  FILL_4__2984_
timestamp 1701859473
transform -1 0 3530 0 -1 3910
box -12 -8 32 272
use FILL  FILL_4__2985_
timestamp 1701859473
transform 1 0 3690 0 1 4430
box -12 -8 32 272
use FILL  FILL_4__2986_
timestamp 1701859473
transform -1 0 5890 0 -1 4430
box -12 -8 32 272
use FILL  FILL_4__2987_
timestamp 1701859473
transform -1 0 5710 0 1 4430
box -12 -8 32 272
use FILL  FILL_4__2988_
timestamp 1701859473
transform 1 0 9370 0 1 6510
box -12 -8 32 272
use FILL  FILL_4__2989_
timestamp 1701859473
transform 1 0 5990 0 1 6510
box -12 -8 32 272
use FILL  FILL_4__2990_
timestamp 1701859473
transform -1 0 6250 0 1 6510
box -12 -8 32 272
use FILL  FILL_4__2991_
timestamp 1701859473
transform 1 0 7150 0 1 6510
box -12 -8 32 272
use FILL  FILL_4__2992_
timestamp 1701859473
transform 1 0 9670 0 1 7030
box -12 -8 32 272
use FILL  FILL_4__2993_
timestamp 1701859473
transform 1 0 9870 0 1 7030
box -12 -8 32 272
use FILL  FILL_4__2994_
timestamp 1701859473
transform -1 0 10790 0 -1 7550
box -12 -8 32 272
use FILL  FILL_4__2995_
timestamp 1701859473
transform -1 0 7590 0 -1 7550
box -12 -8 32 272
use FILL  FILL_4__2996_
timestamp 1701859473
transform 1 0 7490 0 1 7550
box -12 -8 32 272
use FILL  FILL_4__2997_
timestamp 1701859473
transform -1 0 7370 0 -1 7550
box -12 -8 32 272
use FILL  FILL_4__2998_
timestamp 1701859473
transform -1 0 6430 0 -1 7550
box -12 -8 32 272
use FILL  FILL_4__2999_
timestamp 1701859473
transform 1 0 6150 0 1 7550
box -12 -8 32 272
use FILL  FILL_4__3000_
timestamp 1701859473
transform -1 0 5990 0 -1 7550
box -12 -8 32 272
use FILL  FILL_4__3001_
timestamp 1701859473
transform -1 0 5770 0 -1 7550
box -12 -8 32 272
use FILL  FILL_4__3002_
timestamp 1701859473
transform -1 0 6190 0 -1 7550
box -12 -8 32 272
use FILL  FILL_4__3003_
timestamp 1701859473
transform -1 0 6370 0 1 7550
box -12 -8 32 272
use FILL  FILL_4__3004_
timestamp 1701859473
transform 1 0 8170 0 1 7550
box -12 -8 32 272
use FILL  FILL_4__3005_
timestamp 1701859473
transform 1 0 10990 0 -1 7550
box -12 -8 32 272
use FILL  FILL_4__3006_
timestamp 1701859473
transform -1 0 10470 0 1 7550
box -12 -8 32 272
use FILL  FILL_4__3007_
timestamp 1701859473
transform 1 0 6990 0 1 7030
box -12 -8 32 272
use FILL  FILL_4__3008_
timestamp 1701859473
transform -1 0 6550 0 1 7030
box -12 -8 32 272
use FILL  FILL_4__3009_
timestamp 1701859473
transform -1 0 5950 0 -1 7030
box -12 -8 32 272
use FILL  FILL_4__3010_
timestamp 1701859473
transform 1 0 6170 0 -1 7030
box -12 -8 32 272
use FILL  FILL_4__3011_
timestamp 1701859473
transform 1 0 6750 0 1 7030
box -12 -8 32 272
use FILL  FILL_4__3012_
timestamp 1701859473
transform -1 0 7870 0 -1 7030
box -12 -8 32 272
use FILL  FILL_4__3013_
timestamp 1701859473
transform 1 0 8310 0 -1 7030
box -12 -8 32 272
use FILL  FILL_4__3014_
timestamp 1701859473
transform 1 0 10670 0 1 7550
box -12 -8 32 272
use FILL  FILL_4__3015_
timestamp 1701859473
transform -1 0 6390 0 -1 7030
box -12 -8 32 272
use FILL  FILL_4__3016_
timestamp 1701859473
transform -1 0 7270 0 1 7030
box -12 -8 32 272
use FILL  FILL_4__3017_
timestamp 1701859473
transform 1 0 6610 0 -1 7030
box -12 -8 32 272
use FILL  FILL_4__3018_
timestamp 1701859473
transform -1 0 6910 0 -1 7030
box -12 -8 32 272
use FILL  FILL_4__3019_
timestamp 1701859473
transform -1 0 7150 0 -1 7030
box -12 -8 32 272
use FILL  FILL_4__3020_
timestamp 1701859473
transform 1 0 8310 0 1 7030
box -12 -8 32 272
use FILL  FILL_4__3021_
timestamp 1701859473
transform -1 0 9370 0 -1 8070
box -12 -8 32 272
use FILL  FILL_4__3022_
timestamp 1701859473
transform 1 0 9550 0 -1 8070
box -12 -8 32 272
use FILL  FILL_4__3023_
timestamp 1701859473
transform -1 0 5770 0 1 6510
box -12 -8 32 272
use FILL  FILL_4__3024_
timestamp 1701859473
transform 1 0 5510 0 1 6510
box -12 -8 32 272
use FILL  FILL_4__3025_
timestamp 1701859473
transform -1 0 5530 0 -1 6510
box -12 -8 32 272
use FILL  FILL_4__3026_
timestamp 1701859473
transform 1 0 10950 0 -1 5990
box -12 -8 32 272
use FILL  FILL_4__3027_
timestamp 1701859473
transform -1 0 11190 0 -1 5990
box -12 -8 32 272
use FILL  FILL_4__3028_
timestamp 1701859473
transform -1 0 9810 0 -1 8070
box -12 -8 32 272
use FILL  FILL_4__3029_
timestamp 1701859473
transform -1 0 7130 0 -1 7550
box -12 -8 32 272
use FILL  FILL_4__3030_
timestamp 1701859473
transform -1 0 8110 0 -1 7030
box -12 -8 32 272
use FILL  FILL_4__3031_
timestamp 1701859473
transform 1 0 8090 0 1 7030
box -12 -8 32 272
use FILL  FILL_4__3032_
timestamp 1701859473
transform 1 0 7710 0 1 7550
box -12 -8 32 272
use FILL  FILL_4__3033_
timestamp 1701859473
transform -1 0 6790 0 1 8070
box -12 -8 32 272
use FILL  FILL_4__3034_
timestamp 1701859473
transform -1 0 7770 0 -1 8070
box -12 -8 32 272
use FILL  FILL_4__3035_
timestamp 1701859473
transform 1 0 7510 0 -1 8070
box -12 -8 32 272
use FILL  FILL_4__3036_
timestamp 1701859473
transform -1 0 6990 0 1 8070
box -12 -8 32 272
use FILL  FILL_4__3037_
timestamp 1701859473
transform -1 0 6550 0 1 8070
box -12 -8 32 272
use FILL  FILL_4__3038_
timestamp 1701859473
transform -1 0 7170 0 1 8070
box -12 -8 32 272
use FILL  FILL_4__3039_
timestamp 1701859473
transform 1 0 7390 0 1 8070
box -12 -8 32 272
use FILL  FILL_4__3040_
timestamp 1701859473
transform 1 0 9730 0 1 7550
box -12 -8 32 272
use FILL  FILL_4__3041_
timestamp 1701859473
transform -1 0 9590 0 -1 6510
box -12 -8 32 272
use FILL  FILL_4__3042_
timestamp 1701859473
transform 1 0 7290 0 -1 8070
box -12 -8 32 272
use FILL  FILL_4__3043_
timestamp 1701859473
transform -1 0 6610 0 1 7550
box -12 -8 32 272
use FILL  FILL_4__3044_
timestamp 1701859473
transform -1 0 6650 0 -1 7550
box -12 -8 32 272
use FILL  FILL_4__3045_
timestamp 1701859473
transform 1 0 6870 0 -1 7550
box -12 -8 32 272
use FILL  FILL_4__3046_
timestamp 1701859473
transform -1 0 7830 0 1 6510
box -12 -8 32 272
use FILL  FILL_4__3047_
timestamp 1701859473
transform 1 0 9170 0 1 6510
box -12 -8 32 272
use FILL  FILL_4__3048_
timestamp 1701859473
transform 1 0 9790 0 -1 6510
box -12 -8 32 272
use FILL  FILL_4__3049_
timestamp 1701859473
transform -1 0 6870 0 1 7550
box -12 -8 32 272
use FILL  FILL_4__3050_
timestamp 1701859473
transform -1 0 7090 0 1 7550
box -12 -8 32 272
use FILL  FILL_4__3051_
timestamp 1701859473
transform -1 0 7830 0 1 7030
box -12 -8 32 272
use FILL  FILL_4__3052_
timestamp 1701859473
transform 1 0 7530 0 1 7030
box -12 -8 32 272
use FILL  FILL_4__3053_
timestamp 1701859473
transform 1 0 7370 0 -1 7030
box -12 -8 32 272
use FILL  FILL_4__3054_
timestamp 1701859473
transform -1 0 7630 0 -1 7030
box -12 -8 32 272
use FILL  FILL_4__3055_
timestamp 1701859473
transform 1 0 8050 0 1 6510
box -12 -8 32 272
use FILL  FILL_4__3056_
timestamp 1701859473
transform -1 0 9570 0 1 5470
box -12 -8 32 272
use FILL  FILL_4__3057_
timestamp 1701859473
transform -1 0 9330 0 1 5470
box -12 -8 32 272
use FILL  FILL_4__3058_
timestamp 1701859473
transform 1 0 8750 0 -1 7550
box -12 -8 32 272
use FILL  FILL_4__3059_
timestamp 1701859473
transform -1 0 8630 0 -1 5990
box -12 -8 32 272
use FILL  FILL_4__3060_
timestamp 1701859473
transform 1 0 9810 0 1 6510
box -12 -8 32 272
use FILL  FILL_4__3061_
timestamp 1701859473
transform 1 0 10050 0 1 6510
box -12 -8 32 272
use FILL  FILL_4__3062_
timestamp 1701859473
transform -1 0 9670 0 -1 7550
box -12 -8 32 272
use FILL  FILL_4__3063_
timestamp 1701859473
transform 1 0 9410 0 -1 7550
box -12 -8 32 272
use FILL  FILL_4__3064_
timestamp 1701859473
transform -1 0 10370 0 -1 7030
box -12 -8 32 272
use FILL  FILL_4__3065_
timestamp 1701859473
transform -1 0 10610 0 -1 7030
box -12 -8 32 272
use FILL  FILL_4__3066_
timestamp 1701859473
transform -1 0 8530 0 -1 7550
box -12 -8 32 272
use FILL  FILL_4__3067_
timestamp 1701859473
transform 1 0 8270 0 -1 7550
box -12 -8 32 272
use FILL  FILL_4__3068_
timestamp 1701859473
transform 1 0 10230 0 -1 5990
box -12 -8 32 272
use FILL  FILL_4__3069_
timestamp 1701859473
transform 1 0 10470 0 -1 5990
box -12 -8 32 272
use FILL  FILL_4__3070_
timestamp 1701859473
transform 1 0 8930 0 -1 7550
box -12 -8 32 272
use FILL  FILL_4__3071_
timestamp 1701859473
transform -1 0 9190 0 -1 7550
box -12 -8 32 272
use FILL  FILL_4__3072_
timestamp 1701859473
transform -1 0 9810 0 1 5990
box -12 -8 32 272
use FILL  FILL_4__3073_
timestamp 1701859473
transform -1 0 10030 0 1 5990
box -12 -8 32 272
use FILL  FILL_4__3074_
timestamp 1701859473
transform 1 0 8850 0 1 5990
box -12 -8 32 272
use FILL  FILL_4__3075_
timestamp 1701859473
transform 1 0 8850 0 -1 5990
box -12 -8 32 272
use FILL  FILL_4__3076_
timestamp 1701859473
transform 1 0 10750 0 1 6510
box -12 -8 32 272
use FILL  FILL_4__3077_
timestamp 1701859473
transform 1 0 10950 0 1 6510
box -12 -8 32 272
use FILL  FILL_4__3078_
timestamp 1701859473
transform -1 0 8750 0 -1 7030
box -12 -8 32 272
use FILL  FILL_4__3079_
timestamp 1701859473
transform -1 0 8530 0 -1 7030
box -12 -8 32 272
use FILL  FILL_4__3080_
timestamp 1701859473
transform 1 0 11010 0 -1 8590
box -12 -8 32 272
use FILL  FILL_4__3081_
timestamp 1701859473
transform -1 0 11010 0 -1 270
box -12 -8 32 272
use FILL  FILL_4__3082_
timestamp 1701859473
transform 1 0 10110 0 -1 8590
box -12 -8 32 272
use FILL  FILL_4__3083_
timestamp 1701859473
transform -1 0 9890 0 -1 8590
box -12 -8 32 272
use FILL  FILL_4__3084_
timestamp 1701859473
transform -1 0 9070 0 1 7550
box -12 -8 32 272
use FILL  FILL_4__3085_
timestamp 1701859473
transform 1 0 8970 0 1 7030
box -12 -8 32 272
use FILL  FILL_4__3086_
timestamp 1701859473
transform -1 0 10730 0 1 5990
box -12 -8 32 272
use FILL  FILL_4__3087_
timestamp 1701859473
transform 1 0 10930 0 1 5990
box -12 -8 32 272
use FILL  FILL_4__3088_
timestamp 1701859473
transform 1 0 8290 0 1 8070
box -12 -8 32 272
use FILL  FILL_4__3089_
timestamp 1701859473
transform -1 0 8070 0 1 8070
box -12 -8 32 272
use FILL  FILL_4__3090_
timestamp 1701859473
transform -1 0 11170 0 1 4950
box -12 -8 32 272
use FILL  FILL_4__3091_
timestamp 1701859473
transform 1 0 10910 0 1 4950
box -12 -8 32 272
use FILL  FILL_4__3092_
timestamp 1701859473
transform 1 0 8830 0 -1 5470
box -12 -8 32 272
use FILL  FILL_4__3093_
timestamp 1701859473
transform -1 0 9070 0 -1 5470
box -12 -8 32 272
use FILL  FILL_4__3094_
timestamp 1701859473
transform -1 0 10270 0 -1 5470
box -12 -8 32 272
use FILL  FILL_4__3095_
timestamp 1701859473
transform 1 0 10210 0 1 5470
box -12 -8 32 272
use FILL  FILL_4__3096_
timestamp 1701859473
transform 1 0 8950 0 1 6510
box -12 -8 32 272
use FILL  FILL_4__3097_
timestamp 1701859473
transform -1 0 8730 0 1 6510
box -12 -8 32 272
use FILL  FILL_4__3098_
timestamp 1701859473
transform -1 0 10430 0 1 8070
box -12 -8 32 272
use FILL  FILL_4__3099_
timestamp 1701859473
transform -1 0 11190 0 -1 8070
box -12 -8 32 272
use FILL  FILL_4__3100_
timestamp 1701859473
transform 1 0 10190 0 1 8070
box -12 -8 32 272
use FILL  FILL_4__3101_
timestamp 1701859473
transform 1 0 10330 0 -1 8590
box -12 -8 32 272
use FILL  FILL_4__3102_
timestamp 1701859473
transform 1 0 8410 0 -1 8070
box -12 -8 32 272
use FILL  FILL_4__3103_
timestamp 1701859473
transform -1 0 8390 0 1 7550
box -12 -8 32 272
use FILL  FILL_4__3104_
timestamp 1701859473
transform -1 0 11190 0 1 6510
box -12 -8 32 272
use FILL  FILL_4__3105_
timestamp 1701859473
transform -1 0 10990 0 -1 4950
box -12 -8 32 272
use FILL  FILL_4__3106_
timestamp 1701859473
transform 1 0 9410 0 -1 8590
box -12 -8 32 272
use FILL  FILL_4__3107_
timestamp 1701859473
transform -1 0 9650 0 -1 8590
box -12 -8 32 272
use FILL  FILL_4__3108_
timestamp 1701859473
transform 1 0 10010 0 1 5470
box -12 -8 32 272
use FILL  FILL_4__3109_
timestamp 1701859473
transform -1 0 9790 0 1 5470
box -12 -8 32 272
use FILL  FILL_4__3110_
timestamp 1701859473
transform 1 0 8430 0 -1 6510
box -12 -8 32 272
use FILL  FILL_4__3111_
timestamp 1701859473
transform -1 0 8210 0 -1 6510
box -12 -8 32 272
use FILL  FILL_4__3112_
timestamp 1701859473
transform 1 0 550 0 -1 2870
box -12 -8 32 272
use FILL  FILL_4__3113_
timestamp 1701859473
transform 1 0 90 0 -1 2870
box -12 -8 32 272
use FILL  FILL_4__3114_
timestamp 1701859473
transform -1 0 350 0 -1 2870
box -12 -8 32 272
use FILL  FILL_4__3115_
timestamp 1701859473
transform -1 0 1230 0 1 2350
box -12 -8 32 272
use FILL  FILL_4__3116_
timestamp 1701859473
transform 1 0 990 0 -1 2350
box -12 -8 32 272
use FILL  FILL_4__3117_
timestamp 1701859473
transform 1 0 2070 0 -1 1310
box -12 -8 32 272
use FILL  FILL_4__3118_
timestamp 1701859473
transform -1 0 1450 0 -1 2350
box -12 -8 32 272
use FILL  FILL_4__3119_
timestamp 1701859473
transform -1 0 1210 0 -1 2350
box -12 -8 32 272
use FILL  FILL_4__3120_
timestamp 1701859473
transform -1 0 510 0 1 2350
box -12 -8 32 272
use FILL  FILL_4__3121_
timestamp 1701859473
transform 1 0 290 0 1 2870
box -12 -8 32 272
use FILL  FILL_4__3122_
timestamp 1701859473
transform 1 0 2550 0 -1 3390
box -12 -8 32 272
use FILL  FILL_4__3123_
timestamp 1701859473
transform 1 0 570 0 1 3390
box -12 -8 32 272
use FILL  FILL_4__3124_
timestamp 1701859473
transform -1 0 350 0 1 3390
box -12 -8 32 272
use FILL  FILL_4__3125_
timestamp 1701859473
transform -1 0 770 0 -1 2350
box -12 -8 32 272
use FILL  FILL_4__3126_
timestamp 1701859473
transform -1 0 1470 0 1 2350
box -12 -8 32 272
use FILL  FILL_4__3127_
timestamp 1701859473
transform -1 0 990 0 1 2350
box -12 -8 32 272
use FILL  FILL_4__3128_
timestamp 1701859473
transform -1 0 1930 0 1 2350
box -12 -8 32 272
use FILL  FILL_4__3129_
timestamp 1701859473
transform -1 0 1690 0 -1 2350
box -12 -8 32 272
use FILL  FILL_4__3130_
timestamp 1701859473
transform -1 0 1710 0 1 2350
box -12 -8 32 272
use FILL  FILL_4__3131_
timestamp 1701859473
transform -1 0 750 0 1 2350
box -12 -8 32 272
use FILL  FILL_4__3132_
timestamp 1701859473
transform 1 0 510 0 1 2870
box -12 -8 32 272
use FILL  FILL_4__3133_
timestamp 1701859473
transform 1 0 570 0 -1 3910
box -12 -8 32 272
use FILL  FILL_4__3134_
timestamp 1701859473
transform -1 0 1250 0 1 3390
box -12 -8 32 272
use FILL  FILL_4__3135_
timestamp 1701859473
transform 1 0 1010 0 1 3390
box -12 -8 32 272
use FILL  FILL_4__3136_
timestamp 1701859473
transform -1 0 590 0 -1 3390
box -12 -8 32 272
use FILL  FILL_4__3137_
timestamp 1701859473
transform 1 0 310 0 -1 3390
box -12 -8 32 272
use FILL  FILL_4__3138_
timestamp 1701859473
transform -1 0 1710 0 1 4430
box -12 -8 32 272
use FILL  FILL_4__3139_
timestamp 1701859473
transform -1 0 1910 0 -1 3390
box -12 -8 32 272
use FILL  FILL_4__3140_
timestamp 1701859473
transform -1 0 330 0 1 3910
box -12 -8 32 272
use FILL  FILL_4__3141_
timestamp 1701859473
transform 1 0 770 0 1 4430
box -12 -8 32 272
use FILL  FILL_4__3142_
timestamp 1701859473
transform 1 0 1010 0 1 4430
box -12 -8 32 272
use FILL  FILL_4__3143_
timestamp 1701859473
transform 1 0 1030 0 -1 4430
box -12 -8 32 272
use FILL  FILL_4__3144_
timestamp 1701859473
transform -1 0 1270 0 -1 4430
box -12 -8 32 272
use FILL  FILL_4__3145_
timestamp 1701859473
transform -1 0 550 0 1 3910
box -12 -8 32 272
use FILL  FILL_4__3146_
timestamp 1701859473
transform -1 0 770 0 1 3910
box -12 -8 32 272
use FILL  FILL_4__3147_
timestamp 1701859473
transform 1 0 550 0 -1 4430
box -12 -8 32 272
use FILL  FILL_4__3148_
timestamp 1701859473
transform -1 0 810 0 -1 4430
box -12 -8 32 272
use FILL  FILL_4__3149_
timestamp 1701859473
transform -1 0 110 0 -1 3910
box -12 -8 32 272
use FILL  FILL_4__3150_
timestamp 1701859473
transform -1 0 970 0 1 3910
box -12 -8 32 272
use FILL  FILL_4__3151_
timestamp 1701859473
transform 1 0 90 0 1 3910
box -12 -8 32 272
use FILL  FILL_4__3152_
timestamp 1701859473
transform 1 0 90 0 -1 4430
box -12 -8 32 272
use FILL  FILL_4__3153_
timestamp 1701859473
transform -1 0 330 0 -1 4430
box -12 -8 32 272
use FILL  FILL_4__3154_
timestamp 1701859473
transform -1 0 830 0 -1 3390
box -12 -8 32 272
use FILL  FILL_4__3155_
timestamp 1701859473
transform -1 0 110 0 1 2870
box -12 -8 32 272
use FILL  FILL_4__3156_
timestamp 1701859473
transform 1 0 90 0 -1 3390
box -12 -8 32 272
use FILL  FILL_4__3157_
timestamp 1701859473
transform -1 0 110 0 1 3390
box -12 -8 32 272
use FILL  FILL_4__3158_
timestamp 1701859473
transform 1 0 90 0 1 4430
box -12 -8 32 272
use FILL  FILL_4__3159_
timestamp 1701859473
transform 1 0 310 0 1 4430
box -12 -8 32 272
use FILL  FILL_4__3160_
timestamp 1701859473
transform -1 0 550 0 1 4430
box -12 -8 32 272
use FILL  FILL_4__3161_
timestamp 1701859473
transform 1 0 4190 0 -1 7030
box -12 -8 32 272
use FILL  FILL_4__3162_
timestamp 1701859473
transform -1 0 4430 0 -1 7030
box -12 -8 32 272
use FILL  FILL_4__3163_
timestamp 1701859473
transform 1 0 4650 0 -1 7030
box -12 -8 32 272
use FILL  FILL_4__3164_
timestamp 1701859473
transform 1 0 4890 0 1 7030
box -12 -8 32 272
use FILL  FILL_4__3165_
timestamp 1701859473
transform 1 0 4150 0 1 7550
box -12 -8 32 272
use FILL  FILL_4__3166_
timestamp 1701859473
transform -1 0 4390 0 1 7550
box -12 -8 32 272
use FILL  FILL_4__3167_
timestamp 1701859473
transform 1 0 4870 0 -1 10150
box -12 -8 32 272
use FILL  FILL_4__3168_
timestamp 1701859473
transform 1 0 5070 0 -1 10150
box -12 -8 32 272
use FILL  FILL_4__3169_
timestamp 1701859473
transform -1 0 3710 0 -1 10670
box -12 -8 32 272
use FILL  FILL_4__3170_
timestamp 1701859473
transform -1 0 3930 0 -1 10670
box -12 -8 32 272
use FILL  FILL_4__3171_
timestamp 1701859473
transform 1 0 4350 0 -1 10670
box -12 -8 32 272
use FILL  FILL_4__3172_
timestamp 1701859473
transform -1 0 4590 0 -1 10670
box -12 -8 32 272
use FILL  FILL_4__3173_
timestamp 1701859473
transform 1 0 4190 0 1 10150
box -12 -8 32 272
use FILL  FILL_4__3174_
timestamp 1701859473
transform -1 0 4430 0 1 10150
box -12 -8 32 272
use FILL  FILL_4__3175_
timestamp 1701859473
transform 1 0 5530 0 1 10150
box -12 -8 32 272
use FILL  FILL_4__3176_
timestamp 1701859473
transform 1 0 5290 0 1 10150
box -12 -8 32 272
use FILL  FILL_4__3177_
timestamp 1701859473
transform -1 0 1770 0 -1 5990
box -12 -8 32 272
use FILL  FILL_4__3178_
timestamp 1701859473
transform 1 0 2210 0 -1 5990
box -12 -8 32 272
use FILL  FILL_4__3179_
timestamp 1701859473
transform -1 0 1490 0 1 6510
box -12 -8 32 272
use FILL  FILL_4__3180_
timestamp 1701859473
transform -1 0 1710 0 1 6510
box -12 -8 32 272
use FILL  FILL_4__3181_
timestamp 1701859473
transform -1 0 570 0 -1 6510
box -12 -8 32 272
use FILL  FILL_4__3182_
timestamp 1701859473
transform -1 0 970 0 -1 6510
box -12 -8 32 272
use FILL  FILL_4__3183_
timestamp 1701859473
transform 1 0 330 0 1 8070
box -12 -8 32 272
use FILL  FILL_4__3184_
timestamp 1701859473
transform -1 0 570 0 1 8070
box -12 -8 32 272
use FILL  FILL_4__3185_
timestamp 1701859473
transform -1 0 110 0 -1 8590
box -12 -8 32 272
use FILL  FILL_4__3186_
timestamp 1701859473
transform -1 0 110 0 1 8070
box -12 -8 32 272
use FILL  FILL_4__3187_
timestamp 1701859473
transform 1 0 730 0 -1 9110
box -12 -8 32 272
use FILL  FILL_4__3188_
timestamp 1701859473
transform 1 0 950 0 -1 9110
box -12 -8 32 272
use FILL  FILL_4__3189_
timestamp 1701859473
transform 1 0 2130 0 -1 9630
box -12 -8 32 272
use FILL  FILL_4__3190_
timestamp 1701859473
transform 1 0 2370 0 1 9110
box -12 -8 32 272
use FILL  FILL_4__3191_
timestamp 1701859473
transform 1 0 1430 0 -1 9110
box -12 -8 32 272
use FILL  FILL_4__3192_
timestamp 1701859473
transform -1 0 1670 0 -1 9110
box -12 -8 32 272
use FILL  FILL_4__3324_
timestamp 1701859473
transform 1 0 5610 0 1 8070
box -12 -8 32 272
use FILL  FILL_4__3325_
timestamp 1701859473
transform -1 0 6330 0 1 8070
box -12 -8 32 272
use FILL  FILL_4__3326_
timestamp 1701859473
transform -1 0 6230 0 -1 8070
box -12 -8 32 272
use FILL  FILL_4__3327_
timestamp 1701859473
transform -1 0 6190 0 -1 8590
box -12 -8 32 272
use FILL  FILL_4__3328_
timestamp 1701859473
transform -1 0 6090 0 1 8070
box -12 -8 32 272
use FILL  FILL_4__3329_
timestamp 1701859473
transform 1 0 5850 0 1 8070
box -12 -8 32 272
use FILL  FILL_4__3330_
timestamp 1701859473
transform -1 0 7030 0 1 8590
box -12 -8 32 272
use FILL  FILL_4__3331_
timestamp 1701859473
transform 1 0 7310 0 -1 8590
box -12 -8 32 272
use FILL  FILL_4__3332_
timestamp 1701859473
transform 1 0 7030 0 -1 8590
box -12 -8 32 272
use FILL  FILL_4__3333_
timestamp 1701859473
transform 1 0 10230 0 1 8590
box -12 -8 32 272
use FILL  FILL_4__3334_
timestamp 1701859473
transform 1 0 9350 0 1 8590
box -12 -8 32 272
use FILL  FILL_4__3335_
timestamp 1701859473
transform 1 0 7890 0 -1 10150
box -12 -8 32 272
use FILL  FILL_4__3336_
timestamp 1701859473
transform -1 0 6730 0 1 9630
box -12 -8 32 272
use FILL  FILL_4__3337_
timestamp 1701859473
transform -1 0 6250 0 1 9630
box -12 -8 32 272
use FILL  FILL_4__3338_
timestamp 1701859473
transform 1 0 7210 0 -1 10150
box -12 -8 32 272
use FILL  FILL_4__3339_
timestamp 1701859473
transform -1 0 8090 0 1 10150
box -12 -8 32 272
use FILL  FILL_4__3340_
timestamp 1701859473
transform 1 0 7850 0 1 10150
box -12 -8 32 272
use FILL  FILL_4__3341_
timestamp 1701859473
transform 1 0 7610 0 1 10150
box -12 -8 32 272
use FILL  FILL_4__3342_
timestamp 1701859473
transform 1 0 6830 0 -1 11190
box -12 -8 32 272
use FILL  FILL_4__3343_
timestamp 1701859473
transform -1 0 7430 0 -1 10150
box -12 -8 32 272
use FILL  FILL_4__3344_
timestamp 1701859473
transform 1 0 7650 0 -1 10150
box -12 -8 32 272
use FILL  FILL_4__3345_
timestamp 1701859473
transform -1 0 9030 0 1 9630
box -12 -8 32 272
use FILL  FILL_4__3346_
timestamp 1701859473
transform 1 0 8550 0 1 10150
box -12 -8 32 272
use FILL  FILL_4__3347_
timestamp 1701859473
transform -1 0 8330 0 1 10150
box -12 -8 32 272
use FILL  FILL_4__3348_
timestamp 1701859473
transform 1 0 9150 0 -1 10670
box -12 -8 32 272
use FILL  FILL_4__3349_
timestamp 1701859473
transform 1 0 7890 0 1 9630
box -12 -8 32 272
use FILL  FILL_4__3350_
timestamp 1701859473
transform 1 0 7590 0 -1 8590
box -12 -8 32 272
use FILL  FILL_4__3351_
timestamp 1701859473
transform -1 0 7770 0 1 8590
box -12 -8 32 272
use FILL  FILL_4__3352_
timestamp 1701859473
transform -1 0 8230 0 -1 9110
box -12 -8 32 272
use FILL  FILL_4__3353_
timestamp 1701859473
transform 1 0 8110 0 -1 10150
box -12 -8 32 272
use FILL  FILL_4__3354_
timestamp 1701859473
transform 1 0 7790 0 -1 10670
box -12 -8 32 272
use FILL  FILL_4__3355_
timestamp 1701859473
transform -1 0 7570 0 -1 10670
box -12 -8 32 272
use FILL  FILL_4__3356_
timestamp 1701859473
transform 1 0 7350 0 -1 10670
box -12 -8 32 272
use FILL  FILL_4__3357_
timestamp 1701859473
transform 1 0 7170 0 1 10670
box -12 -8 32 272
use FILL  FILL_4__3358_
timestamp 1701859473
transform 1 0 7430 0 1 10670
box -12 -8 32 272
use FILL  FILL_4__3359_
timestamp 1701859473
transform 1 0 7670 0 1 10670
box -12 -8 32 272
use FILL  FILL_4__3360_
timestamp 1701859473
transform -1 0 7930 0 1 10670
box -12 -8 32 272
use FILL  FILL_4__3361_
timestamp 1701859473
transform 1 0 8950 0 -1 10670
box -12 -8 32 272
use FILL  FILL_4__3362_
timestamp 1701859473
transform 1 0 8010 0 -1 10670
box -12 -8 32 272
use FILL  FILL_4__3363_
timestamp 1701859473
transform 1 0 8130 0 1 10670
box -12 -8 32 272
use FILL  FILL_4__3364_
timestamp 1701859473
transform 1 0 7970 0 -1 11190
box -12 -8 32 272
use FILL  FILL_4__3365_
timestamp 1701859473
transform -1 0 7510 0 -1 11190
box -12 -8 32 272
use FILL  FILL_4__3366_
timestamp 1701859473
transform 1 0 7030 0 -1 11190
box -12 -8 32 272
use FILL  FILL_4__3367_
timestamp 1701859473
transform 1 0 6910 0 1 10670
box -12 -8 32 272
use FILL  FILL_4__3368_
timestamp 1701859473
transform 1 0 7250 0 -1 11190
box -12 -8 32 272
use FILL  FILL_4__3369_
timestamp 1701859473
transform 1 0 7730 0 -1 11190
box -12 -8 32 272
use FILL  FILL_4__3370_
timestamp 1701859473
transform 1 0 8250 0 -1 10670
box -12 -8 32 272
use FILL  FILL_4__3371_
timestamp 1701859473
transform 1 0 8350 0 1 10670
box -12 -8 32 272
use FILL  FILL_4__3372_
timestamp 1701859473
transform 1 0 9530 0 1 10670
box -12 -8 32 272
use FILL  FILL_4__3373_
timestamp 1701859473
transform -1 0 6630 0 -1 11190
box -12 -8 32 272
use FILL  FILL_4__3374_
timestamp 1701859473
transform 1 0 5730 0 1 10670
box -12 -8 32 272
use FILL  FILL_4__3375_
timestamp 1701859473
transform -1 0 5990 0 1 10670
box -12 -8 32 272
use FILL  FILL_4__3376_
timestamp 1701859473
transform -1 0 6210 0 1 10670
box -12 -8 32 272
use FILL  FILL_4__3377_
timestamp 1701859473
transform 1 0 6450 0 1 10670
box -12 -8 32 272
use FILL  FILL_4__3378_
timestamp 1701859473
transform 1 0 6390 0 -1 11190
box -12 -8 32 272
use FILL  FILL_4__3379_
timestamp 1701859473
transform 1 0 8710 0 -1 10670
box -12 -8 32 272
use FILL  FILL_4__3380_
timestamp 1701859473
transform 1 0 8830 0 1 10670
box -12 -8 32 272
use FILL  FILL_4__3381_
timestamp 1701859473
transform -1 0 6710 0 1 10670
box -12 -8 32 272
use FILL  FILL_4__3382_
timestamp 1701859473
transform 1 0 6170 0 -1 10670
box -12 -8 32 272
use FILL  FILL_4__3383_
timestamp 1701859473
transform -1 0 6430 0 -1 10670
box -12 -8 32 272
use FILL  FILL_4__3384_
timestamp 1701859473
transform -1 0 6870 0 -1 10670
box -12 -8 32 272
use FILL  FILL_4__3385_
timestamp 1701859473
transform 1 0 6630 0 -1 10670
box -12 -8 32 272
use FILL  FILL_4__3386_
timestamp 1701859473
transform 1 0 7110 0 -1 10670
box -12 -8 32 272
use FILL  FILL_4__3387_
timestamp 1701859473
transform 1 0 8470 0 -1 10670
box -12 -8 32 272
use FILL  FILL_4__3388_
timestamp 1701859473
transform 1 0 8590 0 1 10670
box -12 -8 32 272
use FILL  FILL_4__3389_
timestamp 1701859473
transform 1 0 10250 0 -1 10670
box -12 -8 32 272
use FILL  FILL_4__3390_
timestamp 1701859473
transform 1 0 9810 0 -1 10670
box -12 -8 32 272
use FILL  FILL_4__3391_
timestamp 1701859473
transform 1 0 10010 0 -1 10670
box -12 -8 32 272
use FILL  FILL_4__3392_
timestamp 1701859473
transform 1 0 10470 0 -1 10670
box -12 -8 32 272
use FILL  FILL_4__3393_
timestamp 1701859473
transform -1 0 11210 0 -1 10150
box -12 -8 32 272
use FILL  FILL_4__3394_
timestamp 1701859473
transform 1 0 7390 0 1 10150
box -12 -8 32 272
use FILL  FILL_4__3395_
timestamp 1701859473
transform 1 0 6450 0 1 10150
box -12 -8 32 272
use FILL  FILL_4__3396_
timestamp 1701859473
transform -1 0 6710 0 1 10150
box -12 -8 32 272
use FILL  FILL_4__3397_
timestamp 1701859473
transform -1 0 7030 0 -1 10150
box -12 -8 32 272
use FILL  FILL_4__3398_
timestamp 1701859473
transform 1 0 6310 0 -1 10150
box -12 -8 32 272
use FILL  FILL_4__3399_
timestamp 1701859473
transform -1 0 6790 0 -1 10150
box -12 -8 32 272
use FILL  FILL_4__3400_
timestamp 1701859473
transform -1 0 6970 0 1 10150
box -12 -8 32 272
use FILL  FILL_4__3401_
timestamp 1701859473
transform 1 0 7150 0 1 10150
box -12 -8 32 272
use FILL  FILL_4__3402_
timestamp 1701859473
transform -1 0 9090 0 1 10150
box -12 -8 32 272
use FILL  FILL_4__3403_
timestamp 1701859473
transform 1 0 9530 0 1 10150
box -12 -8 32 272
use FILL  FILL_4__3404_
timestamp 1701859473
transform -1 0 5790 0 1 9630
box -12 -8 32 272
use FILL  FILL_4__3405_
timestamp 1701859473
transform -1 0 6070 0 -1 10150
box -12 -8 32 272
use FILL  FILL_4__3406_
timestamp 1701859473
transform 1 0 6430 0 -1 9630
box -12 -8 32 272
use FILL  FILL_4__3407_
timestamp 1701859473
transform -1 0 6650 0 -1 9630
box -12 -8 32 272
use FILL  FILL_4__3408_
timestamp 1701859473
transform 1 0 6910 0 1 9630
box -12 -8 32 272
use FILL  FILL_4__3409_
timestamp 1701859473
transform -1 0 6530 0 -1 10150
box -12 -8 32 272
use FILL  FILL_4__3410_
timestamp 1701859473
transform 1 0 9270 0 -1 10150
box -12 -8 32 272
use FILL  FILL_4__3411_
timestamp 1701859473
transform 1 0 9290 0 1 10150
box -12 -8 32 272
use FILL  FILL_4__3412_
timestamp 1701859473
transform 1 0 10010 0 1 10150
box -12 -8 32 272
use FILL  FILL_4__3413_
timestamp 1701859473
transform -1 0 6030 0 1 9630
box -12 -8 32 272
use FILL  FILL_4__3414_
timestamp 1701859473
transform 1 0 8170 0 1 9110
box -12 -8 32 272
use FILL  FILL_4__3415_
timestamp 1701859473
transform 1 0 6450 0 1 9630
box -12 -8 32 272
use FILL  FILL_4__3416_
timestamp 1701859473
transform 1 0 7290 0 1 8590
box -12 -8 32 272
use FILL  FILL_4__3417_
timestamp 1701859473
transform 1 0 7370 0 -1 9110
box -12 -8 32 272
use FILL  FILL_4__3418_
timestamp 1701859473
transform -1 0 7510 0 -1 9630
box -12 -8 32 272
use FILL  FILL_4__3419_
timestamp 1701859473
transform 1 0 7270 0 -1 9630
box -12 -8 32 272
use FILL  FILL_4__3420_
timestamp 1701859473
transform -1 0 6850 0 -1 9630
box -12 -8 32 272
use FILL  FILL_4__3421_
timestamp 1701859473
transform -1 0 7070 0 -1 9630
box -12 -8 32 272
use FILL  FILL_4__3422_
timestamp 1701859473
transform -1 0 7170 0 1 9630
box -12 -8 32 272
use FILL  FILL_4__3423_
timestamp 1701859473
transform -1 0 8230 0 -1 9630
box -12 -8 32 272
use FILL  FILL_4__3424_
timestamp 1701859473
transform -1 0 7750 0 -1 9630
box -12 -8 32 272
use FILL  FILL_4__3425_
timestamp 1701859473
transform -1 0 7410 0 1 9630
box -12 -8 32 272
use FILL  FILL_4__3426_
timestamp 1701859473
transform -1 0 9050 0 -1 10150
box -12 -8 32 272
use FILL  FILL_4__3427_
timestamp 1701859473
transform 1 0 8810 0 -1 10150
box -12 -8 32 272
use FILL  FILL_4__3428_
timestamp 1701859473
transform 1 0 7490 0 1 8590
box -12 -8 32 272
use FILL  FILL_4__3429_
timestamp 1701859473
transform 1 0 7570 0 -1 9110
box -12 -8 32 272
use FILL  FILL_4__3430_
timestamp 1701859473
transform -1 0 7790 0 -1 9110
box -12 -8 32 272
use FILL  FILL_4__3431_
timestamp 1701859473
transform 1 0 7710 0 1 9110
box -12 -8 32 272
use FILL  FILL_4__3432_
timestamp 1701859473
transform 1 0 7950 0 1 9110
box -12 -8 32 272
use FILL  FILL_4__3433_
timestamp 1701859473
transform -1 0 7990 0 -1 9630
box -12 -8 32 272
use FILL  FILL_4__3434_
timestamp 1701859473
transform 1 0 7630 0 1 9630
box -12 -8 32 272
use FILL  FILL_4__3435_
timestamp 1701859473
transform 1 0 10250 0 1 10150
box -12 -8 32 272
use FILL  FILL_4__3436_
timestamp 1701859473
transform -1 0 10250 0 -1 10150
box -12 -8 32 272
use FILL  FILL_4__3437_
timestamp 1701859473
transform 1 0 10690 0 1 10150
box -12 -8 32 272
use FILL  FILL_4__3438_
timestamp 1701859473
transform 1 0 10470 0 1 10150
box -12 -8 32 272
use FILL  FILL_4__3439_
timestamp 1701859473
transform 1 0 10910 0 1 10150
box -12 -8 32 272
use FILL  FILL_4__3440_
timestamp 1701859473
transform -1 0 10730 0 -1 10150
box -12 -8 32 272
use FILL  FILL_4__3441_
timestamp 1701859473
transform -1 0 10590 0 1 9630
box -12 -8 32 272
use FILL  FILL_4__3442_
timestamp 1701859473
transform -1 0 10470 0 -1 10150
box -12 -8 32 272
use FILL  FILL_4__3443_
timestamp 1701859473
transform -1 0 11030 0 1 9630
box -12 -8 32 272
use FILL  FILL_4__3444_
timestamp 1701859473
transform -1 0 8430 0 -1 9630
box -12 -8 32 272
use FILL  FILL_4__3445_
timestamp 1701859473
transform -1 0 8130 0 1 9630
box -12 -8 32 272
use FILL  FILL_4__3446_
timestamp 1701859473
transform 1 0 8570 0 1 9630
box -12 -8 32 272
use FILL  FILL_4__3447_
timestamp 1701859473
transform 1 0 8350 0 1 9630
box -12 -8 32 272
use FILL  FILL_4__3448_
timestamp 1701859473
transform -1 0 8790 0 1 9630
box -12 -8 32 272
use FILL  FILL_4__3449_
timestamp 1701859473
transform -1 0 9830 0 1 10150
box -12 -8 32 272
use FILL  FILL_4__3450_
timestamp 1701859473
transform -1 0 9790 0 -1 10150
box -12 -8 32 272
use FILL  FILL_4__3451_
timestamp 1701859473
transform 1 0 9510 0 -1 10150
box -12 -8 32 272
use FILL  FILL_4__3452_
timestamp 1701859473
transform -1 0 9250 0 1 9630
box -12 -8 32 272
use FILL  FILL_4__3453_
timestamp 1701859473
transform -1 0 10010 0 -1 10150
box -12 -8 32 272
use FILL  FILL_4__3454_
timestamp 1701859473
transform 1 0 9450 0 1 9630
box -12 -8 32 272
use FILL  FILL_4__3455_
timestamp 1701859473
transform 1 0 9670 0 1 9630
box -12 -8 32 272
use FILL  FILL_4__3456_
timestamp 1701859473
transform -1 0 10370 0 1 9630
box -12 -8 32 272
use FILL  FILL_4__3457_
timestamp 1701859473
transform -1 0 9910 0 1 9630
box -12 -8 32 272
use FILL  FILL_4__3458_
timestamp 1701859473
transform -1 0 10150 0 1 9630
box -12 -8 32 272
use FILL  FILL_4__3459_
timestamp 1701859473
transform -1 0 10290 0 -1 9630
box -12 -8 32 272
use FILL  FILL_4__3460_
timestamp 1701859473
transform 1 0 10950 0 -1 10150
box -12 -8 32 272
use FILL  FILL_4__3461_
timestamp 1701859473
transform -1 0 11190 0 -1 9630
box -12 -8 32 272
use FILL  FILL_4__3462_
timestamp 1701859473
transform -1 0 10730 0 -1 9630
box -12 -8 32 272
use FILL  FILL_4__3463_
timestamp 1701859473
transform 1 0 10410 0 -1 11190
box -12 -8 32 272
use FILL  FILL_4__3464_
timestamp 1701859473
transform 1 0 9750 0 -1 11190
box -12 -8 32 272
use FILL  FILL_4__3465_
timestamp 1701859473
transform 1 0 9990 0 -1 11190
box -12 -8 32 272
use FILL  FILL_4__3466_
timestamp 1701859473
transform 1 0 10170 0 -1 11190
box -12 -8 32 272
use FILL  FILL_4__3467_
timestamp 1701859473
transform -1 0 11150 0 1 10670
box -12 -8 32 272
use FILL  FILL_4__3468_
timestamp 1701859473
transform 1 0 10650 0 1 10670
box -12 -8 32 272
use FILL  FILL_4__3469_
timestamp 1701859473
transform 1 0 9370 0 -1 10670
box -12 -8 32 272
use FILL  FILL_4__3470_
timestamp 1701859473
transform 1 0 9610 0 -1 10670
box -12 -8 32 272
use FILL  FILL_4__3471_
timestamp 1701859473
transform 1 0 9750 0 1 10670
box -12 -8 32 272
use FILL  FILL_4__3472_
timestamp 1701859473
transform -1 0 10010 0 1 10670
box -12 -8 32 272
use FILL  FILL_4__3473_
timestamp 1701859473
transform 1 0 8630 0 -1 11190
box -12 -8 32 272
use FILL  FILL_4__3474_
timestamp 1701859473
transform 1 0 8190 0 -1 11190
box -12 -8 32 272
use FILL  FILL_4__3475_
timestamp 1701859473
transform 1 0 8430 0 -1 11190
box -12 -8 32 272
use FILL  FILL_4__3476_
timestamp 1701859473
transform -1 0 8870 0 -1 11190
box -12 -8 32 272
use FILL  FILL_4__3477_
timestamp 1701859473
transform 1 0 9090 0 -1 11190
box -12 -8 32 272
use FILL  FILL_4__3478_
timestamp 1701859473
transform 1 0 9070 0 1 10670
box -12 -8 32 272
use FILL  FILL_4__3479_
timestamp 1701859473
transform 1 0 8350 0 -1 10150
box -12 -8 32 272
use FILL  FILL_4__3480_
timestamp 1701859473
transform -1 0 8610 0 -1 10150
box -12 -8 32 272
use FILL  FILL_4__3481_
timestamp 1701859473
transform -1 0 8390 0 1 9110
box -12 -8 32 272
use FILL  FILL_4__3482_
timestamp 1701859473
transform -1 0 8610 0 1 9110
box -12 -8 32 272
use FILL  FILL_4__3483_
timestamp 1701859473
transform 1 0 8790 0 1 10150
box -12 -8 32 272
use FILL  FILL_4__3484_
timestamp 1701859473
transform -1 0 10090 0 -1 9630
box -12 -8 32 272
use FILL  FILL_4__3485_
timestamp 1701859473
transform 1 0 11110 0 1 10150
box -12 -8 32 272
use FILL  FILL_4__3486_
timestamp 1701859473
transform 1 0 10450 0 1 9110
box -12 -8 32 272
use FILL  FILL_4__3487_
timestamp 1701859473
transform 1 0 10490 0 -1 9630
box -12 -8 32 272
use FILL  FILL_4__3488_
timestamp 1701859473
transform -1 0 10790 0 1 9630
box -12 -8 32 272
use FILL  FILL_4__3489_
timestamp 1701859473
transform 1 0 10630 0 -1 11190
box -12 -8 32 272
use FILL  FILL_4__3490_
timestamp 1701859473
transform 1 0 11090 0 -1 11190
box -12 -8 32 272
use FILL  FILL_4__3491_
timestamp 1701859473
transform -1 0 10890 0 -1 11190
box -12 -8 32 272
use FILL  FILL_4__3492_
timestamp 1701859473
transform -1 0 10450 0 1 10670
box -12 -8 32 272
use FILL  FILL_4__3493_
timestamp 1701859473
transform -1 0 10230 0 1 10670
box -12 -8 32 272
use FILL  FILL_4__3494_
timestamp 1701859473
transform 1 0 9330 0 1 10670
box -12 -8 32 272
use FILL  FILL_4__3495_
timestamp 1701859473
transform -1 0 9530 0 -1 11190
box -12 -8 32 272
use FILL  FILL_4__3496_
timestamp 1701859473
transform 1 0 9290 0 -1 11190
box -12 -8 32 272
use FILL  FILL_4__3497_
timestamp 1701859473
transform -1 0 9390 0 -1 9630
box -12 -8 32 272
use FILL  FILL_4__3498_
timestamp 1701859473
transform -1 0 8890 0 1 9110
box -12 -8 32 272
use FILL  FILL_4__3499_
timestamp 1701859473
transform 1 0 8410 0 -1 9110
box -12 -8 32 272
use FILL  FILL_4__3500_
timestamp 1701859473
transform 1 0 9790 0 1 9110
box -12 -8 32 272
use FILL  FILL_4__3501_
timestamp 1701859473
transform -1 0 10030 0 1 9110
box -12 -8 32 272
use FILL  FILL_4__3502_
timestamp 1701859473
transform -1 0 8290 0 -1 8590
box -12 -8 32 272
use FILL  FILL_4__3503_
timestamp 1701859473
transform -1 0 8670 0 -1 9630
box -12 -8 32 272
use FILL  FILL_4__3504_
timestamp 1701859473
transform 1 0 8890 0 -1 9630
box -12 -8 32 272
use FILL  FILL_4__3505_
timestamp 1701859473
transform -1 0 9150 0 -1 9630
box -12 -8 32 272
use FILL  FILL_4__3506_
timestamp 1701859473
transform -1 0 8670 0 1 8590
box -12 -8 32 272
use FILL  FILL_4__3507_
timestamp 1701859473
transform 1 0 10750 0 -1 9110
box -12 -8 32 272
use FILL  FILL_4__3508_
timestamp 1701859473
transform 1 0 10510 0 -1 9110
box -12 -8 32 272
use FILL  FILL_4__3509_
timestamp 1701859473
transform 1 0 8450 0 1 8590
box -12 -8 32 272
use FILL  FILL_4__3510_
timestamp 1701859473
transform -1 0 8910 0 1 8590
box -12 -8 32 272
use FILL  FILL_4__3511_
timestamp 1701859473
transform 1 0 9970 0 -1 270
box -12 -8 32 272
use FILL  FILL_4__3512_
timestamp 1701859473
transform 1 0 10970 0 -1 9110
box -12 -8 32 272
use FILL  FILL_4__3513_
timestamp 1701859473
transform 1 0 10950 0 -1 9630
box -12 -8 32 272
use FILL  FILL_4__3514_
timestamp 1701859473
transform 1 0 10910 0 1 10670
box -12 -8 32 272
use FILL  FILL_4__3515_
timestamp 1701859473
transform -1 0 10710 0 -1 10670
box -12 -8 32 272
use FILL  FILL_4__3516_
timestamp 1701859473
transform 1 0 10930 0 -1 10670
box -12 -8 32 272
use FILL  FILL_4__3517_
timestamp 1701859473
transform 1 0 9610 0 -1 9630
box -12 -8 32 272
use FILL  FILL_4__3518_
timestamp 1701859473
transform 1 0 9830 0 -1 9630
box -12 -8 32 272
use FILL  FILL_4__3519_
timestamp 1701859473
transform 1 0 9110 0 1 9110
box -12 -8 32 272
use FILL  FILL_4__3520_
timestamp 1701859473
transform -1 0 9350 0 1 9110
box -12 -8 32 272
use FILL  FILL_4__3521_
timestamp 1701859473
transform 1 0 6590 0 1 8590
box -12 -8 32 272
use FILL  FILL_4__3522_
timestamp 1701859473
transform 1 0 7990 0 -1 9110
box -12 -8 32 272
use FILL  FILL_4__3523_
timestamp 1701859473
transform 1 0 6790 0 1 8590
box -12 -8 32 272
use FILL  FILL_4__3524_
timestamp 1701859473
transform 1 0 7510 0 1 9110
box -12 -8 32 272
use FILL  FILL_4__3525_
timestamp 1701859473
transform 1 0 7050 0 1 9110
box -12 -8 32 272
use FILL  FILL_4__3526_
timestamp 1701859473
transform -1 0 7290 0 1 9110
box -12 -8 32 272
use FILL  FILL_4__3539_
timestamp 1701859473
transform 1 0 11150 0 -1 7030
box -12 -8 32 272
use FILL  FILL_4__3540_
timestamp 1701859473
transform 1 0 4650 0 1 10670
box -12 -8 32 272
use FILL  FILL_4__3541_
timestamp 1701859473
transform -1 0 110 0 1 5990
box -12 -8 32 272
use FILL  FILL_4__3542_
timestamp 1701859473
transform -1 0 110 0 -1 8070
box -12 -8 32 272
use FILL  FILL_4__3543_
timestamp 1701859473
transform -1 0 110 0 1 8590
box -12 -8 32 272
use FILL  FILL_4__3544_
timestamp 1701859473
transform -1 0 110 0 1 9110
box -12 -8 32 272
use FILL  FILL_4__3545_
timestamp 1701859473
transform -1 0 1950 0 -1 11190
box -12 -8 32 272
use FILL  FILL_4__3546_
timestamp 1701859473
transform -1 0 570 0 1 9110
box -12 -8 32 272
use FILL  FILL_4__3547_
timestamp 1701859473
transform 1 0 4690 0 -1 11190
box -12 -8 32 272
use FILL  FILL_4__3548_
timestamp 1701859473
transform 1 0 5290 0 1 10670
box -12 -8 32 272
use FILL  FILL_4__3549_
timestamp 1701859473
transform -1 0 4290 0 -1 11190
box -12 -8 32 272
use FILL  FILL_4__3550_
timestamp 1701859473
transform -1 0 5130 0 -1 11190
box -12 -8 32 272
use FILL  FILL_4__3551_
timestamp 1701859473
transform 1 0 5530 0 -1 11190
box -12 -8 32 272
use FILL  FILL_4__3552_
timestamp 1701859473
transform 1 0 5310 0 -1 11190
box -12 -8 32 272
use FILL  FILL_4__3553_
timestamp 1701859473
transform -1 0 110 0 -1 5990
box -12 -8 32 272
use FILL  FILL_4__3554_
timestamp 1701859473
transform -1 0 310 0 1 7030
box -12 -8 32 272
use FILL  FILL_4__3555_
timestamp 1701859473
transform -1 0 5090 0 1 10670
box -12 -8 32 272
use FILL  FILL_4__3556_
timestamp 1701859473
transform 1 0 6230 0 1 10150
box -12 -8 32 272
use FILL  FILL_4__3557_
timestamp 1701859473
transform -1 0 5770 0 -1 11190
box -12 -8 32 272
use FILL  FILL_4__3558_
timestamp 1701859473
transform 1 0 6170 0 -1 11190
box -12 -8 32 272
use FILL  FILL_4__3559_
timestamp 1701859473
transform -1 0 4830 0 -1 10670
box -12 -8 32 272
use FILL  FILL_4__3560_
timestamp 1701859473
transform 1 0 5510 0 1 10670
box -12 -8 32 272
use FILL  FILL_4__3561_
timestamp 1701859473
transform 1 0 5950 0 -1 11190
box -12 -8 32 272
use FILL  FILL_4__3562_
timestamp 1701859473
transform 1 0 5750 0 1 10150
box -12 -8 32 272
use FILL  FILL_4__3563_
timestamp 1701859473
transform 1 0 5210 0 1 3390
box -12 -8 32 272
use FILL  FILL_4_BUFX2_insert0
timestamp 1701859473
transform 1 0 5830 0 -1 10150
box -12 -8 32 272
use FILL  FILL_4_BUFX2_insert1
timestamp 1701859473
transform 1 0 6590 0 1 2350
box -12 -8 32 272
use FILL  FILL_4_BUFX2_insert2
timestamp 1701859473
transform 1 0 5430 0 -1 1830
box -12 -8 32 272
use FILL  FILL_4_BUFX2_insert3
timestamp 1701859473
transform -1 0 570 0 -1 5470
box -12 -8 32 272
use FILL  FILL_4_BUFX2_insert4
timestamp 1701859473
transform 1 0 3310 0 1 4950
box -12 -8 32 272
use FILL  FILL_4_BUFX2_insert5
timestamp 1701859473
transform 1 0 1370 0 -1 1830
box -12 -8 32 272
use FILL  FILL_4_BUFX2_insert6
timestamp 1701859473
transform -1 0 110 0 -1 11190
box -12 -8 32 272
use FILL  FILL_4_BUFX2_insert7
timestamp 1701859473
transform 1 0 1670 0 1 10670
box -12 -8 32 272
use FILL  FILL_4_BUFX2_insert8
timestamp 1701859473
transform 1 0 1630 0 1 1830
box -12 -8 32 272
use FILL  FILL_4_BUFX2_insert9
timestamp 1701859473
transform 1 0 1930 0 -1 3910
box -12 -8 32 272
use FILL  FILL_4_BUFX2_insert10
timestamp 1701859473
transform 1 0 1750 0 -1 4430
box -12 -8 32 272
use FILL  FILL_4_BUFX2_insert11
timestamp 1701859473
transform -1 0 1730 0 -1 3910
box -12 -8 32 272
use FILL  FILL_4_BUFX2_insert12
timestamp 1701859473
transform -1 0 1510 0 -1 3910
box -12 -8 32 272
use FILL  FILL_4_BUFX2_insert13
timestamp 1701859473
transform -1 0 1410 0 -1 1310
box -12 -8 32 272
use FILL  FILL_4_BUFX2_insert14
timestamp 1701859473
transform -1 0 3650 0 1 3390
box -12 -8 32 272
use FILL  FILL_4_BUFX2_insert15
timestamp 1701859473
transform 1 0 4530 0 -1 5470
box -12 -8 32 272
use FILL  FILL_4_BUFX2_insert16
timestamp 1701859473
transform 1 0 1330 0 -1 4950
box -12 -8 32 272
use FILL  FILL_4_BUFX2_insert17
timestamp 1701859473
transform 1 0 3610 0 1 1310
box -12 -8 32 272
use FILL  FILL_4_BUFX2_insert18
timestamp 1701859473
transform -1 0 9750 0 1 2350
box -12 -8 32 272
use FILL  FILL_4_BUFX2_insert19
timestamp 1701859473
transform -1 0 8490 0 -1 790
box -12 -8 32 272
use FILL  FILL_4_BUFX2_insert20
timestamp 1701859473
transform 1 0 9950 0 1 2350
box -12 -8 32 272
use FILL  FILL_4_BUFX2_insert21
timestamp 1701859473
transform -1 0 7790 0 -1 1310
box -12 -8 32 272
use FILL  FILL_4_BUFX2_insert22
timestamp 1701859473
transform -1 0 3190 0 -1 2870
box -12 -8 32 272
use FILL  FILL_4_BUFX2_insert23
timestamp 1701859473
transform -1 0 2730 0 -1 4950
box -12 -8 32 272
use FILL  FILL_4_BUFX2_insert24
timestamp 1701859473
transform -1 0 3630 0 -1 4430
box -12 -8 32 272
use FILL  FILL_4_BUFX2_insert25
timestamp 1701859473
transform 1 0 4370 0 1 4430
box -12 -8 32 272
use FILL  FILL_4_BUFX2_insert26
timestamp 1701859473
transform 1 0 4190 0 1 2870
box -12 -8 32 272
use FILL  FILL_4_BUFX2_insert27
timestamp 1701859473
transform 1 0 9590 0 1 4950
box -12 -8 32 272
use FILL  FILL_4_BUFX2_insert28
timestamp 1701859473
transform -1 0 7470 0 -1 5990
box -12 -8 32 272
use FILL  FILL_4_BUFX2_insert29
timestamp 1701859473
transform -1 0 1270 0 1 6510
box -12 -8 32 272
use FILL  FILL_4_BUFX2_insert30
timestamp 1701859473
transform -1 0 8770 0 -1 3910
box -12 -8 32 272
use FILL  FILL_4_BUFX2_insert31
timestamp 1701859473
transform -1 0 9550 0 1 3910
box -12 -8 32 272
use FILL  FILL_4_BUFX2_insert32
timestamp 1701859473
transform 1 0 5850 0 -1 3910
box -12 -8 32 272
use FILL  FILL_4_BUFX2_insert33
timestamp 1701859473
transform -1 0 9530 0 -1 4950
box -12 -8 32 272
use FILL  FILL_4_BUFX2_insert34
timestamp 1701859473
transform 1 0 5190 0 1 8590
box -12 -8 32 272
use FILL  FILL_4_BUFX2_insert35
timestamp 1701859473
transform -1 0 5950 0 1 7550
box -12 -8 32 272
use FILL  FILL_4_BUFX2_insert36
timestamp 1701859473
transform -1 0 1190 0 1 8590
box -12 -8 32 272
use FILL  FILL_4_BUFX2_insert37
timestamp 1701859473
transform -1 0 9570 0 1 8590
box -12 -8 32 272
use FILL  FILL_4_BUFX2_insert49
timestamp 1701859473
transform -1 0 3030 0 1 6510
box -12 -8 32 272
use FILL  FILL_4_BUFX2_insert50
timestamp 1701859473
transform 1 0 2330 0 -1 8590
box -12 -8 32 272
use FILL  FILL_4_BUFX2_insert51
timestamp 1701859473
transform 1 0 3190 0 -1 8590
box -12 -8 32 272
use FILL  FILL_4_BUFX2_insert52
timestamp 1701859473
transform 1 0 3370 0 1 5470
box -12 -8 32 272
use FILL  FILL_4_BUFX2_insert53
timestamp 1701859473
transform -1 0 11210 0 1 9110
box -12 -8 32 272
use FILL  FILL_4_BUFX2_insert54
timestamp 1701859473
transform -1 0 9150 0 1 8590
box -12 -8 32 272
use FILL  FILL_4_BUFX2_insert55
timestamp 1701859473
transform -1 0 9590 0 1 9110
box -12 -8 32 272
use FILL  FILL_4_BUFX2_insert56
timestamp 1701859473
transform -1 0 10250 0 1 9110
box -12 -8 32 272
use FILL  FILL_4_BUFX2_insert57
timestamp 1701859473
transform -1 0 11210 0 -1 2350
box -12 -8 32 272
use FILL  FILL_4_BUFX2_insert58
timestamp 1701859473
transform -1 0 8950 0 1 2870
box -12 -8 32 272
use FILL  FILL_4_BUFX2_insert59
timestamp 1701859473
transform -1 0 7530 0 1 1830
box -12 -8 32 272
use FILL  FILL_4_BUFX2_insert60
timestamp 1701859473
transform 1 0 10870 0 1 1830
box -12 -8 32 272
use FILL  FILL_4_BUFX2_insert61
timestamp 1701859473
transform -1 0 11150 0 1 2870
box -12 -8 32 272
use FILL  FILL_4_BUFX2_insert62
timestamp 1701859473
transform 1 0 2190 0 1 3910
box -12 -8 32 272
use FILL  FILL_4_BUFX2_insert63
timestamp 1701859473
transform 1 0 2110 0 1 3390
box -12 -8 32 272
use FILL  FILL_4_BUFX2_insert64
timestamp 1701859473
transform -1 0 1770 0 1 3910
box -12 -8 32 272
use FILL  FILL_4_BUFX2_insert65
timestamp 1701859473
transform -1 0 1710 0 1 3390
box -12 -8 32 272
use FILL  FILL_4_BUFX2_insert66
timestamp 1701859473
transform -1 0 4290 0 1 1310
box -12 -8 32 272
use FILL  FILL_4_BUFX2_insert67
timestamp 1701859473
transform -1 0 3590 0 -1 10150
box -12 -8 32 272
use FILL  FILL_4_BUFX2_insert68
timestamp 1701859473
transform -1 0 7150 0 1 2870
box -12 -8 32 272
use FILL  FILL_4_BUFX2_insert69
timestamp 1701859473
transform -1 0 5630 0 -1 3390
box -12 -8 32 272
use FILL  FILL_4_BUFX2_insert70
timestamp 1701859473
transform -1 0 3650 0 -1 1830
box -12 -8 32 272
use FILL  FILL_4_BUFX2_insert71
timestamp 1701859473
transform -1 0 7290 0 1 2350
box -12 -8 32 272
use FILL  FILL_4_BUFX2_insert72
timestamp 1701859473
transform -1 0 6470 0 1 1310
box -12 -8 32 272
use FILL  FILL_4_BUFX2_insert73
timestamp 1701859473
transform 1 0 3590 0 1 5470
box -12 -8 32 272
use FILL  FILL_4_BUFX2_insert74
timestamp 1701859473
transform 1 0 7550 0 -1 2350
box -12 -8 32 272
use FILL  FILL_4_BUFX2_insert75
timestamp 1701859473
transform 1 0 7570 0 1 2870
box -12 -8 32 272
use FILL  FILL_4_BUFX2_insert76
timestamp 1701859473
transform 1 0 7350 0 1 2870
box -12 -8 32 272
use FILL  FILL_4_BUFX2_insert77
timestamp 1701859473
transform -1 0 3410 0 -1 2870
box -12 -8 32 272
use FILL  FILL_4_BUFX2_insert78
timestamp 1701859473
transform 1 0 1910 0 -1 2870
box -12 -8 32 272
use FILL  FILL_4_BUFX2_insert79
timestamp 1701859473
transform -1 0 2150 0 -1 2870
box -12 -8 32 272
use FILL  FILL_4_BUFX2_insert80
timestamp 1701859473
transform 1 0 2390 0 1 4430
box -12 -8 32 272
use FILL  FILL_4_BUFX2_insert81
timestamp 1701859473
transform -1 0 1990 0 1 3910
box -12 -8 32 272
use FILL  FILL_4_BUFX2_insert82
timestamp 1701859473
transform -1 0 310 0 1 8590
box -12 -8 32 272
use FILL  FILL_4_BUFX2_insert83
timestamp 1701859473
transform 1 0 4190 0 -1 10150
box -12 -8 32 272
use FILL  FILL_4_BUFX2_insert84
timestamp 1701859473
transform 1 0 4150 0 -1 7550
box -12 -8 32 272
use FILL  FILL_4_BUFX2_insert85
timestamp 1701859473
transform -1 0 110 0 -1 6510
box -12 -8 32 272
use FILL  FILL_4_BUFX2_insert86
timestamp 1701859473
transform 1 0 1910 0 -1 10150
box -12 -8 32 272
use FILL  FILL_4_CLKBUF1_insert38
timestamp 1701859473
transform 1 0 2910 0 -1 7550
box -12 -8 32 272
use FILL  FILL_4_CLKBUF1_insert39
timestamp 1701859473
transform -1 0 4710 0 -1 6510
box -12 -8 32 272
use FILL  FILL_4_CLKBUF1_insert40
timestamp 1701859473
transform -1 0 1010 0 -1 4950
box -12 -8 32 272
use FILL  FILL_4_CLKBUF1_insert41
timestamp 1701859473
transform -1 0 10670 0 -1 270
box -12 -8 32 272
use FILL  FILL_4_CLKBUF1_insert42
timestamp 1701859473
transform 1 0 9730 0 -1 4950
box -12 -8 32 272
use FILL  FILL_4_CLKBUF1_insert43
timestamp 1701859473
transform -1 0 11050 0 1 7030
box -12 -8 32 272
use FILL  FILL_4_CLKBUF1_insert44
timestamp 1701859473
transform -1 0 10790 0 1 4430
box -12 -8 32 272
use FILL  FILL_4_CLKBUF1_insert45
timestamp 1701859473
transform 1 0 5710 0 -1 6510
box -12 -8 32 272
use FILL  FILL_4_CLKBUF1_insert46
timestamp 1701859473
transform 1 0 4030 0 1 5990
box -12 -8 32 272
use FILL  FILL_4_CLKBUF1_insert47
timestamp 1701859473
transform -1 0 2150 0 1 7550
box -12 -8 32 272
use FILL  FILL_4_CLKBUF1_insert48
timestamp 1701859473
transform -1 0 10830 0 -1 7030
box -12 -8 32 272
use FILL  FILL_5__1668_
timestamp 1701859473
transform 1 0 6790 0 -1 3390
box -12 -8 32 272
use FILL  FILL_5__1669_
timestamp 1701859473
transform -1 0 6830 0 -1 790
box -12 -8 32 272
use FILL  FILL_5__1670_
timestamp 1701859473
transform 1 0 6610 0 -1 2870
box -12 -8 32 272
use FILL  FILL_5__1671_
timestamp 1701859473
transform -1 0 6410 0 -1 8590
box -12 -8 32 272
use FILL  FILL_5__1672_
timestamp 1701859473
transform 1 0 5970 0 -1 10670
box -12 -8 32 272
use FILL  FILL_5__1673_
timestamp 1701859473
transform 1 0 6370 0 1 8590
box -12 -8 32 272
use FILL  FILL_5__1674_
timestamp 1701859473
transform -1 0 6450 0 -1 9110
box -12 -8 32 272
use FILL  FILL_5__1675_
timestamp 1701859473
transform 1 0 110 0 -1 5470
box -12 -8 32 272
use FILL  FILL_5__1676_
timestamp 1701859473
transform -1 0 350 0 -1 5470
box -12 -8 32 272
use FILL  FILL_5__1677_
timestamp 1701859473
transform -1 0 590 0 1 5470
box -12 -8 32 272
use FILL  FILL_5__1678_
timestamp 1701859473
transform 1 0 110 0 -1 10670
box -12 -8 32 272
use FILL  FILL_5__1679_
timestamp 1701859473
transform -1 0 330 0 -1 11190
box -12 -8 32 272
use FILL  FILL_5__1680_
timestamp 1701859473
transform 1 0 310 0 -1 10670
box -12 -8 32 272
use FILL  FILL_5__1681_
timestamp 1701859473
transform -1 0 130 0 -1 7030
box -12 -8 32 272
use FILL  FILL_5__1682_
timestamp 1701859473
transform -1 0 130 0 1 7030
box -12 -8 32 272
use FILL  FILL_5__1683_
timestamp 1701859473
transform 1 0 110 0 1 6510
box -12 -8 32 272
use FILL  FILL_5__1684_
timestamp 1701859473
transform 1 0 990 0 -1 11190
box -12 -8 32 272
use FILL  FILL_5__1685_
timestamp 1701859473
transform -1 0 1250 0 -1 11190
box -12 -8 32 272
use FILL  FILL_5__1686_
timestamp 1701859473
transform -1 0 1050 0 1 10670
box -12 -8 32 272
use FILL  FILL_5__1687_
timestamp 1701859473
transform 1 0 1470 0 -1 11190
box -12 -8 32 272
use FILL  FILL_5__1688_
timestamp 1701859473
transform -1 0 1730 0 -1 11190
box -12 -8 32 272
use FILL  FILL_5__1689_
timestamp 1701859473
transform -1 0 1990 0 1 10150
box -12 -8 32 272
use FILL  FILL_5__1690_
timestamp 1701859473
transform 1 0 2150 0 1 9110
box -12 -8 32 272
use FILL  FILL_5__1691_
timestamp 1701859473
transform -1 0 2170 0 -1 9110
box -12 -8 32 272
use FILL  FILL_5__1692_
timestamp 1701859473
transform 1 0 110 0 1 790
box -12 -8 32 272
use FILL  FILL_5__1693_
timestamp 1701859473
transform 1 0 110 0 -1 1310
box -12 -8 32 272
use FILL  FILL_5__1694_
timestamp 1701859473
transform 1 0 530 0 -1 270
box -12 -8 32 272
use FILL  FILL_5__1695_
timestamp 1701859473
transform -1 0 750 0 -1 270
box -12 -8 32 272
use FILL  FILL_5__1696_
timestamp 1701859473
transform 1 0 1170 0 1 2870
box -12 -8 32 272
use FILL  FILL_5__1697_
timestamp 1701859473
transform -1 0 2830 0 -1 2870
box -12 -8 32 272
use FILL  FILL_5__1698_
timestamp 1701859473
transform -1 0 1930 0 1 3390
box -12 -8 32 272
use FILL  FILL_5__1699_
timestamp 1701859473
transform 1 0 3850 0 1 3390
box -12 -8 32 272
use FILL  FILL_5__1700_
timestamp 1701859473
transform -1 0 2650 0 -1 3910
box -12 -8 32 272
use FILL  FILL_5__1701_
timestamp 1701859473
transform -1 0 1190 0 1 270
box -12 -8 32 272
use FILL  FILL_5__1702_
timestamp 1701859473
transform 1 0 950 0 1 270
box -12 -8 32 272
use FILL  FILL_5__1703_
timestamp 1701859473
transform -1 0 1430 0 1 1830
box -12 -8 32 272
use FILL  FILL_5__1704_
timestamp 1701859473
transform -1 0 9190 0 1 2870
box -12 -8 32 272
use FILL  FILL_5__1705_
timestamp 1701859473
transform 1 0 9810 0 -1 790
box -12 -8 32 272
use FILL  FILL_5__1706_
timestamp 1701859473
transform -1 0 8030 0 -1 4950
box -12 -8 32 272
use FILL  FILL_5__1707_
timestamp 1701859473
transform 1 0 8470 0 -1 4950
box -12 -8 32 272
use FILL  FILL_5__1708_
timestamp 1701859473
transform 1 0 5090 0 -1 5990
box -12 -8 32 272
use FILL  FILL_5__1709_
timestamp 1701859473
transform -1 0 11190 0 1 5990
box -12 -8 32 272
use FILL  FILL_5__1710_
timestamp 1701859473
transform 1 0 5470 0 -1 5470
box -12 -8 32 272
use FILL  FILL_5__1711_
timestamp 1701859473
transform -1 0 5310 0 -1 5990
box -12 -8 32 272
use FILL  FILL_5__1712_
timestamp 1701859473
transform -1 0 5130 0 1 5470
box -12 -8 32 272
use FILL  FILL_5__1713_
timestamp 1701859473
transform 1 0 7990 0 1 4430
box -12 -8 32 272
use FILL  FILL_5__1714_
timestamp 1701859473
transform 1 0 7790 0 1 4950
box -12 -8 32 272
use FILL  FILL_5__1715_
timestamp 1701859473
transform -1 0 8030 0 1 4950
box -12 -8 32 272
use FILL  FILL_5__1716_
timestamp 1701859473
transform -1 0 8250 0 1 4430
box -12 -8 32 272
use FILL  FILL_5__1717_
timestamp 1701859473
transform -1 0 8030 0 1 1310
box -12 -8 32 272
use FILL  FILL_5__1718_
timestamp 1701859473
transform -1 0 5970 0 1 5990
box -12 -8 32 272
use FILL  FILL_5__1719_
timestamp 1701859473
transform -1 0 6830 0 -1 5990
box -12 -8 32 272
use FILL  FILL_5__1720_
timestamp 1701859473
transform -1 0 6810 0 1 5470
box -12 -8 32 272
use FILL  FILL_5__1721_
timestamp 1701859473
transform -1 0 7050 0 1 5470
box -12 -8 32 272
use FILL  FILL_5__1722_
timestamp 1701859473
transform -1 0 7750 0 1 4430
box -12 -8 32 272
use FILL  FILL_5__1723_
timestamp 1701859473
transform 1 0 7970 0 1 1830
box -12 -8 32 272
use FILL  FILL_5__1724_
timestamp 1701859473
transform -1 0 8010 0 -1 1310
box -12 -8 32 272
use FILL  FILL_5__1725_
timestamp 1701859473
transform 1 0 6610 0 1 5990
box -12 -8 32 272
use FILL  FILL_5__1726_
timestamp 1701859473
transform 1 0 6810 0 1 5990
box -12 -8 32 272
use FILL  FILL_5__1727_
timestamp 1701859473
transform -1 0 7050 0 1 5990
box -12 -8 32 272
use FILL  FILL_5__1728_
timestamp 1701859473
transform 1 0 7750 0 1 5990
box -12 -8 32 272
use FILL  FILL_5__1729_
timestamp 1701859473
transform -1 0 7690 0 -1 5990
box -12 -8 32 272
use FILL  FILL_5__1730_
timestamp 1701859473
transform -1 0 8170 0 1 3390
box -12 -8 32 272
use FILL  FILL_5__1731_
timestamp 1701859473
transform -1 0 8030 0 -1 270
box -12 -8 32 272
use FILL  FILL_5__1732_
timestamp 1701859473
transform -1 0 7990 0 1 5470
box -12 -8 32 272
use FILL  FILL_5__1733_
timestamp 1701859473
transform -1 0 8210 0 1 5470
box -12 -8 32 272
use FILL  FILL_5__1734_
timestamp 1701859473
transform 1 0 8170 0 -1 5470
box -12 -8 32 272
use FILL  FILL_5__1735_
timestamp 1701859473
transform 1 0 8630 0 -1 5470
box -12 -8 32 272
use FILL  FILL_5__1736_
timestamp 1701859473
transform 1 0 8470 0 1 4950
box -12 -8 32 272
use FILL  FILL_5__1737_
timestamp 1701859473
transform -1 0 8550 0 -1 3910
box -12 -8 32 272
use FILL  FILL_5__1738_
timestamp 1701859473
transform 1 0 8950 0 1 790
box -12 -8 32 272
use FILL  FILL_5__1739_
timestamp 1701859473
transform -1 0 9170 0 -1 790
box -12 -8 32 272
use FILL  FILL_5__1740_
timestamp 1701859473
transform 1 0 6530 0 1 270
box -12 -8 32 272
use FILL  FILL_5__1741_
timestamp 1701859473
transform 1 0 6430 0 1 790
box -12 -8 32 272
use FILL  FILL_5__1742_
timestamp 1701859473
transform -1 0 6370 0 -1 790
box -12 -8 32 272
use FILL  FILL_5__1743_
timestamp 1701859473
transform -1 0 2370 0 -1 3390
box -12 -8 32 272
use FILL  FILL_5__1744_
timestamp 1701859473
transform 1 0 350 0 -1 4950
box -12 -8 32 272
use FILL  FILL_5__1745_
timestamp 1701859473
transform 1 0 2170 0 -1 3910
box -12 -8 32 272
use FILL  FILL_5__1746_
timestamp 1701859473
transform -1 0 5190 0 -1 3390
box -12 -8 32 272
use FILL  FILL_5__1747_
timestamp 1701859473
transform -1 0 350 0 -1 270
box -12 -8 32 272
use FILL  FILL_5__1748_
timestamp 1701859473
transform -1 0 550 0 1 270
box -12 -8 32 272
use FILL  FILL_5__1749_
timestamp 1701859473
transform -1 0 990 0 1 1310
box -12 -8 32 272
use FILL  FILL_5__1750_
timestamp 1701859473
transform -1 0 1210 0 1 1310
box -12 -8 32 272
use FILL  FILL_5__1751_
timestamp 1701859473
transform -1 0 4570 0 -1 2870
box -12 -8 32 272
use FILL  FILL_5__1752_
timestamp 1701859473
transform 1 0 4770 0 -1 2870
box -12 -8 32 272
use FILL  FILL_5__1753_
timestamp 1701859473
transform -1 0 4390 0 1 790
box -12 -8 32 272
use FILL  FILL_5__1754_
timestamp 1701859473
transform 1 0 330 0 -1 790
box -12 -8 32 272
use FILL  FILL_5__1755_
timestamp 1701859473
transform -1 0 550 0 -1 790
box -12 -8 32 272
use FILL  FILL_5__1756_
timestamp 1701859473
transform -1 0 130 0 -1 270
box -12 -8 32 272
use FILL  FILL_5__1757_
timestamp 1701859473
transform 1 0 730 0 -1 790
box -12 -8 32 272
use FILL  FILL_5__1758_
timestamp 1701859473
transform 1 0 110 0 1 2350
box -12 -8 32 272
use FILL  FILL_5__1759_
timestamp 1701859473
transform -1 0 2610 0 -1 2870
box -12 -8 32 272
use FILL  FILL_5__1760_
timestamp 1701859473
transform 1 0 2990 0 -1 2870
box -12 -8 32 272
use FILL  FILL_5__1761_
timestamp 1701859473
transform -1 0 3310 0 -1 3390
box -12 -8 32 272
use FILL  FILL_5__1762_
timestamp 1701859473
transform -1 0 130 0 1 270
box -12 -8 32 272
use FILL  FILL_5__1763_
timestamp 1701859473
transform 1 0 110 0 -1 790
box -12 -8 32 272
use FILL  FILL_5__1764_
timestamp 1701859473
transform 1 0 550 0 1 1310
box -12 -8 32 272
use FILL  FILL_5__1765_
timestamp 1701859473
transform 1 0 1410 0 1 1310
box -12 -8 32 272
use FILL  FILL_5__1766_
timestamp 1701859473
transform -1 0 3210 0 -1 1830
box -12 -8 32 272
use FILL  FILL_5__1767_
timestamp 1701859473
transform 1 0 1510 0 -1 4430
box -12 -8 32 272
use FILL  FILL_5__1768_
timestamp 1701859473
transform 1 0 330 0 -1 1310
box -12 -8 32 272
use FILL  FILL_5__1769_
timestamp 1701859473
transform -1 0 550 0 1 1830
box -12 -8 32 272
use FILL  FILL_5__1770_
timestamp 1701859473
transform 1 0 2150 0 -1 3390
box -12 -8 32 272
use FILL  FILL_5__1771_
timestamp 1701859473
transform -1 0 2410 0 -1 3910
box -12 -8 32 272
use FILL  FILL_5__1772_
timestamp 1701859473
transform -1 0 3070 0 -1 3910
box -12 -8 32 272
use FILL  FILL_5__1773_
timestamp 1701859473
transform 1 0 3970 0 1 2870
box -12 -8 32 272
use FILL  FILL_5__1774_
timestamp 1701859473
transform -1 0 5350 0 -1 2350
box -12 -8 32 272
use FILL  FILL_5__1775_
timestamp 1701859473
transform 1 0 310 0 1 790
box -12 -8 32 272
use FILL  FILL_5__1776_
timestamp 1701859473
transform -1 0 350 0 1 1310
box -12 -8 32 272
use FILL  FILL_5__1777_
timestamp 1701859473
transform 1 0 770 0 -1 1830
box -12 -8 32 272
use FILL  FILL_5__1778_
timestamp 1701859473
transform -1 0 4490 0 1 5470
box -12 -8 32 272
use FILL  FILL_5__1779_
timestamp 1701859473
transform -1 0 6130 0 -1 5470
box -12 -8 32 272
use FILL  FILL_5__1780_
timestamp 1701859473
transform 1 0 4850 0 1 2870
box -12 -8 32 272
use FILL  FILL_5__1781_
timestamp 1701859473
transform 1 0 4430 0 1 2870
box -12 -8 32 272
use FILL  FILL_5__1782_
timestamp 1701859473
transform -1 0 130 0 1 1310
box -12 -8 32 272
use FILL  FILL_5__1783_
timestamp 1701859473
transform -1 0 1410 0 1 2870
box -12 -8 32 272
use FILL  FILL_5__1784_
timestamp 1701859473
transform -1 0 5110 0 1 2870
box -12 -8 32 272
use FILL  FILL_5__1785_
timestamp 1701859473
transform 1 0 5030 0 -1 2870
box -12 -8 32 272
use FILL  FILL_5__1786_
timestamp 1701859473
transform -1 0 5110 0 -1 2350
box -12 -8 32 272
use FILL  FILL_5__1787_
timestamp 1701859473
transform 1 0 5090 0 1 2350
box -12 -8 32 272
use FILL  FILL_5__1788_
timestamp 1701859473
transform -1 0 4890 0 -1 2350
box -12 -8 32 272
use FILL  FILL_5__1789_
timestamp 1701859473
transform 1 0 110 0 1 1830
box -12 -8 32 272
use FILL  FILL_5__1790_
timestamp 1701859473
transform -1 0 350 0 -1 2350
box -12 -8 32 272
use FILL  FILL_5__1791_
timestamp 1701859473
transform -1 0 2150 0 -1 2350
box -12 -8 32 272
use FILL  FILL_5__1792_
timestamp 1701859473
transform -1 0 3530 0 -1 2350
box -12 -8 32 272
use FILL  FILL_5__1793_
timestamp 1701859473
transform -1 0 4630 0 1 1830
box -12 -8 32 272
use FILL  FILL_5__1794_
timestamp 1701859473
transform 1 0 950 0 1 1830
box -12 -8 32 272
use FILL  FILL_5__1795_
timestamp 1701859473
transform -1 0 2210 0 1 2350
box -12 -8 32 272
use FILL  FILL_5__1796_
timestamp 1701859473
transform -1 0 1830 0 -1 1830
box -12 -8 32 272
use FILL  FILL_5__1797_
timestamp 1701859473
transform 1 0 2050 0 -1 1830
box -12 -8 32 272
use FILL  FILL_5__1798_
timestamp 1701859473
transform 1 0 970 0 -1 1310
box -12 -8 32 272
use FILL  FILL_5__1799_
timestamp 1701859473
transform 1 0 3790 0 1 3910
box -12 -8 32 272
use FILL  FILL_5__1800_
timestamp 1701859473
transform 1 0 3470 0 1 1830
box -12 -8 32 272
use FILL  FILL_5__1801_
timestamp 1701859473
transform -1 0 1210 0 1 1830
box -12 -8 32 272
use FILL  FILL_5__1802_
timestamp 1701859473
transform -1 0 3750 0 1 2350
box -12 -8 32 272
use FILL  FILL_5__1803_
timestamp 1701859473
transform -1 0 3970 0 1 2350
box -12 -8 32 272
use FILL  FILL_5__1804_
timestamp 1701859473
transform -1 0 4210 0 1 2350
box -12 -8 32 272
use FILL  FILL_5__1805_
timestamp 1701859473
transform 1 0 5510 0 1 2350
box -12 -8 32 272
use FILL  FILL_5__1806_
timestamp 1701859473
transform -1 0 4910 0 1 2350
box -12 -8 32 272
use FILL  FILL_5__1807_
timestamp 1701859473
transform -1 0 5310 0 1 2350
box -12 -8 32 272
use FILL  FILL_5__1808_
timestamp 1701859473
transform 1 0 4830 0 1 1830
box -12 -8 32 272
use FILL  FILL_5__1809_
timestamp 1701859473
transform -1 0 7190 0 -1 270
box -12 -8 32 272
use FILL  FILL_5__1810_
timestamp 1701859473
transform -1 0 7170 0 1 1310
box -12 -8 32 272
use FILL  FILL_5__1811_
timestamp 1701859473
transform 1 0 7510 0 -1 1830
box -12 -8 32 272
use FILL  FILL_5__1812_
timestamp 1701859473
transform -1 0 7590 0 -1 1310
box -12 -8 32 272
use FILL  FILL_5__1813_
timestamp 1701859473
transform 1 0 9170 0 1 790
box -12 -8 32 272
use FILL  FILL_5__1814_
timestamp 1701859473
transform -1 0 8210 0 -1 1830
box -12 -8 32 272
use FILL  FILL_5__1815_
timestamp 1701859473
transform 1 0 8410 0 1 2350
box -12 -8 32 272
use FILL  FILL_5__1816_
timestamp 1701859473
transform -1 0 9690 0 -1 2350
box -12 -8 32 272
use FILL  FILL_5__1817_
timestamp 1701859473
transform -1 0 9410 0 1 1310
box -12 -8 32 272
use FILL  FILL_5__1818_
timestamp 1701859473
transform -1 0 9610 0 1 270
box -12 -8 32 272
use FILL  FILL_5__1819_
timestamp 1701859473
transform -1 0 8430 0 -1 1830
box -12 -8 32 272
use FILL  FILL_5__1820_
timestamp 1701859473
transform -1 0 8510 0 1 1310
box -12 -8 32 272
use FILL  FILL_5__1821_
timestamp 1701859473
transform -1 0 4950 0 1 1310
box -12 -8 32 272
use FILL  FILL_5__1822_
timestamp 1701859473
transform -1 0 4750 0 -1 790
box -12 -8 32 272
use FILL  FILL_5__1823_
timestamp 1701859473
transform -1 0 4290 0 -1 790
box -12 -8 32 272
use FILL  FILL_5__1824_
timestamp 1701859473
transform 1 0 4670 0 1 2350
box -12 -8 32 272
use FILL  FILL_5__1825_
timestamp 1701859473
transform 1 0 5730 0 1 1830
box -12 -8 32 272
use FILL  FILL_5__1826_
timestamp 1701859473
transform 1 0 8230 0 -1 270
box -12 -8 32 272
use FILL  FILL_5__1827_
timestamp 1701859473
transform 1 0 9370 0 -1 790
box -12 -8 32 272
use FILL  FILL_5__1828_
timestamp 1701859473
transform 1 0 8530 0 1 270
box -12 -8 32 272
use FILL  FILL_5__1829_
timestamp 1701859473
transform 1 0 5830 0 1 270
box -12 -8 32 272
use FILL  FILL_5__1830_
timestamp 1701859473
transform 1 0 3270 0 1 4430
box -12 -8 32 272
use FILL  FILL_5__1831_
timestamp 1701859473
transform -1 0 8050 0 -1 790
box -12 -8 32 272
use FILL  FILL_5__1832_
timestamp 1701859473
transform 1 0 6550 0 -1 790
box -12 -8 32 272
use FILL  FILL_5__1833_
timestamp 1701859473
transform -1 0 750 0 1 270
box -12 -8 32 272
use FILL  FILL_5__1834_
timestamp 1701859473
transform 1 0 1190 0 -1 1310
box -12 -8 32 272
use FILL  FILL_5__1835_
timestamp 1701859473
transform -1 0 2570 0 -1 1310
box -12 -8 32 272
use FILL  FILL_5__1836_
timestamp 1701859473
transform 1 0 1130 0 1 790
box -12 -8 32 272
use FILL  FILL_5__1837_
timestamp 1701859473
transform -1 0 2530 0 1 790
box -12 -8 32 272
use FILL  FILL_5__1838_
timestamp 1701859473
transform 1 0 2270 0 1 790
box -12 -8 32 272
use FILL  FILL_5__1839_
timestamp 1701859473
transform -1 0 330 0 1 270
box -12 -8 32 272
use FILL  FILL_5__1840_
timestamp 1701859473
transform -1 0 970 0 1 2870
box -12 -8 32 272
use FILL  FILL_5__1841_
timestamp 1701859473
transform 1 0 3750 0 1 2870
box -12 -8 32 272
use FILL  FILL_5__1842_
timestamp 1701859473
transform -1 0 3010 0 -1 1830
box -12 -8 32 272
use FILL  FILL_5__1843_
timestamp 1701859473
transform -1 0 3970 0 -1 2350
box -12 -8 32 272
use FILL  FILL_5__1844_
timestamp 1701859473
transform 1 0 3870 0 -1 2870
box -12 -8 32 272
use FILL  FILL_5__1845_
timestamp 1701859473
transform -1 0 1810 0 -1 4950
box -12 -8 32 272
use FILL  FILL_5__1846_
timestamp 1701859473
transform 1 0 4170 0 1 4430
box -12 -8 32 272
use FILL  FILL_5__1847_
timestamp 1701859473
transform 1 0 3490 0 1 4430
box -12 -8 32 272
use FILL  FILL_5__1848_
timestamp 1701859473
transform 1 0 3930 0 1 4430
box -12 -8 32 272
use FILL  FILL_5__1849_
timestamp 1701859473
transform -1 0 4130 0 -1 2870
box -12 -8 32 272
use FILL  FILL_5__1850_
timestamp 1701859473
transform -1 0 950 0 1 790
box -12 -8 32 272
use FILL  FILL_5__1851_
timestamp 1701859473
transform 1 0 1610 0 -1 1830
box -12 -8 32 272
use FILL  FILL_5__1852_
timestamp 1701859473
transform -1 0 2430 0 1 2350
box -12 -8 32 272
use FILL  FILL_5__1853_
timestamp 1701859473
transform 1 0 110 0 -1 2350
box -12 -8 32 272
use FILL  FILL_5__1854_
timestamp 1701859473
transform 1 0 2350 0 -1 2350
box -12 -8 32 272
use FILL  FILL_5__1855_
timestamp 1701859473
transform -1 0 2610 0 -1 2350
box -12 -8 32 272
use FILL  FILL_5__1856_
timestamp 1701859473
transform 1 0 1510 0 -1 790
box -12 -8 32 272
use FILL  FILL_5__1857_
timestamp 1701859473
transform -1 0 2710 0 -1 790
box -12 -8 32 272
use FILL  FILL_5__1858_
timestamp 1701859473
transform 1 0 2450 0 -1 790
box -12 -8 32 272
use FILL  FILL_5__1859_
timestamp 1701859473
transform 1 0 2230 0 -1 790
box -12 -8 32 272
use FILL  FILL_5__1860_
timestamp 1701859473
transform -1 0 1770 0 -1 790
box -12 -8 32 272
use FILL  FILL_5__1861_
timestamp 1701859473
transform -1 0 2010 0 -1 790
box -12 -8 32 272
use FILL  FILL_5__1862_
timestamp 1701859473
transform -1 0 2090 0 1 270
box -12 -8 32 272
use FILL  FILL_5__1863_
timestamp 1701859473
transform 1 0 2310 0 1 270
box -12 -8 32 272
use FILL  FILL_5__1864_
timestamp 1701859473
transform 1 0 3550 0 1 270
box -12 -8 32 272
use FILL  FILL_5__1865_
timestamp 1701859473
transform 1 0 7350 0 -1 1310
box -12 -8 32 272
use FILL  FILL_5__1866_
timestamp 1701859473
transform 1 0 3710 0 -1 1310
box -12 -8 32 272
use FILL  FILL_5__1867_
timestamp 1701859473
transform 1 0 1170 0 -1 1830
box -12 -8 32 272
use FILL  FILL_5__1868_
timestamp 1701859473
transform 1 0 1610 0 1 1310
box -12 -8 32 272
use FILL  FILL_5__1869_
timestamp 1701859473
transform 1 0 2030 0 1 1310
box -12 -8 32 272
use FILL  FILL_5__1870_
timestamp 1701859473
transform -1 0 1650 0 -1 1310
box -12 -8 32 272
use FILL  FILL_5__1871_
timestamp 1701859473
transform -1 0 2770 0 -1 1310
box -12 -8 32 272
use FILL  FILL_5__1872_
timestamp 1701859473
transform -1 0 550 0 1 790
box -12 -8 32 272
use FILL  FILL_5__1873_
timestamp 1701859473
transform 1 0 730 0 1 790
box -12 -8 32 272
use FILL  FILL_5__1874_
timestamp 1701859473
transform -1 0 1370 0 1 790
box -12 -8 32 272
use FILL  FILL_5__1875_
timestamp 1701859473
transform 1 0 950 0 -1 790
box -12 -8 32 272
use FILL  FILL_5__1876_
timestamp 1701859473
transform 1 0 1270 0 -1 790
box -12 -8 32 272
use FILL  FILL_5__1877_
timestamp 1701859473
transform 1 0 2210 0 1 4950
box -12 -8 32 272
use FILL  FILL_5__1878_
timestamp 1701859473
transform 1 0 550 0 -1 1310
box -12 -8 32 272
use FILL  FILL_5__1879_
timestamp 1701859473
transform 1 0 770 0 1 1310
box -12 -8 32 272
use FILL  FILL_5__1880_
timestamp 1701859473
transform -1 0 2030 0 -1 4950
box -12 -8 32 272
use FILL  FILL_5__1881_
timestamp 1701859473
transform -1 0 2270 0 -1 4950
box -12 -8 32 272
use FILL  FILL_5__1882_
timestamp 1701859473
transform 1 0 1590 0 -1 3390
box -12 -8 32 272
use FILL  FILL_5__1883_
timestamp 1701859473
transform 1 0 1070 0 -1 3390
box -12 -8 32 272
use FILL  FILL_5__1884_
timestamp 1701859473
transform -1 0 4090 0 1 3390
box -12 -8 32 272
use FILL  FILL_5__1885_
timestamp 1701859473
transform -1 0 3810 0 -1 3390
box -12 -8 32 272
use FILL  FILL_5__1886_
timestamp 1701859473
transform 1 0 3550 0 -1 3390
box -12 -8 32 272
use FILL  FILL_5__1887_
timestamp 1701859473
transform -1 0 3530 0 1 2870
box -12 -8 32 272
use FILL  FILL_5__1888_
timestamp 1701859473
transform -1 0 2570 0 1 270
box -12 -8 32 272
use FILL  FILL_5__1889_
timestamp 1701859473
transform 1 0 1710 0 -1 2870
box -12 -8 32 272
use FILL  FILL_5__1890_
timestamp 1701859473
transform -1 0 350 0 -1 1830
box -12 -8 32 272
use FILL  FILL_5__1891_
timestamp 1701859473
transform 1 0 110 0 -1 1830
box -12 -8 32 272
use FILL  FILL_5__1892_
timestamp 1701859473
transform 1 0 4950 0 -1 3390
box -12 -8 32 272
use FILL  FILL_5__1893_
timestamp 1701859473
transform 1 0 3950 0 1 1830
box -12 -8 32 272
use FILL  FILL_5__1894_
timestamp 1701859473
transform 1 0 4150 0 1 1830
box -12 -8 32 272
use FILL  FILL_5__1895_
timestamp 1701859473
transform -1 0 1890 0 1 1830
box -12 -8 32 272
use FILL  FILL_5__1896_
timestamp 1701859473
transform 1 0 1910 0 -1 2350
box -12 -8 32 272
use FILL  FILL_5__1897_
timestamp 1701859473
transform 1 0 3530 0 1 2350
box -12 -8 32 272
use FILL  FILL_5__1898_
timestamp 1701859473
transform 1 0 3310 0 1 2350
box -12 -8 32 272
use FILL  FILL_5__1899_
timestamp 1701859473
transform -1 0 3290 0 -1 2350
box -12 -8 32 272
use FILL  FILL_5__1900_
timestamp 1701859473
transform -1 0 4130 0 -1 1830
box -12 -8 32 272
use FILL  FILL_5__1901_
timestamp 1701859473
transform -1 0 770 0 1 1830
box -12 -8 32 272
use FILL  FILL_5__1902_
timestamp 1701859473
transform 1 0 5070 0 1 1830
box -12 -8 32 272
use FILL  FILL_5__1903_
timestamp 1701859473
transform 1 0 3390 0 1 1310
box -12 -8 32 272
use FILL  FILL_5__1904_
timestamp 1701859473
transform -1 0 3490 0 -1 1310
box -12 -8 32 272
use FILL  FILL_5__1905_
timestamp 1701859473
transform 1 0 3030 0 1 270
box -12 -8 32 272
use FILL  FILL_5__1906_
timestamp 1701859473
transform 1 0 310 0 1 2350
box -12 -8 32 272
use FILL  FILL_5__1907_
timestamp 1701859473
transform -1 0 3070 0 -1 2350
box -12 -8 32 272
use FILL  FILL_5__1908_
timestamp 1701859473
transform 1 0 6490 0 -1 2350
box -12 -8 32 272
use FILL  FILL_5__1909_
timestamp 1701859473
transform -1 0 6090 0 -1 2350
box -12 -8 32 272
use FILL  FILL_5__1910_
timestamp 1701859473
transform -1 0 5590 0 -1 2350
box -12 -8 32 272
use FILL  FILL_5__1911_
timestamp 1701859473
transform -1 0 750 0 1 2870
box -12 -8 32 272
use FILL  FILL_5__1912_
timestamp 1701859473
transform -1 0 3350 0 1 3910
box -12 -8 32 272
use FILL  FILL_5__1913_
timestamp 1701859473
transform -1 0 1070 0 -1 2870
box -12 -8 32 272
use FILL  FILL_5__1914_
timestamp 1701859473
transform -1 0 1510 0 1 3390
box -12 -8 32 272
use FILL  FILL_5__1915_
timestamp 1701859473
transform 1 0 2590 0 1 3390
box -12 -8 32 272
use FILL  FILL_5__1916_
timestamp 1701859473
transform -1 0 3450 0 1 3390
box -12 -8 32 272
use FILL  FILL_5__1917_
timestamp 1701859473
transform -1 0 4730 0 -1 3390
box -12 -8 32 272
use FILL  FILL_5__1918_
timestamp 1701859473
transform 1 0 1770 0 1 4950
box -12 -8 32 272
use FILL  FILL_5__1919_
timestamp 1701859473
transform -1 0 1290 0 -1 2870
box -12 -8 32 272
use FILL  FILL_5__1920_
timestamp 1701859473
transform -1 0 5070 0 1 4430
box -12 -8 32 272
use FILL  FILL_5__1921_
timestamp 1701859473
transform 1 0 4830 0 1 4430
box -12 -8 32 272
use FILL  FILL_5__1922_
timestamp 1701859473
transform -1 0 4630 0 1 4430
box -12 -8 32 272
use FILL  FILL_5__1923_
timestamp 1701859473
transform 1 0 4490 0 -1 3390
box -12 -8 32 272
use FILL  FILL_5__1924_
timestamp 1701859473
transform 1 0 1990 0 1 4950
box -12 -8 32 272
use FILL  FILL_5__1925_
timestamp 1701859473
transform 1 0 6130 0 -1 4430
box -12 -8 32 272
use FILL  FILL_5__1926_
timestamp 1701859473
transform 1 0 750 0 -1 1310
box -12 -8 32 272
use FILL  FILL_5__1927_
timestamp 1701859473
transform 1 0 2990 0 -1 1310
box -12 -8 32 272
use FILL  FILL_5__1928_
timestamp 1701859473
transform -1 0 3250 0 -1 1310
box -12 -8 32 272
use FILL  FILL_5__1929_
timestamp 1701859473
transform 1 0 3430 0 1 790
box -12 -8 32 272
use FILL  FILL_5__1930_
timestamp 1701859473
transform 1 0 3250 0 1 270
box -12 -8 32 272
use FILL  FILL_5__1931_
timestamp 1701859473
transform 1 0 3850 0 1 270
box -12 -8 32 272
use FILL  FILL_5__1932_
timestamp 1701859473
transform -1 0 4090 0 1 270
box -12 -8 32 272
use FILL  FILL_5__1933_
timestamp 1701859473
transform -1 0 1890 0 1 270
box -12 -8 32 272
use FILL  FILL_5__1934_
timestamp 1701859473
transform -1 0 5510 0 1 790
box -12 -8 32 272
use FILL  FILL_5__1935_
timestamp 1701859473
transform 1 0 5630 0 -1 270
box -12 -8 32 272
use FILL  FILL_5__1936_
timestamp 1701859473
transform -1 0 8390 0 1 3390
box -12 -8 32 272
use FILL  FILL_5__1937_
timestamp 1701859473
transform -1 0 7610 0 -1 270
box -12 -8 32 272
use FILL  FILL_5__1938_
timestamp 1701859473
transform -1 0 7810 0 -1 270
box -12 -8 32 272
use FILL  FILL_5__1939_
timestamp 1701859473
transform -1 0 6730 0 -1 270
box -12 -8 32 272
use FILL  FILL_5__1940_
timestamp 1701859473
transform -1 0 5850 0 -1 270
box -12 -8 32 272
use FILL  FILL_5__1941_
timestamp 1701859473
transform 1 0 5870 0 -1 790
box -12 -8 32 272
use FILL  FILL_5__1942_
timestamp 1701859473
transform 1 0 4850 0 -1 1310
box -12 -8 32 272
use FILL  FILL_5__1943_
timestamp 1701859473
transform 1 0 8110 0 1 270
box -12 -8 32 272
use FILL  FILL_5__1944_
timestamp 1701859473
transform -1 0 8350 0 1 270
box -12 -8 32 272
use FILL  FILL_5__1945_
timestamp 1701859473
transform 1 0 7890 0 1 270
box -12 -8 32 272
use FILL  FILL_5__1946_
timestamp 1701859473
transform -1 0 6090 0 1 270
box -12 -8 32 272
use FILL  FILL_5__1947_
timestamp 1701859473
transform -1 0 6110 0 -1 790
box -12 -8 32 272
use FILL  FILL_5__1948_
timestamp 1701859473
transform 1 0 5390 0 -1 790
box -12 -8 32 272
use FILL  FILL_5__1949_
timestamp 1701859473
transform 1 0 4630 0 -1 1310
box -12 -8 32 272
use FILL  FILL_5__1950_
timestamp 1701859473
transform -1 0 8270 0 -1 790
box -12 -8 32 272
use FILL  FILL_5__1951_
timestamp 1701859473
transform 1 0 550 0 -1 2350
box -12 -8 32 272
use FILL  FILL_5__1952_
timestamp 1701859473
transform -1 0 5730 0 1 2350
box -12 -8 32 272
use FILL  FILL_5__1953_
timestamp 1701859473
transform 1 0 5830 0 -1 2350
box -12 -8 32 272
use FILL  FILL_5__1954_
timestamp 1701859473
transform 1 0 8210 0 -1 1310
box -12 -8 32 272
use FILL  FILL_5__1955_
timestamp 1701859473
transform -1 0 8750 0 1 1310
box -12 -8 32 272
use FILL  FILL_5__1956_
timestamp 1701859473
transform -1 0 6290 0 -1 1310
box -12 -8 32 272
use FILL  FILL_5__1957_
timestamp 1701859473
transform -1 0 6050 0 -1 1310
box -12 -8 32 272
use FILL  FILL_5__1958_
timestamp 1701859473
transform 1 0 5310 0 -1 1310
box -12 -8 32 272
use FILL  FILL_5__1959_
timestamp 1701859473
transform 1 0 5750 0 -1 2870
box -12 -8 32 272
use FILL  FILL_5__1960_
timestamp 1701859473
transform -1 0 6190 0 -1 2870
box -12 -8 32 272
use FILL  FILL_5__1961_
timestamp 1701859473
transform -1 0 4450 0 1 2350
box -12 -8 32 272
use FILL  FILL_5__1962_
timestamp 1701859473
transform 1 0 5910 0 1 2350
box -12 -8 32 272
use FILL  FILL_5__1963_
timestamp 1701859473
transform 1 0 5370 0 1 1310
box -12 -8 32 272
use FILL  FILL_5__1964_
timestamp 1701859473
transform 1 0 9190 0 1 1310
box -12 -8 32 272
use FILL  FILL_5__1965_
timestamp 1701859473
transform 1 0 7590 0 1 790
box -12 -8 32 272
use FILL  FILL_5__1966_
timestamp 1701859473
transform -1 0 7710 0 1 270
box -12 -8 32 272
use FILL  FILL_5__1967_
timestamp 1701859473
transform -1 0 6770 0 1 270
box -12 -8 32 272
use FILL  FILL_5__1968_
timestamp 1701859473
transform 1 0 5550 0 -1 1310
box -12 -8 32 272
use FILL  FILL_5__1969_
timestamp 1701859473
transform 1 0 5750 0 1 2870
box -12 -8 32 272
use FILL  FILL_5__1970_
timestamp 1701859473
transform 1 0 5390 0 -1 3390
box -12 -8 32 272
use FILL  FILL_5__1971_
timestamp 1701859473
transform 1 0 5830 0 1 3910
box -12 -8 32 272
use FILL  FILL_5__1972_
timestamp 1701859473
transform 1 0 5770 0 1 4950
box -12 -8 32 272
use FILL  FILL_5__1973_
timestamp 1701859473
transform -1 0 6110 0 -1 3910
box -12 -8 32 272
use FILL  FILL_5__1974_
timestamp 1701859473
transform 1 0 6290 0 -1 3910
box -12 -8 32 272
use FILL  FILL_5__1975_
timestamp 1701859473
transform -1 0 6090 0 1 3910
box -12 -8 32 272
use FILL  FILL_5__1976_
timestamp 1701859473
transform -1 0 6550 0 -1 3910
box -12 -8 32 272
use FILL  FILL_5__1977_
timestamp 1701859473
transform 1 0 6870 0 1 2870
box -12 -8 32 272
use FILL  FILL_5__1978_
timestamp 1701859473
transform -1 0 6410 0 -1 2870
box -12 -8 32 272
use FILL  FILL_5__1979_
timestamp 1701859473
transform 1 0 6450 0 1 2870
box -12 -8 32 272
use FILL  FILL_5__1980_
timestamp 1701859473
transform 1 0 6650 0 1 2870
box -12 -8 32 272
use FILL  FILL_5__1981_
timestamp 1701859473
transform 1 0 6230 0 1 2870
box -12 -8 32 272
use FILL  FILL_5__1982_
timestamp 1701859473
transform -1 0 5690 0 -1 1830
box -12 -8 32 272
use FILL  FILL_5__1983_
timestamp 1701859473
transform -1 0 4790 0 -1 270
box -12 -8 32 272
use FILL  FILL_5__1984_
timestamp 1701859473
transform -1 0 6490 0 -1 1310
box -12 -8 32 272
use FILL  FILL_5__1985_
timestamp 1701859473
transform 1 0 5050 0 -1 1310
box -12 -8 32 272
use FILL  FILL_5__1986_
timestamp 1701859473
transform 1 0 8250 0 1 790
box -12 -8 32 272
use FILL  FILL_5__1987_
timestamp 1701859473
transform 1 0 6930 0 1 1310
box -12 -8 32 272
use FILL  FILL_5__1988_
timestamp 1701859473
transform -1 0 7390 0 1 1310
box -12 -8 32 272
use FILL  FILL_5__1989_
timestamp 1701859473
transform 1 0 2750 0 -1 5470
box -12 -8 32 272
use FILL  FILL_5__1990_
timestamp 1701859473
transform 1 0 2070 0 1 1830
box -12 -8 32 272
use FILL  FILL_5__1991_
timestamp 1701859473
transform -1 0 2790 0 1 1830
box -12 -8 32 272
use FILL  FILL_5__1992_
timestamp 1701859473
transform -1 0 4190 0 -1 2350
box -12 -8 32 272
use FILL  FILL_5__1993_
timestamp 1701859473
transform -1 0 4430 0 -1 2350
box -12 -8 32 272
use FILL  FILL_5__1994_
timestamp 1701859473
transform 1 0 2530 0 1 1830
box -12 -8 32 272
use FILL  FILL_5__1995_
timestamp 1701859473
transform 1 0 3010 0 1 1830
box -12 -8 32 272
use FILL  FILL_5__1996_
timestamp 1701859473
transform -1 0 6690 0 1 790
box -12 -8 32 272
use FILL  FILL_5__1997_
timestamp 1701859473
transform -1 0 5030 0 1 790
box -12 -8 32 272
use FILL  FILL_5__1998_
timestamp 1701859473
transform 1 0 4290 0 1 270
box -12 -8 32 272
use FILL  FILL_5__1999_
timestamp 1701859473
transform -1 0 3890 0 -1 270
box -12 -8 32 272
use FILL  FILL_5__2000_
timestamp 1701859473
transform -1 0 4570 0 -1 270
box -12 -8 32 272
use FILL  FILL_5__2001_
timestamp 1701859473
transform -1 0 5950 0 -1 2870
box -12 -8 32 272
use FILL  FILL_5__2002_
timestamp 1701859473
transform -1 0 1890 0 1 2870
box -12 -8 32 272
use FILL  FILL_5__2003_
timestamp 1701859473
transform 1 0 1390 0 -1 3390
box -12 -8 32 272
use FILL  FILL_5__2004_
timestamp 1701859473
transform 1 0 2810 0 -1 3390
box -12 -8 32 272
use FILL  FILL_5__2005_
timestamp 1701859473
transform -1 0 3090 0 1 2870
box -12 -8 32 272
use FILL  FILL_5__2006_
timestamp 1701859473
transform 1 0 2830 0 1 2870
box -12 -8 32 272
use FILL  FILL_5__2007_
timestamp 1701859473
transform 1 0 6850 0 -1 2870
box -12 -8 32 272
use FILL  FILL_5__2008_
timestamp 1701859473
transform 1 0 530 0 -1 1830
box -12 -8 32 272
use FILL  FILL_5__2009_
timestamp 1701859473
transform -1 0 4050 0 -1 3390
box -12 -8 32 272
use FILL  FILL_5__2010_
timestamp 1701859473
transform -1 0 4350 0 -1 2870
box -12 -8 32 272
use FILL  FILL_5__2011_
timestamp 1701859473
transform -1 0 2090 0 1 790
box -12 -8 32 272
use FILL  FILL_5__2012_
timestamp 1701859473
transform 1 0 1590 0 1 790
box -12 -8 32 272
use FILL  FILL_5__2013_
timestamp 1701859473
transform -1 0 1850 0 1 790
box -12 -8 32 272
use FILL  FILL_5__2014_
timestamp 1701859473
transform 1 0 4510 0 1 1310
box -12 -8 32 272
use FILL  FILL_5__2015_
timestamp 1701859473
transform 1 0 3230 0 1 1830
box -12 -8 32 272
use FILL  FILL_5__2016_
timestamp 1701859473
transform -1 0 3730 0 1 1830
box -12 -8 32 272
use FILL  FILL_5__2017_
timestamp 1701859473
transform -1 0 5250 0 -1 1830
box -12 -8 32 272
use FILL  FILL_5__2018_
timestamp 1701859473
transform 1 0 5010 0 -1 1830
box -12 -8 32 272
use FILL  FILL_5__2019_
timestamp 1701859473
transform -1 0 5530 0 -1 2870
box -12 -8 32 272
use FILL  FILL_5__2020_
timestamp 1701859473
transform -1 0 5290 0 -1 2870
box -12 -8 32 272
use FILL  FILL_5__2021_
timestamp 1701859473
transform -1 0 6930 0 -1 1310
box -12 -8 32 272
use FILL  FILL_5__2022_
timestamp 1701859473
transform -1 0 7170 0 1 790
box -12 -8 32 272
use FILL  FILL_5__2023_
timestamp 1701859473
transform 1 0 8210 0 1 1830
box -12 -8 32 272
use FILL  FILL_5__2024_
timestamp 1701859473
transform -1 0 8430 0 1 1830
box -12 -8 32 272
use FILL  FILL_5__2025_
timestamp 1701859473
transform 1 0 9590 0 -1 790
box -12 -8 32 272
use FILL  FILL_5__2026_
timestamp 1701859473
transform -1 0 8730 0 1 790
box -12 -8 32 272
use FILL  FILL_5__2027_
timestamp 1701859473
transform -1 0 6930 0 1 790
box -12 -8 32 272
use FILL  FILL_5__2028_
timestamp 1701859473
transform 1 0 7030 0 -1 790
box -12 -8 32 272
use FILL  FILL_5__2029_
timestamp 1701859473
transform 1 0 7470 0 1 270
box -12 -8 32 272
use FILL  FILL_5__2030_
timestamp 1701859473
transform -1 0 7150 0 -1 1310
box -12 -8 32 272
use FILL  FILL_5__2031_
timestamp 1701859473
transform 1 0 7470 0 -1 790
box -12 -8 32 272
use FILL  FILL_5__2032_
timestamp 1701859473
transform -1 0 8770 0 1 270
box -12 -8 32 272
use FILL  FILL_5__2033_
timestamp 1701859473
transform 1 0 8250 0 1 1310
box -12 -8 32 272
use FILL  FILL_5__2034_
timestamp 1701859473
transform -1 0 8930 0 -1 1310
box -12 -8 32 272
use FILL  FILL_5__2035_
timestamp 1701859473
transform -1 0 8510 0 1 790
box -12 -8 32 272
use FILL  FILL_5__2036_
timestamp 1701859473
transform -1 0 8670 0 -1 1830
box -12 -8 32 272
use FILL  FILL_5__2037_
timestamp 1701859473
transform -1 0 8730 0 -1 790
box -12 -8 32 272
use FILL  FILL_5__2038_
timestamp 1701859473
transform 1 0 8030 0 1 790
box -12 -8 32 272
use FILL  FILL_5__2039_
timestamp 1701859473
transform 1 0 7810 0 1 790
box -12 -8 32 272
use FILL  FILL_5__2040_
timestamp 1701859473
transform -1 0 7730 0 -1 790
box -12 -8 32 272
use FILL  FILL_5__2041_
timestamp 1701859473
transform -1 0 6950 0 -1 270
box -12 -8 32 272
use FILL  FILL_5__2042_
timestamp 1701859473
transform 1 0 8930 0 -1 790
box -12 -8 32 272
use FILL  FILL_5__2043_
timestamp 1701859473
transform 1 0 7250 0 1 270
box -12 -8 32 272
use FILL  FILL_5__2044_
timestamp 1701859473
transform 1 0 6990 0 1 270
box -12 -8 32 272
use FILL  FILL_5__2045_
timestamp 1701859473
transform -1 0 6310 0 1 270
box -12 -8 32 272
use FILL  FILL_5__2046_
timestamp 1701859473
transform 1 0 6490 0 -1 270
box -12 -8 32 272
use FILL  FILL_5__2047_
timestamp 1701859473
transform -1 0 6270 0 -1 270
box -12 -8 32 272
use FILL  FILL_5__2048_
timestamp 1701859473
transform -1 0 6070 0 -1 270
box -12 -8 32 272
use FILL  FILL_5__2049_
timestamp 1701859473
transform -1 0 7250 0 -1 790
box -12 -8 32 272
use FILL  FILL_5__2050_
timestamp 1701859473
transform 1 0 1490 0 -1 2870
box -12 -8 32 272
use FILL  FILL_5__2051_
timestamp 1701859473
transform 1 0 6290 0 -1 2350
box -12 -8 32 272
use FILL  FILL_5__2052_
timestamp 1701859473
transform -1 0 6190 0 1 790
box -12 -8 32 272
use FILL  FILL_5__2053_
timestamp 1701859473
transform -1 0 4410 0 1 1830
box -12 -8 32 272
use FILL  FILL_5__2054_
timestamp 1701859473
transform 1 0 2910 0 1 1310
box -12 -8 32 272
use FILL  FILL_5__2055_
timestamp 1701859473
transform -1 0 3170 0 1 1310
box -12 -8 32 272
use FILL  FILL_5__2056_
timestamp 1701859473
transform -1 0 1890 0 -1 1310
box -12 -8 32 272
use FILL  FILL_5__2057_
timestamp 1701859473
transform 1 0 2750 0 1 790
box -12 -8 32 272
use FILL  FILL_5__2058_
timestamp 1701859473
transform 1 0 3670 0 1 790
box -12 -8 32 272
use FILL  FILL_5__2059_
timestamp 1701859473
transform 1 0 3910 0 1 790
box -12 -8 32 272
use FILL  FILL_5__2060_
timestamp 1701859473
transform -1 0 4150 0 1 790
box -12 -8 32 272
use FILL  FILL_5__2061_
timestamp 1701859473
transform -1 0 3010 0 -1 270
box -12 -8 32 272
use FILL  FILL_5__2062_
timestamp 1701859473
transform 1 0 2790 0 1 270
box -12 -8 32 272
use FILL  FILL_5__2063_
timestamp 1701859473
transform 1 0 3170 0 -1 270
box -12 -8 32 272
use FILL  FILL_5__2064_
timestamp 1701859473
transform 1 0 3410 0 -1 270
box -12 -8 32 272
use FILL  FILL_5__2065_
timestamp 1701859473
transform -1 0 3650 0 -1 270
box -12 -8 32 272
use FILL  FILL_5__2066_
timestamp 1701859473
transform -1 0 5430 0 -1 270
box -12 -8 32 272
use FILL  FILL_5__2067_
timestamp 1701859473
transform 1 0 7370 0 1 790
box -12 -8 32 272
use FILL  FILL_5__2068_
timestamp 1701859473
transform 1 0 5930 0 1 790
box -12 -8 32 272
use FILL  FILL_5__2069_
timestamp 1701859473
transform 1 0 3410 0 -1 1830
box -12 -8 32 272
use FILL  FILL_5__2070_
timestamp 1701859473
transform -1 0 3890 0 -1 1830
box -12 -8 32 272
use FILL  FILL_5__2071_
timestamp 1701859473
transform -1 0 5730 0 1 790
box -12 -8 32 272
use FILL  FILL_5__2072_
timestamp 1701859473
transform -1 0 7790 0 1 1310
box -12 -8 32 272
use FILL  FILL_5__2073_
timestamp 1701859473
transform 1 0 6670 0 1 1310
box -12 -8 32 272
use FILL  FILL_5__2074_
timestamp 1701859473
transform 1 0 1810 0 1 1310
box -12 -8 32 272
use FILL  FILL_5__2075_
timestamp 1701859473
transform -1 0 2290 0 1 1310
box -12 -8 32 272
use FILL  FILL_5__2076_
timestamp 1701859473
transform -1 0 2330 0 -1 1310
box -12 -8 32 272
use FILL  FILL_5__2077_
timestamp 1701859473
transform 1 0 4190 0 -1 1310
box -12 -8 32 272
use FILL  FILL_5__2078_
timestamp 1701859473
transform -1 0 2330 0 1 1830
box -12 -8 32 272
use FILL  FILL_5__2079_
timestamp 1701859473
transform -1 0 970 0 -1 1830
box -12 -8 32 272
use FILL  FILL_5__2080_
timestamp 1701859473
transform 1 0 2290 0 -1 1830
box -12 -8 32 272
use FILL  FILL_5__2081_
timestamp 1701859473
transform 1 0 2530 0 -1 1830
box -12 -8 32 272
use FILL  FILL_5__2082_
timestamp 1701859473
transform -1 0 2750 0 -1 1830
box -12 -8 32 272
use FILL  FILL_5__2083_
timestamp 1701859473
transform 1 0 4430 0 -1 1310
box -12 -8 32 272
use FILL  FILL_5__2084_
timestamp 1701859473
transform -1 0 5270 0 1 790
box -12 -8 32 272
use FILL  FILL_5__2085_
timestamp 1701859473
transform -1 0 5110 0 -1 270
box -12 -8 32 272
use FILL  FILL_5__2086_
timestamp 1701859473
transform -1 0 4330 0 -1 270
box -12 -8 32 272
use FILL  FILL_5__2087_
timestamp 1701859473
transform -1 0 4810 0 1 790
box -12 -8 32 272
use FILL  FILL_5__2088_
timestamp 1701859473
transform -1 0 5650 0 1 270
box -12 -8 32 272
use FILL  FILL_5__2089_
timestamp 1701859473
transform 1 0 5410 0 1 270
box -12 -8 32 272
use FILL  FILL_5__2090_
timestamp 1701859473
transform -1 0 4990 0 -1 790
box -12 -8 32 272
use FILL  FILL_5__2091_
timestamp 1701859473
transform 1 0 3210 0 1 790
box -12 -8 32 272
use FILL  FILL_5__2092_
timestamp 1701859473
transform 1 0 2770 0 -1 270
box -12 -8 32 272
use FILL  FILL_5__2093_
timestamp 1701859473
transform -1 0 2930 0 -1 790
box -12 -8 32 272
use FILL  FILL_5__2094_
timestamp 1701859473
transform 1 0 2330 0 -1 270
box -12 -8 32 272
use FILL  FILL_5__2095_
timestamp 1701859473
transform 1 0 2530 0 -1 270
box -12 -8 32 272
use FILL  FILL_5__2096_
timestamp 1701859473
transform -1 0 4990 0 1 270
box -12 -8 32 272
use FILL  FILL_5__2097_
timestamp 1701859473
transform -1 0 5210 0 1 270
box -12 -8 32 272
use FILL  FILL_5__2098_
timestamp 1701859473
transform 1 0 4750 0 1 270
box -12 -8 32 272
use FILL  FILL_5__2099_
timestamp 1701859473
transform 1 0 4070 0 -1 270
box -12 -8 32 272
use FILL  FILL_5__2100_
timestamp 1701859473
transform -1 0 5930 0 -1 1830
box -12 -8 32 272
use FILL  FILL_5__2101_
timestamp 1701859473
transform -1 0 5850 0 1 1310
box -12 -8 32 272
use FILL  FILL_5__2102_
timestamp 1701859473
transform -1 0 6250 0 1 1310
box -12 -8 32 272
use FILL  FILL_5__2103_
timestamp 1701859473
transform 1 0 5810 0 -1 1310
box -12 -8 32 272
use FILL  FILL_5__2104_
timestamp 1701859473
transform -1 0 6050 0 1 1310
box -12 -8 32 272
use FILL  FILL_5__2105_
timestamp 1701859473
transform -1 0 4350 0 -1 1830
box -12 -8 32 272
use FILL  FILL_5__2106_
timestamp 1701859473
transform 1 0 4030 0 -1 790
box -12 -8 32 272
use FILL  FILL_5__2107_
timestamp 1701859473
transform -1 0 3610 0 -1 790
box -12 -8 32 272
use FILL  FILL_5__2108_
timestamp 1701859473
transform 1 0 2970 0 1 790
box -12 -8 32 272
use FILL  FILL_5__2109_
timestamp 1701859473
transform -1 0 3390 0 -1 790
box -12 -8 32 272
use FILL  FILL_5__2110_
timestamp 1701859473
transform 1 0 3150 0 -1 790
box -12 -8 32 272
use FILL  FILL_5__2111_
timestamp 1701859473
transform -1 0 3830 0 -1 790
box -12 -8 32 272
use FILL  FILL_5__2112_
timestamp 1701859473
transform -1 0 5190 0 -1 790
box -12 -8 32 272
use FILL  FILL_5__2113_
timestamp 1701859473
transform -1 0 5170 0 1 1310
box -12 -8 32 272
use FILL  FILL_5__2114_
timestamp 1701859473
transform -1 0 5610 0 1 1310
box -12 -8 32 272
use FILL  FILL_5__2115_
timestamp 1701859473
transform -1 0 5650 0 -1 790
box -12 -8 32 272
use FILL  FILL_5__2116_
timestamp 1701859473
transform 1 0 2470 0 1 1310
box -12 -8 32 272
use FILL  FILL_5__2117_
timestamp 1701859473
transform 1 0 2670 0 1 1310
box -12 -8 32 272
use FILL  FILL_5__2118_
timestamp 1701859473
transform 1 0 3850 0 1 1310
box -12 -8 32 272
use FILL  FILL_5__2119_
timestamp 1701859473
transform -1 0 4110 0 1 1310
box -12 -8 32 272
use FILL  FILL_5__2120_
timestamp 1701859473
transform 1 0 3970 0 -1 1310
box -12 -8 32 272
use FILL  FILL_5__2121_
timestamp 1701859473
transform -1 0 4550 0 1 270
box -12 -8 32 272
use FILL  FILL_5__2122_
timestamp 1701859473
transform -1 0 2890 0 1 2350
box -12 -8 32 272
use FILL  FILL_5__2123_
timestamp 1701859473
transform 1 0 2830 0 -1 2350
box -12 -8 32 272
use FILL  FILL_5__2124_
timestamp 1701859473
transform -1 0 3730 0 -1 2350
box -12 -8 32 272
use FILL  FILL_5__2125_
timestamp 1701859473
transform 1 0 5850 0 -1 3390
box -12 -8 32 272
use FILL  FILL_5__2126_
timestamp 1701859473
transform 1 0 5530 0 1 2870
box -12 -8 32 272
use FILL  FILL_5__2127_
timestamp 1701859473
transform -1 0 6010 0 1 2870
box -12 -8 32 272
use FILL  FILL_5__2128_
timestamp 1701859473
transform 1 0 4630 0 1 2870
box -12 -8 32 272
use FILL  FILL_5__2129_
timestamp 1701859473
transform 1 0 5310 0 1 2870
box -12 -8 32 272
use FILL  FILL_5__2130_
timestamp 1701859473
transform -1 0 4670 0 -1 2350
box -12 -8 32 272
use FILL  FILL_5__2131_
timestamp 1701859473
transform 1 0 4710 0 1 1310
box -12 -8 32 272
use FILL  FILL_5__2132_
timestamp 1701859473
transform -1 0 4590 0 1 790
box -12 -8 32 272
use FILL  FILL_5__2133_
timestamp 1701859473
transform 1 0 4510 0 -1 790
box -12 -8 32 272
use FILL  FILL_5__2134_
timestamp 1701859473
transform 1 0 3630 0 -1 2870
box -12 -8 32 272
use FILL  FILL_5__2135_
timestamp 1701859473
transform 1 0 4250 0 -1 3390
box -12 -8 32 272
use FILL  FILL_5__2136_
timestamp 1701859473
transform -1 0 2790 0 1 3390
box -12 -8 32 272
use FILL  FILL_5__2137_
timestamp 1701859473
transform 1 0 2350 0 1 3390
box -12 -8 32 272
use FILL  FILL_5__2138_
timestamp 1701859473
transform 1 0 3150 0 -1 4430
box -12 -8 32 272
use FILL  FILL_5__2139_
timestamp 1701859473
transform -1 0 2930 0 -1 4430
box -12 -8 32 272
use FILL  FILL_5__2140_
timestamp 1701859473
transform 1 0 2850 0 1 4430
box -12 -8 32 272
use FILL  FILL_5__2141_
timestamp 1701859473
transform -1 0 3090 0 1 4430
box -12 -8 32 272
use FILL  FILL_5__2142_
timestamp 1701859473
transform 1 0 2970 0 1 3390
box -12 -8 32 272
use FILL  FILL_5__2143_
timestamp 1701859473
transform -1 0 7470 0 -1 3390
box -12 -8 32 272
use FILL  FILL_5__2144_
timestamp 1701859473
transform 1 0 2110 0 1 2870
box -12 -8 32 272
use FILL  FILL_5__2145_
timestamp 1701859473
transform -1 0 10090 0 -1 2870
box -12 -8 32 272
use FILL  FILL_5__2146_
timestamp 1701859473
transform -1 0 7670 0 -1 3390
box -12 -8 32 272
use FILL  FILL_5__2147_
timestamp 1701859473
transform 1 0 7630 0 -1 3910
box -12 -8 32 272
use FILL  FILL_5__2148_
timestamp 1701859473
transform 1 0 7470 0 1 3390
box -12 -8 32 272
use FILL  FILL_5__2149_
timestamp 1701859473
transform 1 0 7670 0 1 3390
box -12 -8 32 272
use FILL  FILL_5__2150_
timestamp 1701859473
transform -1 0 7930 0 1 3390
box -12 -8 32 272
use FILL  FILL_5__2151_
timestamp 1701859473
transform 1 0 7210 0 -1 3390
box -12 -8 32 272
use FILL  FILL_5__2152_
timestamp 1701859473
transform 1 0 6970 0 -1 3390
box -12 -8 32 272
use FILL  FILL_5__2153_
timestamp 1701859473
transform -1 0 6110 0 -1 3390
box -12 -8 32 272
use FILL  FILL_5__2154_
timestamp 1701859473
transform 1 0 2870 0 -1 7030
box -12 -8 32 272
use FILL  FILL_5__2155_
timestamp 1701859473
transform 1 0 6430 0 1 5990
box -12 -8 32 272
use FILL  FILL_5__2156_
timestamp 1701859473
transform -1 0 4650 0 1 3910
box -12 -8 32 272
use FILL  FILL_5__2157_
timestamp 1701859473
transform -1 0 4790 0 -1 4430
box -12 -8 32 272
use FILL  FILL_5__2158_
timestamp 1701859473
transform -1 0 2650 0 1 2350
box -12 -8 32 272
use FILL  FILL_5__2159_
timestamp 1701859473
transform 1 0 3550 0 1 3910
box -12 -8 32 272
use FILL  FILL_5__2160_
timestamp 1701859473
transform -1 0 3870 0 -1 4430
box -12 -8 32 272
use FILL  FILL_5__2161_
timestamp 1701859473
transform -1 0 4010 0 1 3910
box -12 -8 32 272
use FILL  FILL_5__2162_
timestamp 1701859473
transform -1 0 4450 0 1 3910
box -12 -8 32 272
use FILL  FILL_5__2163_
timestamp 1701859473
transform 1 0 3770 0 -1 3910
box -12 -8 32 272
use FILL  FILL_5__2164_
timestamp 1701859473
transform -1 0 590 0 -1 4950
box -12 -8 32 272
use FILL  FILL_5__2165_
timestamp 1701859473
transform -1 0 3290 0 -1 3910
box -12 -8 32 272
use FILL  FILL_5__2166_
timestamp 1701859473
transform 1 0 3990 0 -1 3910
box -12 -8 32 272
use FILL  FILL_5__2167_
timestamp 1701859473
transform 1 0 4190 0 1 3910
box -12 -8 32 272
use FILL  FILL_5__2168_
timestamp 1701859473
transform 1 0 3110 0 1 3910
box -12 -8 32 272
use FILL  FILL_5__2169_
timestamp 1701859473
transform 1 0 2470 0 -1 4430
box -12 -8 32 272
use FILL  FILL_5__2170_
timestamp 1701859473
transform -1 0 2730 0 -1 4430
box -12 -8 32 272
use FILL  FILL_5__2171_
timestamp 1701859473
transform 1 0 4070 0 -1 4430
box -12 -8 32 272
use FILL  FILL_5__2172_
timestamp 1701859473
transform 1 0 4310 0 -1 4430
box -12 -8 32 272
use FILL  FILL_5__2173_
timestamp 1701859473
transform -1 0 4550 0 -1 4430
box -12 -8 32 272
use FILL  FILL_5__2174_
timestamp 1701859473
transform 1 0 6050 0 1 7030
box -12 -8 32 272
use FILL  FILL_5__2175_
timestamp 1701859473
transform -1 0 2550 0 1 8070
box -12 -8 32 272
use FILL  FILL_5__2176_
timestamp 1701859473
transform -1 0 6470 0 -1 8070
box -12 -8 32 272
use FILL  FILL_5__2177_
timestamp 1701859473
transform 1 0 4990 0 1 8070
box -12 -8 32 272
use FILL  FILL_5__2178_
timestamp 1701859473
transform -1 0 4170 0 -1 8590
box -12 -8 32 272
use FILL  FILL_5__2179_
timestamp 1701859473
transform -1 0 5990 0 -1 8070
box -12 -8 32 272
use FILL  FILL_5__2180_
timestamp 1701859473
transform -1 0 3010 0 -1 9630
box -12 -8 32 272
use FILL  FILL_5__2181_
timestamp 1701859473
transform 1 0 5070 0 1 7550
box -12 -8 32 272
use FILL  FILL_5__2182_
timestamp 1701859473
transform 1 0 5590 0 -1 10150
box -12 -8 32 272
use FILL  FILL_5__2183_
timestamp 1701859473
transform -1 0 3570 0 1 10150
box -12 -8 32 272
use FILL  FILL_5__2184_
timestamp 1701859473
transform 1 0 4390 0 1 8070
box -12 -8 32 272
use FILL  FILL_5__2185_
timestamp 1701859473
transform 1 0 5990 0 1 10150
box -12 -8 32 272
use FILL  FILL_5__2186_
timestamp 1701859473
transform 1 0 3550 0 1 10670
box -12 -8 32 272
use FILL  FILL_5__2187_
timestamp 1701859473
transform -1 0 5470 0 -1 10670
box -12 -8 32 272
use FILL  FILL_5__2188_
timestamp 1701859473
transform 1 0 2150 0 -1 10670
box -12 -8 32 272
use FILL  FILL_5__2189_
timestamp 1701859473
transform 1 0 5710 0 -1 10670
box -12 -8 32 272
use FILL  FILL_5__2190_
timestamp 1701859473
transform -1 0 2870 0 1 10150
box -12 -8 32 272
use FILL  FILL_5__2191_
timestamp 1701859473
transform -1 0 5350 0 -1 10150
box -12 -8 32 272
use FILL  FILL_5__2192_
timestamp 1701859473
transform -1 0 11150 0 1 3910
box -12 -8 32 272
use FILL  FILL_5__2193_
timestamp 1701859473
transform 1 0 1270 0 -1 3910
box -12 -8 32 272
use FILL  FILL_5__2194_
timestamp 1701859473
transform 1 0 1070 0 -1 3910
box -12 -8 32 272
use FILL  FILL_5__2195_
timestamp 1701859473
transform 1 0 2650 0 1 3910
box -12 -8 32 272
use FILL  FILL_5__2196_
timestamp 1701859473
transform 1 0 2890 0 1 3910
box -12 -8 32 272
use FILL  FILL_5__2197_
timestamp 1701859473
transform 1 0 5370 0 1 3910
box -12 -8 32 272
use FILL  FILL_5__2198_
timestamp 1701859473
transform 1 0 310 0 1 1830
box -12 -8 32 272
use FILL  FILL_5__2199_
timestamp 1701859473
transform -1 0 2870 0 -1 3910
box -12 -8 32 272
use FILL  FILL_5__2200_
timestamp 1701859473
transform 1 0 5390 0 -1 3910
box -12 -8 32 272
use FILL  FILL_5__2201_
timestamp 1701859473
transform -1 0 5630 0 1 3910
box -12 -8 32 272
use FILL  FILL_5__2202_
timestamp 1701859473
transform -1 0 8210 0 -1 4430
box -12 -8 32 272
use FILL  FILL_5__2203_
timestamp 1701859473
transform -1 0 4930 0 -1 3910
box -12 -8 32 272
use FILL  FILL_5__2204_
timestamp 1701859473
transform 1 0 5150 0 -1 3910
box -12 -8 32 272
use FILL  FILL_5__2205_
timestamp 1701859473
transform -1 0 9010 0 -1 3910
box -12 -8 32 272
use FILL  FILL_5__2206_
timestamp 1701859473
transform 1 0 9090 0 1 3910
box -12 -8 32 272
use FILL  FILL_5__2207_
timestamp 1701859473
transform 1 0 9550 0 -1 3910
box -12 -8 32 272
use FILL  FILL_5__2208_
timestamp 1701859473
transform -1 0 9810 0 -1 3910
box -12 -8 32 272
use FILL  FILL_5__2209_
timestamp 1701859473
transform -1 0 9610 0 1 4430
box -12 -8 32 272
use FILL  FILL_5__2210_
timestamp 1701859473
transform -1 0 10610 0 -1 4950
box -12 -8 32 272
use FILL  FILL_5__2211_
timestamp 1701859473
transform 1 0 9310 0 -1 3910
box -12 -8 32 272
use FILL  FILL_5__2212_
timestamp 1701859473
transform -1 0 8890 0 1 3910
box -12 -8 32 272
use FILL  FILL_5__2213_
timestamp 1701859473
transform -1 0 9330 0 1 3910
box -12 -8 32 272
use FILL  FILL_5__2214_
timestamp 1701859473
transform -1 0 9530 0 -1 4430
box -12 -8 32 272
use FILL  FILL_5__2215_
timestamp 1701859473
transform 1 0 9730 0 -1 4430
box -12 -8 32 272
use FILL  FILL_5__2216_
timestamp 1701859473
transform -1 0 9490 0 -1 7030
box -12 -8 32 272
use FILL  FILL_5__2217_
timestamp 1701859473
transform 1 0 9270 0 -1 4430
box -12 -8 32 272
use FILL  FILL_5__2218_
timestamp 1701859473
transform -1 0 9790 0 1 3910
box -12 -8 32 272
use FILL  FILL_5__2219_
timestamp 1701859473
transform 1 0 9970 0 1 3910
box -12 -8 32 272
use FILL  FILL_5__2220_
timestamp 1701859473
transform 1 0 10350 0 -1 4950
box -12 -8 32 272
use FILL  FILL_5__2221_
timestamp 1701859473
transform -1 0 9730 0 -1 7030
box -12 -8 32 272
use FILL  FILL_5__2222_
timestamp 1701859473
transform 1 0 10090 0 1 4430
box -12 -8 32 272
use FILL  FILL_5__2223_
timestamp 1701859473
transform -1 0 9990 0 -1 4430
box -12 -8 32 272
use FILL  FILL_5__2224_
timestamp 1701859473
transform -1 0 9850 0 1 4430
box -12 -8 32 272
use FILL  FILL_5__2225_
timestamp 1701859473
transform 1 0 10090 0 -1 4950
box -12 -8 32 272
use FILL  FILL_5__2226_
timestamp 1701859473
transform 1 0 8970 0 -1 7030
box -12 -8 32 272
use FILL  FILL_5__2227_
timestamp 1701859473
transform -1 0 9250 0 -1 7030
box -12 -8 32 272
use FILL  FILL_5__2228_
timestamp 1701859473
transform -1 0 5790 0 -1 7030
box -12 -8 32 272
use FILL  FILL_5__2229_
timestamp 1701859473
transform 1 0 4350 0 1 3390
box -12 -8 32 272
use FILL  FILL_5__2230_
timestamp 1701859473
transform -1 0 4450 0 -1 3910
box -12 -8 32 272
use FILL  FILL_5__2231_
timestamp 1701859473
transform -1 0 4230 0 -1 3910
box -12 -8 32 272
use FILL  FILL_5__2232_
timestamp 1701859473
transform 1 0 1630 0 1 2870
box -12 -8 32 272
use FILL  FILL_5__2233_
timestamp 1701859473
transform 1 0 2350 0 1 2870
box -12 -8 32 272
use FILL  FILL_5__2234_
timestamp 1701859473
transform -1 0 2610 0 1 2870
box -12 -8 32 272
use FILL  FILL_5__2235_
timestamp 1701859473
transform 1 0 6370 0 1 3390
box -12 -8 32 272
use FILL  FILL_5__2236_
timestamp 1701859473
transform -1 0 5650 0 -1 3910
box -12 -8 32 272
use FILL  FILL_5__2237_
timestamp 1701859473
transform -1 0 4690 0 -1 3910
box -12 -8 32 272
use FILL  FILL_5__2238_
timestamp 1701859473
transform 1 0 4750 0 -1 4950
box -12 -8 32 272
use FILL  FILL_5__2239_
timestamp 1701859473
transform 1 0 2870 0 1 4950
box -12 -8 32 272
use FILL  FILL_5__2240_
timestamp 1701859473
transform 1 0 2430 0 1 3910
box -12 -8 32 272
use FILL  FILL_5__2241_
timestamp 1701859473
transform -1 0 2450 0 1 4950
box -12 -8 32 272
use FILL  FILL_5__2242_
timestamp 1701859473
transform 1 0 2490 0 -1 4950
box -12 -8 32 272
use FILL  FILL_5__2243_
timestamp 1701859473
transform 1 0 2670 0 1 4950
box -12 -8 32 272
use FILL  FILL_5__2244_
timestamp 1701859473
transform 1 0 3090 0 1 4950
box -12 -8 32 272
use FILL  FILL_5__2245_
timestamp 1701859473
transform 1 0 2930 0 1 5990
box -12 -8 32 272
use FILL  FILL_5__2246_
timestamp 1701859473
transform 1 0 2950 0 -1 4950
box -12 -8 32 272
use FILL  FILL_5__2247_
timestamp 1701859473
transform -1 0 3070 0 -1 6510
box -12 -8 32 272
use FILL  FILL_5__2248_
timestamp 1701859473
transform 1 0 3530 0 -1 7030
box -12 -8 32 272
use FILL  FILL_5__2249_
timestamp 1701859473
transform 1 0 6310 0 1 7030
box -12 -8 32 272
use FILL  FILL_5__2250_
timestamp 1701859473
transform -1 0 10610 0 -1 7550
box -12 -8 32 272
use FILL  FILL_5__2251_
timestamp 1701859473
transform -1 0 10670 0 1 8070
box -12 -8 32 272
use FILL  FILL_5__2252_
timestamp 1701859473
transform -1 0 10970 0 -1 8070
box -12 -8 32 272
use FILL  FILL_5__2253_
timestamp 1701859473
transform -1 0 10730 0 -1 8070
box -12 -8 32 272
use FILL  FILL_5__2254_
timestamp 1701859473
transform 1 0 5430 0 1 8070
box -12 -8 32 272
use FILL  FILL_5__2255_
timestamp 1701859473
transform 1 0 3050 0 1 7030
box -12 -8 32 272
use FILL  FILL_5__2256_
timestamp 1701859473
transform -1 0 5170 0 1 7030
box -12 -8 32 272
use FILL  FILL_5__2257_
timestamp 1701859473
transform 1 0 5110 0 -1 7550
box -12 -8 32 272
use FILL  FILL_5__2258_
timestamp 1701859473
transform 1 0 5750 0 -1 8590
box -12 -8 32 272
use FILL  FILL_5__2259_
timestamp 1701859473
transform 1 0 10370 0 -1 7550
box -12 -8 32 272
use FILL  FILL_5__2260_
timestamp 1701859473
transform 1 0 9950 0 1 8070
box -12 -8 32 272
use FILL  FILL_5__2261_
timestamp 1701859473
transform -1 0 10250 0 1 7550
box -12 -8 32 272
use FILL  FILL_5__2262_
timestamp 1701859473
transform -1 0 10010 0 1 7550
box -12 -8 32 272
use FILL  FILL_5__2263_
timestamp 1701859473
transform 1 0 5510 0 1 7550
box -12 -8 32 272
use FILL  FILL_5__2264_
timestamp 1701859473
transform 1 0 1670 0 -1 6510
box -12 -8 32 272
use FILL  FILL_5__2265_
timestamp 1701859473
transform 1 0 1850 0 -1 6510
box -12 -8 32 272
use FILL  FILL_5__2266_
timestamp 1701859473
transform 1 0 3950 0 1 6510
box -12 -8 32 272
use FILL  FILL_5__2267_
timestamp 1701859473
transform -1 0 3710 0 -1 7550
box -12 -8 32 272
use FILL  FILL_5__2268_
timestamp 1701859473
transform 1 0 4390 0 -1 7550
box -12 -8 32 272
use FILL  FILL_5__2269_
timestamp 1701859473
transform 1 0 5710 0 1 7550
box -12 -8 32 272
use FILL  FILL_5__2270_
timestamp 1701859473
transform 1 0 8630 0 1 7550
box -12 -8 32 272
use FILL  FILL_5__2271_
timestamp 1701859473
transform -1 0 8910 0 -1 8070
box -12 -8 32 272
use FILL  FILL_5__2272_
timestamp 1701859473
transform -1 0 9170 0 -1 8070
box -12 -8 32 272
use FILL  FILL_5__2273_
timestamp 1701859473
transform -1 0 8670 0 -1 8070
box -12 -8 32 272
use FILL  FILL_5__2274_
timestamp 1701859473
transform -1 0 6030 0 -1 9630
box -12 -8 32 272
use FILL  FILL_5__2275_
timestamp 1701859473
transform -1 0 2330 0 1 8070
box -12 -8 32 272
use FILL  FILL_5__2276_
timestamp 1701859473
transform -1 0 3210 0 1 8070
box -12 -8 32 272
use FILL  FILL_5__2277_
timestamp 1701859473
transform -1 0 3690 0 -1 8590
box -12 -8 32 272
use FILL  FILL_5__2278_
timestamp 1701859473
transform 1 0 6590 0 1 9110
box -12 -8 32 272
use FILL  FILL_5__2279_
timestamp 1701859473
transform -1 0 10290 0 1 5990
box -12 -8 32 272
use FILL  FILL_5__2280_
timestamp 1701859473
transform 1 0 10470 0 1 5990
box -12 -8 32 272
use FILL  FILL_5__2281_
timestamp 1701859473
transform -1 0 10750 0 -1 5990
box -12 -8 32 272
use FILL  FILL_5__2282_
timestamp 1701859473
transform -1 0 10530 0 -1 6510
box -12 -8 32 272
use FILL  FILL_5__2283_
timestamp 1701859473
transform 1 0 5990 0 -1 8590
box -12 -8 32 272
use FILL  FILL_5__2284_
timestamp 1701859473
transform -1 0 2110 0 1 8070
box -12 -8 32 272
use FILL  FILL_5__2285_
timestamp 1701859473
transform -1 0 4170 0 1 8070
box -12 -8 32 272
use FILL  FILL_5__2286_
timestamp 1701859473
transform 1 0 5070 0 -1 8590
box -12 -8 32 272
use FILL  FILL_5__2287_
timestamp 1701859473
transform -1 0 6150 0 1 8590
box -12 -8 32 272
use FILL  FILL_5__2288_
timestamp 1701859473
transform -1 0 8870 0 1 7550
box -12 -8 32 272
use FILL  FILL_5__2289_
timestamp 1701859473
transform 1 0 8530 0 1 8070
box -12 -8 32 272
use FILL  FILL_5__2290_
timestamp 1701859473
transform -1 0 10030 0 -1 8070
box -12 -8 32 272
use FILL  FILL_5__2291_
timestamp 1701859473
transform -1 0 8810 0 1 8070
box -12 -8 32 272
use FILL  FILL_5__2292_
timestamp 1701859473
transform -1 0 6250 0 -1 9110
box -12 -8 32 272
use FILL  FILL_5__2293_
timestamp 1701859473
transform -1 0 2570 0 -1 8590
box -12 -8 32 272
use FILL  FILL_5__2294_
timestamp 1701859473
transform -1 0 4050 0 1 8590
box -12 -8 32 272
use FILL  FILL_5__2295_
timestamp 1701859473
transform 1 0 4970 0 1 8590
box -12 -8 32 272
use FILL  FILL_5__2296_
timestamp 1701859473
transform 1 0 6690 0 -1 9110
box -12 -8 32 272
use FILL  FILL_5__2297_
timestamp 1701859473
transform -1 0 9590 0 -1 5990
box -12 -8 32 272
use FILL  FILL_5__2298_
timestamp 1701859473
transform -1 0 10030 0 -1 5470
box -12 -8 32 272
use FILL  FILL_5__2299_
timestamp 1701859473
transform -1 0 9370 0 -1 6510
box -12 -8 32 272
use FILL  FILL_5__2300_
timestamp 1701859473
transform 1 0 9570 0 1 5990
box -12 -8 32 272
use FILL  FILL_5__2301_
timestamp 1701859473
transform 1 0 5610 0 1 9630
box -12 -8 32 272
use FILL  FILL_5__2302_
timestamp 1701859473
transform -1 0 3510 0 -1 9110
box -12 -8 32 272
use FILL  FILL_5__2303_
timestamp 1701859473
transform 1 0 2630 0 1 9110
box -12 -8 32 272
use FILL  FILL_5__2304_
timestamp 1701859473
transform 1 0 2830 0 -1 9110
box -12 -8 32 272
use FILL  FILL_5__2305_
timestamp 1701859473
transform -1 0 3810 0 1 8590
box -12 -8 32 272
use FILL  FILL_5__2306_
timestamp 1701859473
transform 1 0 4490 0 1 8590
box -12 -8 32 272
use FILL  FILL_5__2307_
timestamp 1701859473
transform 1 0 6350 0 1 9110
box -12 -8 32 272
use FILL  FILL_5__2308_
timestamp 1701859473
transform -1 0 8930 0 -1 6510
box -12 -8 32 272
use FILL  FILL_5__2309_
timestamp 1701859473
transform -1 0 8630 0 1 5990
box -12 -8 32 272
use FILL  FILL_5__2310_
timestamp 1701859473
transform -1 0 9130 0 -1 6510
box -12 -8 32 272
use FILL  FILL_5__2311_
timestamp 1701859473
transform -1 0 8690 0 -1 6510
box -12 -8 32 272
use FILL  FILL_5__2312_
timestamp 1701859473
transform -1 0 5590 0 -1 9630
box -12 -8 32 272
use FILL  FILL_5__2313_
timestamp 1701859473
transform -1 0 1870 0 1 8590
box -12 -8 32 272
use FILL  FILL_5__2314_
timestamp 1701859473
transform 1 0 1470 0 -1 8590
box -12 -8 32 272
use FILL  FILL_5__2315_
timestamp 1701859473
transform 1 0 1910 0 -1 8590
box -12 -8 32 272
use FILL  FILL_5__2316_
timestamp 1701859473
transform -1 0 4270 0 1 8590
box -12 -8 32 272
use FILL  FILL_5__2317_
timestamp 1701859473
transform 1 0 4730 0 1 8590
box -12 -8 32 272
use FILL  FILL_5__2318_
timestamp 1701859473
transform 1 0 6830 0 1 9110
box -12 -8 32 272
use FILL  FILL_5__2319_
timestamp 1701859473
transform -1 0 11150 0 1 4430
box -12 -8 32 272
use FILL  FILL_5__2320_
timestamp 1701859473
transform 1 0 5130 0 1 3910
box -12 -8 32 272
use FILL  FILL_5__2321_
timestamp 1701859473
transform 1 0 6550 0 1 3910
box -12 -8 32 272
use FILL  FILL_5__2322_
timestamp 1701859473
transform -1 0 7930 0 1 3910
box -12 -8 32 272
use FILL  FILL_5__2323_
timestamp 1701859473
transform 1 0 7970 0 -1 4430
box -12 -8 32 272
use FILL  FILL_5__2324_
timestamp 1701859473
transform -1 0 11190 0 -1 2870
box -12 -8 32 272
use FILL  FILL_5__2325_
timestamp 1701859473
transform -1 0 8170 0 1 3910
box -12 -8 32 272
use FILL  FILL_5__2326_
timestamp 1701859473
transform -1 0 3210 0 -1 4950
box -12 -8 32 272
use FILL  FILL_5__2327_
timestamp 1701859473
transform -1 0 3410 0 -1 4950
box -12 -8 32 272
use FILL  FILL_5__2328_
timestamp 1701859473
transform 1 0 3890 0 -1 5470
box -12 -8 32 272
use FILL  FILL_5__2329_
timestamp 1701859473
transform 1 0 3650 0 -1 5470
box -12 -8 32 272
use FILL  FILL_5__2330_
timestamp 1701859473
transform 1 0 3790 0 1 4950
box -12 -8 32 272
use FILL  FILL_5__2331_
timestamp 1701859473
transform 1 0 4870 0 1 3910
box -12 -8 32 272
use FILL  FILL_5__2332_
timestamp 1701859473
transform -1 0 4210 0 1 4950
box -12 -8 32 272
use FILL  FILL_5__2333_
timestamp 1701859473
transform -1 0 11170 0 -1 4430
box -12 -8 32 272
use FILL  FILL_5__2334_
timestamp 1701859473
transform 1 0 9050 0 -1 4430
box -12 -8 32 272
use FILL  FILL_5__2335_
timestamp 1701859473
transform 1 0 5230 0 -1 5470
box -12 -8 32 272
use FILL  FILL_5__2336_
timestamp 1701859473
transform -1 0 5090 0 1 5990
box -12 -8 32 272
use FILL  FILL_5__2337_
timestamp 1701859473
transform 1 0 4590 0 1 3390
box -12 -8 32 272
use FILL  FILL_5__2338_
timestamp 1701859473
transform 1 0 3190 0 1 3390
box -12 -8 32 272
use FILL  FILL_5__2339_
timestamp 1701859473
transform 1 0 4770 0 1 3390
box -12 -8 32 272
use FILL  FILL_5__2340_
timestamp 1701859473
transform 1 0 5010 0 1 3390
box -12 -8 32 272
use FILL  FILL_5__2341_
timestamp 1701859473
transform -1 0 590 0 1 5990
box -12 -8 32 272
use FILL  FILL_5__2342_
timestamp 1701859473
transform 1 0 2690 0 1 5470
box -12 -8 32 272
use FILL  FILL_5__2343_
timestamp 1701859473
transform -1 0 4630 0 1 6510
box -12 -8 32 272
use FILL  FILL_5__2344_
timestamp 1701859473
transform -1 0 4910 0 1 5470
box -12 -8 32 272
use FILL  FILL_5__2345_
timestamp 1701859473
transform -1 0 4710 0 1 5470
box -12 -8 32 272
use FILL  FILL_5__2346_
timestamp 1701859473
transform -1 0 4870 0 -1 5990
box -12 -8 32 272
use FILL  FILL_5__2347_
timestamp 1701859473
transform -1 0 5730 0 -1 5990
box -12 -8 32 272
use FILL  FILL_5__2348_
timestamp 1701859473
transform 1 0 5290 0 -1 6510
box -12 -8 32 272
use FILL  FILL_5__2349_
timestamp 1701859473
transform -1 0 5070 0 -1 6510
box -12 -8 32 272
use FILL  FILL_5__2350_
timestamp 1701859473
transform -1 0 4490 0 -1 6510
box -12 -8 32 272
use FILL  FILL_5__2351_
timestamp 1701859473
transform 1 0 5630 0 1 7030
box -12 -8 32 272
use FILL  FILL_5__2352_
timestamp 1701859473
transform -1 0 5850 0 1 7030
box -12 -8 32 272
use FILL  FILL_5__2353_
timestamp 1701859473
transform -1 0 790 0 1 7030
box -12 -8 32 272
use FILL  FILL_5__2354_
timestamp 1701859473
transform 1 0 5490 0 -1 5990
box -12 -8 32 272
use FILL  FILL_5__2355_
timestamp 1701859473
transform 1 0 5390 0 1 7030
box -12 -8 32 272
use FILL  FILL_5__2356_
timestamp 1701859473
transform -1 0 4890 0 -1 7550
box -12 -8 32 272
use FILL  FILL_5__2357_
timestamp 1701859473
transform 1 0 4750 0 1 8070
box -12 -8 32 272
use FILL  FILL_5__2358_
timestamp 1701859473
transform 1 0 5230 0 1 8070
box -12 -8 32 272
use FILL  FILL_5__2359_
timestamp 1701859473
transform -1 0 5550 0 -1 8590
box -12 -8 32 272
use FILL  FILL_5__2360_
timestamp 1701859473
transform -1 0 790 0 -1 6510
box -12 -8 32 272
use FILL  FILL_5__2361_
timestamp 1701859473
transform -1 0 5290 0 1 5990
box -12 -8 32 272
use FILL  FILL_5__2362_
timestamp 1701859473
transform 1 0 5290 0 1 6510
box -12 -8 32 272
use FILL  FILL_5__2363_
timestamp 1701859473
transform 1 0 5310 0 -1 7030
box -12 -8 32 272
use FILL  FILL_5__2364_
timestamp 1701859473
transform 1 0 5310 0 -1 8070
box -12 -8 32 272
use FILL  FILL_5__2365_
timestamp 1701859473
transform 1 0 5550 0 -1 8070
box -12 -8 32 272
use FILL  FILL_5__2366_
timestamp 1701859473
transform -1 0 5770 0 -1 8070
box -12 -8 32 272
use FILL  FILL_5__2367_
timestamp 1701859473
transform 1 0 2730 0 -1 7550
box -12 -8 32 272
use FILL  FILL_5__2368_
timestamp 1701859473
transform -1 0 5570 0 -1 7030
box -12 -8 32 272
use FILL  FILL_5__2369_
timestamp 1701859473
transform 1 0 5270 0 1 7550
box -12 -8 32 272
use FILL  FILL_5__2370_
timestamp 1701859473
transform -1 0 5310 0 -1 8590
box -12 -8 32 272
use FILL  FILL_5__2371_
timestamp 1701859473
transform 1 0 5990 0 -1 9110
box -12 -8 32 272
use FILL  FILL_5__2372_
timestamp 1701859473
transform 1 0 6150 0 1 9110
box -12 -8 32 272
use FILL  FILL_5__2373_
timestamp 1701859473
transform -1 0 6230 0 -1 9630
box -12 -8 32 272
use FILL  FILL_5__2374_
timestamp 1701859473
transform 1 0 110 0 -1 9110
box -12 -8 32 272
use FILL  FILL_5__2375_
timestamp 1701859473
transform -1 0 4250 0 1 5470
box -12 -8 32 272
use FILL  FILL_5__2376_
timestamp 1701859473
transform 1 0 4590 0 -1 5990
box -12 -8 32 272
use FILL  FILL_5__2377_
timestamp 1701859473
transform -1 0 4010 0 -1 6510
box -12 -8 32 272
use FILL  FILL_5__2378_
timestamp 1701859473
transform 1 0 3750 0 -1 6510
box -12 -8 32 272
use FILL  FILL_5__2379_
timestamp 1701859473
transform -1 0 5070 0 1 6510
box -12 -8 32 272
use FILL  FILL_5__2380_
timestamp 1701859473
transform -1 0 4850 0 -1 8590
box -12 -8 32 272
use FILL  FILL_5__2381_
timestamp 1701859473
transform 1 0 3910 0 -1 8590
box -12 -8 32 272
use FILL  FILL_5__2382_
timestamp 1701859473
transform -1 0 4610 0 -1 8590
box -12 -8 32 272
use FILL  FILL_5__2383_
timestamp 1701859473
transform -1 0 5690 0 1 8590
box -12 -8 32 272
use FILL  FILL_5__2384_
timestamp 1701859473
transform -1 0 5910 0 1 8590
box -12 -8 32 272
use FILL  FILL_5__2385_
timestamp 1701859473
transform 1 0 1290 0 -1 10150
box -12 -8 32 272
use FILL  FILL_5__2386_
timestamp 1701859473
transform 1 0 5550 0 -1 7550
box -12 -8 32 272
use FILL  FILL_5__2387_
timestamp 1701859473
transform 1 0 5530 0 -1 9110
box -12 -8 32 272
use FILL  FILL_5__2388_
timestamp 1701859473
transform -1 0 5330 0 -1 9110
box -12 -8 32 272
use FILL  FILL_5__2389_
timestamp 1701859473
transform -1 0 5110 0 -1 9630
box -12 -8 32 272
use FILL  FILL_5__2390_
timestamp 1701859473
transform 1 0 5170 0 1 9630
box -12 -8 32 272
use FILL  FILL_5__2391_
timestamp 1701859473
transform -1 0 5390 0 1 9630
box -12 -8 32 272
use FILL  FILL_5__2392_
timestamp 1701859473
transform 1 0 1490 0 -1 10150
box -12 -8 32 272
use FILL  FILL_5__2393_
timestamp 1701859473
transform -1 0 5350 0 -1 7550
box -12 -8 32 272
use FILL  FILL_5__2394_
timestamp 1701859473
transform 1 0 5430 0 1 8590
box -12 -8 32 272
use FILL  FILL_5__2395_
timestamp 1701859473
transform -1 0 5790 0 -1 9110
box -12 -8 32 272
use FILL  FILL_5__2396_
timestamp 1701859473
transform 1 0 5710 0 1 9110
box -12 -8 32 272
use FILL  FILL_5__2397_
timestamp 1701859473
transform 1 0 5950 0 1 9110
box -12 -8 32 272
use FILL  FILL_5__2398_
timestamp 1701859473
transform 1 0 5770 0 -1 9630
box -12 -8 32 272
use FILL  FILL_5__2399_
timestamp 1701859473
transform -1 0 3210 0 -1 5470
box -12 -8 32 272
use FILL  FILL_5__2400_
timestamp 1701859473
transform -1 0 3390 0 1 5990
box -12 -8 32 272
use FILL  FILL_5__2401_
timestamp 1701859473
transform 1 0 3310 0 -1 6510
box -12 -8 32 272
use FILL  FILL_5__2402_
timestamp 1701859473
transform -1 0 2250 0 -1 4430
box -12 -8 32 272
use FILL  FILL_5__2403_
timestamp 1701859473
transform -1 0 2650 0 1 4430
box -12 -8 32 272
use FILL  FILL_5__2404_
timestamp 1701859473
transform -1 0 2970 0 -1 5470
box -12 -8 32 272
use FILL  FILL_5__2405_
timestamp 1701859473
transform 1 0 2350 0 -1 2870
box -12 -8 32 272
use FILL  FILL_5__2406_
timestamp 1701859473
transform 1 0 3050 0 -1 3390
box -12 -8 32 272
use FILL  FILL_5__2407_
timestamp 1701859473
transform -1 0 3190 0 1 5470
box -12 -8 32 272
use FILL  FILL_5__2408_
timestamp 1701859473
transform 1 0 810 0 -1 2870
box -12 -8 32 272
use FILL  FILL_5__2409_
timestamp 1701859473
transform 1 0 830 0 -1 3910
box -12 -8 32 272
use FILL  FILL_5__2410_
timestamp 1701859473
transform 1 0 1230 0 1 4430
box -12 -8 32 272
use FILL  FILL_5__2411_
timestamp 1701859473
transform -1 0 790 0 -1 4950
box -12 -8 32 272
use FILL  FILL_5__2412_
timestamp 1701859473
transform 1 0 2470 0 -1 5990
box -12 -8 32 272
use FILL  FILL_5__2413_
timestamp 1701859473
transform 1 0 2930 0 1 5470
box -12 -8 32 272
use FILL  FILL_5__2414_
timestamp 1701859473
transform 1 0 4090 0 -1 5470
box -12 -8 32 272
use FILL  FILL_5__2415_
timestamp 1701859473
transform -1 0 4030 0 1 7030
box -12 -8 32 272
use FILL  FILL_5__2416_
timestamp 1701859473
transform 1 0 3990 0 1 4950
box -12 -8 32 272
use FILL  FILL_5__2417_
timestamp 1701859473
transform 1 0 4330 0 -1 5470
box -12 -8 32 272
use FILL  FILL_5__2418_
timestamp 1701859473
transform -1 0 1590 0 -1 4950
box -12 -8 32 272
use FILL  FILL_5__2419_
timestamp 1701859473
transform 1 0 2170 0 1 4430
box -12 -8 32 272
use FILL  FILL_5__2420_
timestamp 1701859473
transform 1 0 3830 0 1 5990
box -12 -8 32 272
use FILL  FILL_5__2421_
timestamp 1701859473
transform -1 0 3610 0 1 5990
box -12 -8 32 272
use FILL  FILL_5__2422_
timestamp 1701859473
transform -1 0 3490 0 -1 5990
box -12 -8 32 272
use FILL  FILL_5__2423_
timestamp 1701859473
transform -1 0 3710 0 -1 5990
box -12 -8 32 272
use FILL  FILL_5__2424_
timestamp 1701859473
transform 1 0 3250 0 -1 5990
box -12 -8 32 272
use FILL  FILL_5__2425_
timestamp 1701859473
transform 1 0 4390 0 1 5990
box -12 -8 32 272
use FILL  FILL_5__2426_
timestamp 1701859473
transform 1 0 3990 0 -1 7030
box -12 -8 32 272
use FILL  FILL_5__2427_
timestamp 1701859473
transform 1 0 4810 0 1 5990
box -12 -8 32 272
use FILL  FILL_5__2428_
timestamp 1701859473
transform 1 0 4570 0 1 5990
box -12 -8 32 272
use FILL  FILL_5__2429_
timestamp 1701859473
transform -1 0 4250 0 -1 6510
box -12 -8 32 272
use FILL  FILL_5__2430_
timestamp 1701859473
transform 1 0 4810 0 1 6510
box -12 -8 32 272
use FILL  FILL_5__2431_
timestamp 1701859473
transform -1 0 4910 0 -1 7030
box -12 -8 32 272
use FILL  FILL_5__2432_
timestamp 1701859473
transform 1 0 5130 0 -1 7030
box -12 -8 32 272
use FILL  FILL_5__2433_
timestamp 1701859473
transform -1 0 4390 0 -1 8070
box -12 -8 32 272
use FILL  FILL_5__2434_
timestamp 1701859473
transform 1 0 4870 0 1 7550
box -12 -8 32 272
use FILL  FILL_5__2435_
timestamp 1701859473
transform 1 0 4210 0 1 7030
box -12 -8 32 272
use FILL  FILL_5__2436_
timestamp 1701859473
transform -1 0 4650 0 -1 7550
box -12 -8 32 272
use FILL  FILL_5__2437_
timestamp 1701859473
transform -1 0 4630 0 -1 8070
box -12 -8 32 272
use FILL  FILL_5__2438_
timestamp 1701859473
transform -1 0 4870 0 -1 8070
box -12 -8 32 272
use FILL  FILL_5__2439_
timestamp 1701859473
transform -1 0 5110 0 -1 8070
box -12 -8 32 272
use FILL  FILL_5__2440_
timestamp 1701859473
transform 1 0 4650 0 1 10150
box -12 -8 32 272
use FILL  FILL_5__2441_
timestamp 1701859473
transform 1 0 3930 0 -1 7550
box -12 -8 32 272
use FILL  FILL_5__2442_
timestamp 1701859473
transform -1 0 4150 0 -1 8070
box -12 -8 32 272
use FILL  FILL_5__2443_
timestamp 1701859473
transform -1 0 3930 0 1 8070
box -12 -8 32 272
use FILL  FILL_5__2444_
timestamp 1701859473
transform 1 0 3670 0 1 8070
box -12 -8 32 272
use FILL  FILL_5__2445_
timestamp 1701859473
transform -1 0 4650 0 1 7550
box -12 -8 32 272
use FILL  FILL_5__2446_
timestamp 1701859473
transform 1 0 4570 0 1 8070
box -12 -8 32 272
use FILL  FILL_5__2447_
timestamp 1701859473
transform 1 0 4310 0 1 9110
box -12 -8 32 272
use FILL  FILL_5__2448_
timestamp 1701859473
transform 1 0 4970 0 1 9110
box -12 -8 32 272
use FILL  FILL_5__2449_
timestamp 1701859473
transform 1 0 5230 0 1 9110
box -12 -8 32 272
use FILL  FILL_5__2450_
timestamp 1701859473
transform 1 0 5470 0 1 9110
box -12 -8 32 272
use FILL  FILL_5__2451_
timestamp 1701859473
transform -1 0 5350 0 -1 9630
box -12 -8 32 272
use FILL  FILL_5__2452_
timestamp 1701859473
transform -1 0 5270 0 -1 10670
box -12 -8 32 272
use FILL  FILL_5__2453_
timestamp 1701859473
transform 1 0 3810 0 -1 10150
box -12 -8 32 272
use FILL  FILL_5__2454_
timestamp 1701859473
transform 1 0 3930 0 1 7550
box -12 -8 32 272
use FILL  FILL_5__2455_
timestamp 1701859473
transform 1 0 3890 0 -1 8070
box -12 -8 32 272
use FILL  FILL_5__2456_
timestamp 1701859473
transform -1 0 3670 0 -1 8070
box -12 -8 32 272
use FILL  FILL_5__2457_
timestamp 1701859473
transform 1 0 3430 0 1 8070
box -12 -8 32 272
use FILL  FILL_5__2458_
timestamp 1701859473
transform -1 0 4370 0 -1 8590
box -12 -8 32 272
use FILL  FILL_5__2459_
timestamp 1701859473
transform -1 0 4530 0 -1 11190
box -12 -8 32 272
use FILL  FILL_5__2460_
timestamp 1701859473
transform 1 0 4170 0 -1 10670
box -12 -8 32 272
use FILL  FILL_5__2461_
timestamp 1701859473
transform 1 0 4350 0 -1 9110
box -12 -8 32 272
use FILL  FILL_5__2462_
timestamp 1701859473
transform -1 0 4610 0 -1 9110
box -12 -8 32 272
use FILL  FILL_5__2463_
timestamp 1701859473
transform -1 0 4850 0 -1 9110
box -12 -8 32 272
use FILL  FILL_5__2464_
timestamp 1701859473
transform -1 0 5090 0 -1 9110
box -12 -8 32 272
use FILL  FILL_5__2465_
timestamp 1701859473
transform -1 0 4950 0 -1 11190
box -12 -8 32 272
use FILL  FILL_5__2466_
timestamp 1701859473
transform -1 0 4030 0 -1 10150
box -12 -8 32 272
use FILL  FILL_5__2467_
timestamp 1701859473
transform -1 0 4130 0 -1 9630
box -12 -8 32 272
use FILL  FILL_5__2468_
timestamp 1701859473
transform -1 0 4390 0 -1 9630
box -12 -8 32 272
use FILL  FILL_5__2469_
timestamp 1701859473
transform -1 0 4250 0 1 9630
box -12 -8 32 272
use FILL  FILL_5__2470_
timestamp 1701859473
transform -1 0 4490 0 1 9630
box -12 -8 32 272
use FILL  FILL_5__2471_
timestamp 1701859473
transform -1 0 5070 0 -1 10670
box -12 -8 32 272
use FILL  FILL_5__2472_
timestamp 1701859473
transform 1 0 4030 0 1 9630
box -12 -8 32 272
use FILL  FILL_5__2473_
timestamp 1701859473
transform 1 0 4590 0 -1 9630
box -12 -8 32 272
use FILL  FILL_5__2474_
timestamp 1701859473
transform -1 0 4870 0 -1 9630
box -12 -8 32 272
use FILL  FILL_5__2475_
timestamp 1701859473
transform 1 0 4710 0 1 9630
box -12 -8 32 272
use FILL  FILL_5__2476_
timestamp 1701859473
transform -1 0 4950 0 1 9630
box -12 -8 32 272
use FILL  FILL_5__2477_
timestamp 1701859473
transform 1 0 4890 0 1 10670
box -12 -8 32 272
use FILL  FILL_5__2478_
timestamp 1701859473
transform 1 0 3130 0 1 5990
box -12 -8 32 272
use FILL  FILL_5__2479_
timestamp 1701859473
transform -1 0 2690 0 1 5990
box -12 -8 32 272
use FILL  FILL_5__2480_
timestamp 1701859473
transform -1 0 2710 0 -1 5990
box -12 -8 32 272
use FILL  FILL_5__2481_
timestamp 1701859473
transform -1 0 2950 0 -1 5990
box -12 -8 32 272
use FILL  FILL_5__2482_
timestamp 1701859473
transform 1 0 1530 0 -1 5990
box -12 -8 32 272
use FILL  FILL_5__2483_
timestamp 1701859473
transform 1 0 2350 0 1 6510
box -12 -8 32 272
use FILL  FILL_5__2484_
timestamp 1701859473
transform -1 0 1970 0 1 6510
box -12 -8 32 272
use FILL  FILL_5__2485_
timestamp 1701859473
transform -1 0 2170 0 1 6510
box -12 -8 32 272
use FILL  FILL_5__2486_
timestamp 1701859473
transform 1 0 2370 0 -1 7030
box -12 -8 32 272
use FILL  FILL_5__2487_
timestamp 1701859473
transform 1 0 2130 0 -1 7030
box -12 -8 32 272
use FILL  FILL_5__2488_
timestamp 1701859473
transform -1 0 1930 0 -1 7030
box -12 -8 32 272
use FILL  FILL_5__2489_
timestamp 1701859473
transform 1 0 1430 0 -1 7030
box -12 -8 32 272
use FILL  FILL_5__2490_
timestamp 1701859473
transform -1 0 1030 0 1 5470
box -12 -8 32 272
use FILL  FILL_5__2491_
timestamp 1701859473
transform 1 0 1230 0 1 5470
box -12 -8 32 272
use FILL  FILL_5__2492_
timestamp 1701859473
transform -1 0 2090 0 -1 6510
box -12 -8 32 272
use FILL  FILL_5__2493_
timestamp 1701859473
transform 1 0 1970 0 1 5990
box -12 -8 32 272
use FILL  FILL_5__2494_
timestamp 1701859473
transform -1 0 1530 0 1 5990
box -12 -8 32 272
use FILL  FILL_5__2495_
timestamp 1701859473
transform 1 0 1270 0 1 5990
box -12 -8 32 272
use FILL  FILL_5__2496_
timestamp 1701859473
transform 1 0 1670 0 -1 7030
box -12 -8 32 272
use FILL  FILL_5__2497_
timestamp 1701859473
transform -1 0 1870 0 -1 7550
box -12 -8 32 272
use FILL  FILL_5__2498_
timestamp 1701859473
transform 1 0 810 0 1 8070
box -12 -8 32 272
use FILL  FILL_5__2499_
timestamp 1701859473
transform 1 0 2490 0 1 7550
box -12 -8 32 272
use FILL  FILL_5__2500_
timestamp 1701859473
transform 1 0 1910 0 1 7550
box -12 -8 32 272
use FILL  FILL_5__2501_
timestamp 1701859473
transform 1 0 1690 0 1 7550
box -12 -8 32 272
use FILL  FILL_5__2502_
timestamp 1701859473
transform -1 0 1230 0 1 7550
box -12 -8 32 272
use FILL  FILL_5__2503_
timestamp 1701859473
transform -1 0 1470 0 1 8070
box -12 -8 32 272
use FILL  FILL_5__2504_
timestamp 1701859473
transform -1 0 1890 0 1 8070
box -12 -8 32 272
use FILL  FILL_5__2505_
timestamp 1701859473
transform 1 0 1230 0 1 8070
box -12 -8 32 272
use FILL  FILL_5__2506_
timestamp 1701859473
transform -1 0 1750 0 -1 8070
box -12 -8 32 272
use FILL  FILL_5__2507_
timestamp 1701859473
transform 1 0 1490 0 -1 8070
box -12 -8 32 272
use FILL  FILL_5__2508_
timestamp 1701859473
transform 1 0 1010 0 1 8070
box -12 -8 32 272
use FILL  FILL_5__2509_
timestamp 1701859473
transform 1 0 570 0 -1 8590
box -12 -8 32 272
use FILL  FILL_5__2510_
timestamp 1701859473
transform -1 0 1510 0 1 9110
box -12 -8 32 272
use FILL  FILL_5__2511_
timestamp 1701859473
transform -1 0 1450 0 -1 9630
box -12 -8 32 272
use FILL  FILL_5__2512_
timestamp 1701859473
transform 1 0 1010 0 -1 9630
box -12 -8 32 272
use FILL  FILL_5__2513_
timestamp 1701859473
transform -1 0 1010 0 1 8590
box -12 -8 32 272
use FILL  FILL_5__2514_
timestamp 1701859473
transform 1 0 2090 0 -1 8590
box -12 -8 32 272
use FILL  FILL_5__2515_
timestamp 1701859473
transform 1 0 1210 0 -1 9110
box -12 -8 32 272
use FILL  FILL_5__2516_
timestamp 1701859473
transform -1 0 1050 0 1 9110
box -12 -8 32 272
use FILL  FILL_5__2517_
timestamp 1701859473
transform -1 0 810 0 1 9110
box -12 -8 32 272
use FILL  FILL_5__2518_
timestamp 1701859473
transform 1 0 1670 0 -1 9630
box -12 -8 32 272
use FILL  FILL_5__2519_
timestamp 1701859473
transform 1 0 1770 0 1 9630
box -12 -8 32 272
use FILL  FILL_5__2520_
timestamp 1701859473
transform -1 0 2610 0 -1 9110
box -12 -8 32 272
use FILL  FILL_5__2521_
timestamp 1701859473
transform 1 0 2350 0 -1 9110
box -12 -8 32 272
use FILL  FILL_5__2522_
timestamp 1701859473
transform -1 0 1970 0 1 9630
box -12 -8 32 272
use FILL  FILL_5__2523_
timestamp 1701859473
transform -1 0 2190 0 1 9630
box -12 -8 32 272
use FILL  FILL_5__2524_
timestamp 1701859473
transform -1 0 1930 0 -1 9110
box -12 -8 32 272
use FILL  FILL_5__2525_
timestamp 1701859473
transform 1 0 810 0 -1 8590
box -12 -8 32 272
use FILL  FILL_5__2526_
timestamp 1701859473
transform -1 0 1710 0 -1 8590
box -12 -8 32 272
use FILL  FILL_5__2527_
timestamp 1701859473
transform -1 0 1250 0 -1 8590
box -12 -8 32 272
use FILL  FILL_5__2528_
timestamp 1701859473
transform -1 0 1030 0 -1 8590
box -12 -8 32 272
use FILL  FILL_5__2529_
timestamp 1701859473
transform -1 0 1270 0 1 9110
box -12 -8 32 272
use FILL  FILL_5__2530_
timestamp 1701859473
transform -1 0 7530 0 -1 6510
box -12 -8 32 272
use FILL  FILL_5__2531_
timestamp 1701859473
transform 1 0 7950 0 1 7550
box -12 -8 32 272
use FILL  FILL_5__2532_
timestamp 1701859473
transform -1 0 9850 0 1 2870
box -12 -8 32 272
use FILL  FILL_5__2533_
timestamp 1701859473
transform -1 0 8930 0 1 4430
box -12 -8 32 272
use FILL  FILL_5__2534_
timestamp 1701859473
transform -1 0 9330 0 -1 5470
box -12 -8 32 272
use FILL  FILL_5__2535_
timestamp 1701859473
transform 1 0 110 0 -1 4950
box -12 -8 32 272
use FILL  FILL_5__2536_
timestamp 1701859473
transform 1 0 670 0 1 4950
box -12 -8 32 272
use FILL  FILL_5__2537_
timestamp 1701859473
transform 1 0 810 0 1 3390
box -12 -8 32 272
use FILL  FILL_5__2538_
timestamp 1701859473
transform -1 0 370 0 -1 3910
box -12 -8 32 272
use FILL  FILL_5__2539_
timestamp 1701859473
transform -1 0 130 0 1 4950
box -12 -8 32 272
use FILL  FILL_5__2540_
timestamp 1701859473
transform 1 0 3070 0 1 2350
box -12 -8 32 272
use FILL  FILL_5__2541_
timestamp 1701859473
transform -1 0 3330 0 1 2870
box -12 -8 32 272
use FILL  FILL_5__2542_
timestamp 1701859473
transform -1 0 2330 0 -1 6510
box -12 -8 32 272
use FILL  FILL_5__2543_
timestamp 1701859473
transform 1 0 890 0 1 4950
box -12 -8 32 272
use FILL  FILL_5__2544_
timestamp 1701859473
transform 1 0 1450 0 1 4430
box -12 -8 32 272
use FILL  FILL_5__2545_
timestamp 1701859473
transform 1 0 1310 0 -1 5470
box -12 -8 32 272
use FILL  FILL_5__2546_
timestamp 1701859473
transform -1 0 2050 0 -1 5470
box -12 -8 32 272
use FILL  FILL_5__2547_
timestamp 1701859473
transform 1 0 1990 0 -1 4430
box -12 -8 32 272
use FILL  FILL_5__2548_
timestamp 1701859473
transform 1 0 1110 0 1 4950
box -12 -8 32 272
use FILL  FILL_5__2549_
timestamp 1701859473
transform 1 0 1330 0 1 4950
box -12 -8 32 272
use FILL  FILL_5__2550_
timestamp 1701859473
transform -1 0 1810 0 -1 5470
box -12 -8 32 272
use FILL  FILL_5__2551_
timestamp 1701859473
transform 1 0 2590 0 -1 9630
box -12 -8 32 272
use FILL  FILL_5__2552_
timestamp 1701859473
transform 1 0 3430 0 -1 5470
box -12 -8 32 272
use FILL  FILL_5__2553_
timestamp 1701859473
transform -1 0 2810 0 -1 6510
box -12 -8 32 272
use FILL  FILL_5__2554_
timestamp 1701859473
transform -1 0 3270 0 1 6510
box -12 -8 32 272
use FILL  FILL_5__2555_
timestamp 1701859473
transform -1 0 3510 0 1 6510
box -12 -8 32 272
use FILL  FILL_5__2556_
timestamp 1701859473
transform -1 0 2830 0 1 6510
box -12 -8 32 272
use FILL  FILL_5__2557_
timestamp 1701859473
transform 1 0 2530 0 -1 6510
box -12 -8 32 272
use FILL  FILL_5__2558_
timestamp 1701859473
transform 1 0 3270 0 -1 7550
box -12 -8 32 272
use FILL  FILL_5__2559_
timestamp 1701859473
transform 1 0 3470 0 -1 7550
box -12 -8 32 272
use FILL  FILL_5__2560_
timestamp 1701859473
transform -1 0 3530 0 1 7030
box -12 -8 32 272
use FILL  FILL_5__2561_
timestamp 1701859473
transform -1 0 1550 0 1 4950
box -12 -8 32 272
use FILL  FILL_5__2562_
timestamp 1701859473
transform 1 0 3270 0 1 7030
box -12 -8 32 272
use FILL  FILL_5__2563_
timestamp 1701859473
transform 1 0 3830 0 1 5470
box -12 -8 32 272
use FILL  FILL_5__2564_
timestamp 1701859473
transform -1 0 3710 0 1 6510
box -12 -8 32 272
use FILL  FILL_5__2565_
timestamp 1701859473
transform 1 0 3770 0 1 7030
box -12 -8 32 272
use FILL  FILL_5__2566_
timestamp 1701859473
transform 1 0 3230 0 1 7550
box -12 -8 32 272
use FILL  FILL_5__2567_
timestamp 1701859473
transform 1 0 3190 0 -1 8070
box -12 -8 32 272
use FILL  FILL_5__2568_
timestamp 1701859473
transform -1 0 3010 0 -1 8590
box -12 -8 32 272
use FILL  FILL_5__2569_
timestamp 1701859473
transform 1 0 2770 0 -1 8590
box -12 -8 32 272
use FILL  FILL_5__2570_
timestamp 1701859473
transform 1 0 2950 0 -1 8070
box -12 -8 32 272
use FILL  FILL_5__2571_
timestamp 1701859473
transform -1 0 3910 0 -1 9630
box -12 -8 32 272
use FILL  FILL_5__2572_
timestamp 1701859473
transform -1 0 3930 0 -1 5990
box -12 -8 32 272
use FILL  FILL_5__2573_
timestamp 1701859473
transform -1 0 3790 0 -1 7030
box -12 -8 32 272
use FILL  FILL_5__2574_
timestamp 1701859473
transform 1 0 3510 0 -1 6510
box -12 -8 32 272
use FILL  FILL_5__2575_
timestamp 1701859473
transform 1 0 3410 0 -1 8070
box -12 -8 32 272
use FILL  FILL_5__2576_
timestamp 1701859473
transform -1 0 3450 0 -1 8590
box -12 -8 32 272
use FILL  FILL_5__2577_
timestamp 1701859473
transform 1 0 3330 0 1 9110
box -12 -8 32 272
use FILL  FILL_5__2578_
timestamp 1701859473
transform 1 0 3830 0 1 9110
box -12 -8 32 272
use FILL  FILL_5__2579_
timestamp 1701859473
transform -1 0 2810 0 -1 9630
box -12 -8 32 272
use FILL  FILL_5__2580_
timestamp 1701859473
transform -1 0 4170 0 -1 9110
box -12 -8 32 272
use FILL  FILL_5__2581_
timestamp 1701859473
transform -1 0 4090 0 1 9110
box -12 -8 32 272
use FILL  FILL_5__2582_
timestamp 1701859473
transform 1 0 3590 0 1 9110
box -12 -8 32 272
use FILL  FILL_5__2583_
timestamp 1701859473
transform 1 0 3090 0 1 9110
box -12 -8 32 272
use FILL  FILL_5__2584_
timestamp 1701859473
transform 1 0 2850 0 1 9110
box -12 -8 32 272
use FILL  FILL_5__2585_
timestamp 1701859473
transform 1 0 3950 0 -1 9110
box -12 -8 32 272
use FILL  FILL_5__2586_
timestamp 1701859473
transform 1 0 3110 0 1 9630
box -12 -8 32 272
use FILL  FILL_5__2587_
timestamp 1701859473
transform 1 0 3690 0 -1 9110
box -12 -8 32 272
use FILL  FILL_5__2588_
timestamp 1701859473
transform 1 0 3290 0 1 8590
box -12 -8 32 272
use FILL  FILL_5__2589_
timestamp 1701859473
transform 1 0 3130 0 -1 10150
box -12 -8 32 272
use FILL  FILL_5__2590_
timestamp 1701859473
transform 1 0 2870 0 -1 10150
box -12 -8 32 272
use FILL  FILL_5__2591_
timestamp 1701859473
transform -1 0 3630 0 -1 11190
box -12 -8 32 272
use FILL  FILL_5__2592_
timestamp 1701859473
transform -1 0 3690 0 -1 9630
box -12 -8 32 272
use FILL  FILL_5__2593_
timestamp 1701859473
transform -1 0 3210 0 -1 9630
box -12 -8 32 272
use FILL  FILL_5__2594_
timestamp 1701859473
transform -1 0 3370 0 -1 10150
box -12 -8 32 272
use FILL  FILL_5__2595_
timestamp 1701859473
transform 1 0 3090 0 -1 11190
box -12 -8 32 272
use FILL  FILL_5__2596_
timestamp 1701859473
transform 1 0 3370 0 -1 11190
box -12 -8 32 272
use FILL  FILL_5__2597_
timestamp 1701859473
transform 1 0 2830 0 -1 10670
box -12 -8 32 272
use FILL  FILL_5__2598_
timestamp 1701859473
transform -1 0 3570 0 1 9630
box -12 -8 32 272
use FILL  FILL_5__2599_
timestamp 1701859473
transform -1 0 3350 0 1 9630
box -12 -8 32 272
use FILL  FILL_5__2600_
timestamp 1701859473
transform -1 0 3070 0 1 10150
box -12 -8 32 272
use FILL  FILL_5__2601_
timestamp 1701859473
transform 1 0 3030 0 -1 10670
box -12 -8 32 272
use FILL  FILL_5__2602_
timestamp 1701859473
transform -1 0 3290 0 -1 10670
box -12 -8 32 272
use FILL  FILL_5__2603_
timestamp 1701859473
transform 1 0 3490 0 -1 10670
box -12 -8 32 272
use FILL  FILL_5__2604_
timestamp 1701859473
transform 1 0 3290 0 1 10150
box -12 -8 32 272
use FILL  FILL_5__2605_
timestamp 1701859473
transform 1 0 2410 0 1 10670
box -12 -8 32 272
use FILL  FILL_5__2606_
timestamp 1701859473
transform 1 0 2610 0 1 10670
box -12 -8 32 272
use FILL  FILL_5__2607_
timestamp 1701859473
transform -1 0 2850 0 1 10670
box -12 -8 32 272
use FILL  FILL_5__2608_
timestamp 1701859473
transform -1 0 3810 0 1 9630
box -12 -8 32 272
use FILL  FILL_5__2609_
timestamp 1701859473
transform -1 0 2430 0 1 9630
box -12 -8 32 272
use FILL  FILL_5__2610_
timestamp 1701859473
transform -1 0 2650 0 -1 10150
box -12 -8 32 272
use FILL  FILL_5__2611_
timestamp 1701859473
transform -1 0 2370 0 -1 10670
box -12 -8 32 272
use FILL  FILL_5__2612_
timestamp 1701859473
transform 1 0 2590 0 -1 10670
box -12 -8 32 272
use FILL  FILL_5__2613_
timestamp 1701859473
transform 1 0 1910 0 1 10670
box -12 -8 32 272
use FILL  FILL_5__2614_
timestamp 1701859473
transform 1 0 1910 0 -1 10670
box -12 -8 32 272
use FILL  FILL_5__2615_
timestamp 1701859473
transform -1 0 2430 0 -1 11190
box -12 -8 32 272
use FILL  FILL_5__2616_
timestamp 1701859473
transform -1 0 3450 0 -1 9630
box -12 -8 32 272
use FILL  FILL_5__2617_
timestamp 1701859473
transform 1 0 2350 0 -1 9630
box -12 -8 32 272
use FILL  FILL_5__2618_
timestamp 1701859473
transform -1 0 2630 0 1 10150
box -12 -8 32 272
use FILL  FILL_5__2619_
timestamp 1701859473
transform 1 0 2130 0 1 10670
box -12 -8 32 272
use FILL  FILL_5__2620_
timestamp 1701859473
transform 1 0 2170 0 -1 11190
box -12 -8 32 272
use FILL  FILL_5__2621_
timestamp 1701859473
transform -1 0 1450 0 1 5470
box -12 -8 32 272
use FILL  FILL_5__2622_
timestamp 1701859473
transform -1 0 1290 0 -1 5990
box -12 -8 32 272
use FILL  FILL_5__2623_
timestamp 1701859473
transform 1 0 2510 0 -1 5470
box -12 -8 32 272
use FILL  FILL_5__2624_
timestamp 1701859473
transform -1 0 2470 0 1 5470
box -12 -8 32 272
use FILL  FILL_5__2625_
timestamp 1701859473
transform 1 0 2270 0 -1 5470
box -12 -8 32 272
use FILL  FILL_5__2626_
timestamp 1701859473
transform -1 0 1010 0 -1 5470
box -12 -8 32 272
use FILL  FILL_5__2627_
timestamp 1701859473
transform -1 0 1530 0 1 3910
box -12 -8 32 272
use FILL  FILL_5__2628_
timestamp 1701859473
transform 1 0 1210 0 1 3910
box -12 -8 32 272
use FILL  FILL_5__2629_
timestamp 1701859473
transform -1 0 810 0 -1 5470
box -12 -8 32 272
use FILL  FILL_5__2630_
timestamp 1701859473
transform 1 0 790 0 -1 5990
box -12 -8 32 272
use FILL  FILL_5__2631_
timestamp 1701859473
transform -1 0 790 0 1 5990
box -12 -8 32 272
use FILL  FILL_5__2632_
timestamp 1701859473
transform 1 0 2170 0 1 10150
box -12 -8 32 272
use FILL  FILL_5__2633_
timestamp 1701859473
transform -1 0 2410 0 1 10150
box -12 -8 32 272
use FILL  FILL_5__2634_
timestamp 1701859473
transform 1 0 2370 0 -1 10150
box -12 -8 32 272
use FILL  FILL_5__2635_
timestamp 1701859473
transform 1 0 2150 0 -1 10150
box -12 -8 32 272
use FILL  FILL_5__2636_
timestamp 1701859473
transform -1 0 790 0 -1 10150
box -12 -8 32 272
use FILL  FILL_5__2637_
timestamp 1701859473
transform -1 0 590 0 1 6510
box -12 -8 32 272
use FILL  FILL_5__2638_
timestamp 1701859473
transform -1 0 370 0 1 6510
box -12 -8 32 272
use FILL  FILL_5__2639_
timestamp 1701859473
transform -1 0 350 0 -1 6510
box -12 -8 32 272
use FILL  FILL_5__2640_
timestamp 1701859473
transform -1 0 350 0 1 5990
box -12 -8 32 272
use FILL  FILL_5__2641_
timestamp 1701859473
transform 1 0 110 0 -1 7550
box -12 -8 32 272
use FILL  FILL_5__2642_
timestamp 1701859473
transform -1 0 450 0 1 4950
box -12 -8 32 272
use FILL  FILL_5__2643_
timestamp 1701859473
transform -1 0 2590 0 1 6510
box -12 -8 32 272
use FILL  FILL_5__2644_
timestamp 1701859473
transform 1 0 2630 0 -1 7030
box -12 -8 32 272
use FILL  FILL_5__2645_
timestamp 1701859473
transform 1 0 2810 0 1 7030
box -12 -8 32 272
use FILL  FILL_5__2646_
timestamp 1701859473
transform 1 0 2110 0 1 7030
box -12 -8 32 272
use FILL  FILL_5__2647_
timestamp 1701859473
transform 1 0 790 0 1 7550
box -12 -8 32 272
use FILL  FILL_5__2648_
timestamp 1701859473
transform 1 0 330 0 1 7550
box -12 -8 32 272
use FILL  FILL_5__2649_
timestamp 1701859473
transform 1 0 310 0 -1 7550
box -12 -8 32 272
use FILL  FILL_5__2650_
timestamp 1701859473
transform -1 0 790 0 -1 7550
box -12 -8 32 272
use FILL  FILL_5__2651_
timestamp 1701859473
transform 1 0 530 0 -1 7550
box -12 -8 32 272
use FILL  FILL_5__2652_
timestamp 1701859473
transform 1 0 530 0 1 7030
box -12 -8 32 272
use FILL  FILL_5__2653_
timestamp 1701859473
transform 1 0 110 0 1 7550
box -12 -8 32 272
use FILL  FILL_5__2654_
timestamp 1701859473
transform -1 0 590 0 1 7550
box -12 -8 32 272
use FILL  FILL_5__2655_
timestamp 1701859473
transform 1 0 1910 0 1 7030
box -12 -8 32 272
use FILL  FILL_5__2656_
timestamp 1701859473
transform 1 0 1550 0 -1 5470
box -12 -8 32 272
use FILL  FILL_5__2657_
timestamp 1701859473
transform -1 0 1750 0 1 5990
box -12 -8 32 272
use FILL  FILL_5__2658_
timestamp 1701859473
transform -1 0 2230 0 1 5470
box -12 -8 32 272
use FILL  FILL_5__2659_
timestamp 1701859473
transform 1 0 1990 0 -1 5990
box -12 -8 32 272
use FILL  FILL_5__2660_
timestamp 1701859473
transform -1 0 1990 0 1 5470
box -12 -8 32 272
use FILL  FILL_5__2661_
timestamp 1701859473
transform -1 0 1670 0 1 5470
box -12 -8 32 272
use FILL  FILL_5__2662_
timestamp 1701859473
transform 1 0 770 0 1 5470
box -12 -8 32 272
use FILL  FILL_5__2663_
timestamp 1701859473
transform -1 0 1050 0 -1 5990
box -12 -8 32 272
use FILL  FILL_5__2664_
timestamp 1701859473
transform 1 0 770 0 -1 7030
box -12 -8 32 272
use FILL  FILL_5__2665_
timestamp 1701859473
transform 1 0 1230 0 -1 7030
box -12 -8 32 272
use FILL  FILL_5__2666_
timestamp 1701859473
transform 1 0 1430 0 1 7030
box -12 -8 32 272
use FILL  FILL_5__2667_
timestamp 1701859473
transform 1 0 970 0 -1 7030
box -12 -8 32 272
use FILL  FILL_5__2668_
timestamp 1701859473
transform -1 0 2770 0 1 7550
box -12 -8 32 272
use FILL  FILL_5__2669_
timestamp 1701859473
transform 1 0 2710 0 -1 8070
box -12 -8 32 272
use FILL  FILL_5__2670_
timestamp 1701859473
transform 1 0 1970 0 -1 8070
box -12 -8 32 272
use FILL  FILL_5__2671_
timestamp 1701859473
transform -1 0 1470 0 1 7550
box -12 -8 32 272
use FILL  FILL_5__2672_
timestamp 1701859473
transform 1 0 1190 0 -1 7550
box -12 -8 32 272
use FILL  FILL_5__2673_
timestamp 1701859473
transform -1 0 1390 0 -1 7550
box -12 -8 32 272
use FILL  FILL_5__2674_
timestamp 1701859473
transform 1 0 1670 0 1 7030
box -12 -8 32 272
use FILL  FILL_5__2675_
timestamp 1701859473
transform 1 0 1610 0 -1 7550
box -12 -8 32 272
use FILL  FILL_5__2676_
timestamp 1701859473
transform -1 0 2050 0 -1 7550
box -12 -8 32 272
use FILL  FILL_5__2677_
timestamp 1701859473
transform 1 0 2450 0 -1 8070
box -12 -8 32 272
use FILL  FILL_5__2678_
timestamp 1701859473
transform -1 0 2230 0 -1 8070
box -12 -8 32 272
use FILL  FILL_5__2679_
timestamp 1701859473
transform -1 0 1670 0 1 8070
box -12 -8 32 272
use FILL  FILL_5__2680_
timestamp 1701859473
transform -1 0 350 0 -1 8590
box -12 -8 32 272
use FILL  FILL_5__2681_
timestamp 1701859473
transform 1 0 970 0 -1 7550
box -12 -8 32 272
use FILL  FILL_5__2682_
timestamp 1701859473
transform -1 0 350 0 -1 8070
box -12 -8 32 272
use FILL  FILL_5__2683_
timestamp 1701859473
transform -1 0 130 0 -1 9630
box -12 -8 32 272
use FILL  FILL_5__2684_
timestamp 1701859473
transform -1 0 130 0 1 10150
box -12 -8 32 272
use FILL  FILL_5__2685_
timestamp 1701859473
transform 1 0 1010 0 1 5990
box -12 -8 32 272
use FILL  FILL_5__2686_
timestamp 1701859473
transform 1 0 990 0 1 7550
box -12 -8 32 272
use FILL  FILL_5__2687_
timestamp 1701859473
transform -1 0 990 0 -1 10150
box -12 -8 32 272
use FILL  FILL_5__2688_
timestamp 1701859473
transform 1 0 110 0 -1 10150
box -12 -8 32 272
use FILL  FILL_5__2689_
timestamp 1701859473
transform 1 0 330 0 -1 9630
box -12 -8 32 272
use FILL  FILL_5__2690_
timestamp 1701859473
transform 1 0 330 0 1 9110
box -12 -8 32 272
use FILL  FILL_5__2691_
timestamp 1701859473
transform 1 0 2790 0 1 8590
box -12 -8 32 272
use FILL  FILL_5__2692_
timestamp 1701859473
transform 1 0 2550 0 1 8590
box -12 -8 32 272
use FILL  FILL_5__2693_
timestamp 1701859473
transform -1 0 1210 0 -1 9630
box -12 -8 32 272
use FILL  FILL_5__2694_
timestamp 1701859473
transform 1 0 790 0 -1 9630
box -12 -8 32 272
use FILL  FILL_5__2695_
timestamp 1701859473
transform 1 0 110 0 1 9630
box -12 -8 32 272
use FILL  FILL_5__2696_
timestamp 1701859473
transform -1 0 590 0 -1 10150
box -12 -8 32 272
use FILL  FILL_5__2697_
timestamp 1701859473
transform 1 0 330 0 -1 10150
box -12 -8 32 272
use FILL  FILL_5__2698_
timestamp 1701859473
transform 1 0 350 0 1 9630
box -12 -8 32 272
use FILL  FILL_5__2699_
timestamp 1701859473
transform 1 0 570 0 -1 9630
box -12 -8 32 272
use FILL  FILL_5__2700_
timestamp 1701859473
transform 1 0 590 0 1 9630
box -12 -8 32 272
use FILL  FILL_5__2701_
timestamp 1701859473
transform -1 0 810 0 -1 10670
box -12 -8 32 272
use FILL  FILL_5__2702_
timestamp 1701859473
transform 1 0 3530 0 1 8590
box -12 -8 32 272
use FILL  FILL_5__2703_
timestamp 1701859473
transform -1 0 3070 0 1 8590
box -12 -8 32 272
use FILL  FILL_5__2704_
timestamp 1701859473
transform -1 0 1550 0 1 9630
box -12 -8 32 272
use FILL  FILL_5__2705_
timestamp 1701859473
transform 1 0 1290 0 1 9630
box -12 -8 32 272
use FILL  FILL_5__2706_
timestamp 1701859473
transform 1 0 310 0 1 10150
box -12 -8 32 272
use FILL  FILL_5__2707_
timestamp 1701859473
transform -1 0 550 0 1 10150
box -12 -8 32 272
use FILL  FILL_5__2708_
timestamp 1701859473
transform 1 0 750 0 1 10150
box -12 -8 32 272
use FILL  FILL_5__2709_
timestamp 1701859473
transform -1 0 570 0 -1 10670
box -12 -8 32 272
use FILL  FILL_5__2710_
timestamp 1701859473
transform 1 0 1750 0 1 10150
box -12 -8 32 272
use FILL  FILL_5__2711_
timestamp 1701859473
transform 1 0 2290 0 1 8590
box -12 -8 32 272
use FILL  FILL_5__2712_
timestamp 1701859473
transform -1 0 2070 0 1 8590
box -12 -8 32 272
use FILL  FILL_5__2713_
timestamp 1701859473
transform -1 0 1930 0 -1 9630
box -12 -8 32 272
use FILL  FILL_5__2714_
timestamp 1701859473
transform 1 0 1690 0 -1 10150
box -12 -8 32 272
use FILL  FILL_5__2715_
timestamp 1701859473
transform 1 0 1010 0 1 10150
box -12 -8 32 272
use FILL  FILL_5__2716_
timestamp 1701859473
transform 1 0 1250 0 1 10150
box -12 -8 32 272
use FILL  FILL_5__2717_
timestamp 1701859473
transform 1 0 1510 0 1 10150
box -12 -8 32 272
use FILL  FILL_5__2718_
timestamp 1701859473
transform -1 0 10090 0 1 4950
box -12 -8 32 272
use FILL  FILL_5__2719_
timestamp 1701859473
transform -1 0 9850 0 1 4950
box -12 -8 32 272
use FILL  FILL_5__2720_
timestamp 1701859473
transform -1 0 4630 0 1 4950
box -12 -8 32 272
use FILL  FILL_5__2721_
timestamp 1701859473
transform -1 0 7390 0 -1 2350
box -12 -8 32 272
use FILL  FILL_5__2722_
timestamp 1701859473
transform 1 0 10030 0 -1 790
box -12 -8 32 272
use FILL  FILL_5__2723_
timestamp 1701859473
transform -1 0 7150 0 1 1830
box -12 -8 32 272
use FILL  FILL_5__2724_
timestamp 1701859473
transform -1 0 7150 0 -1 2350
box -12 -8 32 272
use FILL  FILL_5__2725_
timestamp 1701859473
transform 1 0 7010 0 1 3390
box -12 -8 32 272
use FILL  FILL_5__2726_
timestamp 1701859473
transform -1 0 7250 0 1 3390
box -12 -8 32 272
use FILL  FILL_5__2727_
timestamp 1701859473
transform -1 0 5470 0 1 3390
box -12 -8 32 272
use FILL  FILL_5__2728_
timestamp 1701859473
transform -1 0 5690 0 1 3390
box -12 -8 32 272
use FILL  FILL_5__2729_
timestamp 1701859473
transform -1 0 6790 0 -1 3910
box -12 -8 32 272
use FILL  FILL_5__2730_
timestamp 1701859473
transform 1 0 8290 0 -1 3910
box -12 -8 32 272
use FILL  FILL_5__2731_
timestamp 1701859473
transform 1 0 9310 0 1 1830
box -12 -8 32 272
use FILL  FILL_5__2732_
timestamp 1701859473
transform 1 0 7750 0 1 1830
box -12 -8 32 272
use FILL  FILL_5__2733_
timestamp 1701859473
transform 1 0 8630 0 1 2350
box -12 -8 32 272
use FILL  FILL_5__2734_
timestamp 1701859473
transform 1 0 7210 0 -1 5470
box -12 -8 32 272
use FILL  FILL_5__2735_
timestamp 1701859473
transform 1 0 7290 0 -1 2870
box -12 -8 32 272
use FILL  FILL_5__2736_
timestamp 1701859473
transform -1 0 7570 0 1 1310
box -12 -8 32 272
use FILL  FILL_5__2737_
timestamp 1701859473
transform 1 0 8630 0 1 1830
box -12 -8 32 272
use FILL  FILL_5__2738_
timestamp 1701859473
transform -1 0 8010 0 -1 2870
box -12 -8 32 272
use FILL  FILL_5__2739_
timestamp 1701859473
transform -1 0 7830 0 1 2870
box -12 -8 32 272
use FILL  FILL_5__2740_
timestamp 1701859473
transform -1 0 6610 0 -1 1830
box -12 -8 32 272
use FILL  FILL_5__2741_
timestamp 1701859473
transform 1 0 6810 0 -1 1830
box -12 -8 32 272
use FILL  FILL_5__2742_
timestamp 1701859473
transform -1 0 8250 0 -1 2870
box -12 -8 32 272
use FILL  FILL_5__2743_
timestamp 1701859473
transform -1 0 8270 0 1 2870
box -12 -8 32 272
use FILL  FILL_5__2744_
timestamp 1701859473
transform -1 0 7390 0 -1 270
box -12 -8 32 272
use FILL  FILL_5__2745_
timestamp 1701859473
transform -1 0 7350 0 1 1830
box -12 -8 32 272
use FILL  FILL_5__2746_
timestamp 1701859473
transform 1 0 8010 0 1 2870
box -12 -8 32 272
use FILL  FILL_5__2747_
timestamp 1701859473
transform -1 0 7810 0 -1 2350
box -12 -8 32 272
use FILL  FILL_5__2748_
timestamp 1701859473
transform 1 0 7990 0 -1 2350
box -12 -8 32 272
use FILL  FILL_5__2749_
timestamp 1701859473
transform 1 0 5950 0 1 1830
box -12 -8 32 272
use FILL  FILL_5__2750_
timestamp 1701859473
transform -1 0 6710 0 -1 1310
box -12 -8 32 272
use FILL  FILL_5__2751_
timestamp 1701859473
transform -1 0 6430 0 1 1830
box -12 -8 32 272
use FILL  FILL_5__2752_
timestamp 1701859473
transform -1 0 7790 0 1 2350
box -12 -8 32 272
use FILL  FILL_5__2753_
timestamp 1701859473
transform -1 0 7530 0 1 2350
box -12 -8 32 272
use FILL  FILL_5__2754_
timestamp 1701859473
transform 1 0 8870 0 -1 4950
box -12 -8 32 272
use FILL  FILL_5__2755_
timestamp 1701859473
transform 1 0 9770 0 1 790
box -12 -8 32 272
use FILL  FILL_5__2756_
timestamp 1701859473
transform -1 0 10010 0 1 790
box -12 -8 32 272
use FILL  FILL_5__2757_
timestamp 1701859473
transform 1 0 10710 0 -1 2870
box -12 -8 32 272
use FILL  FILL_5__2758_
timestamp 1701859473
transform -1 0 9210 0 -1 2870
box -12 -8 32 272
use FILL  FILL_5__2759_
timestamp 1701859473
transform 1 0 9130 0 1 4430
box -12 -8 32 272
use FILL  FILL_5__2760_
timestamp 1701859473
transform 1 0 10470 0 -1 790
box -12 -8 32 272
use FILL  FILL_5__2761_
timestamp 1701859473
transform 1 0 10230 0 -1 790
box -12 -8 32 272
use FILL  FILL_5__2762_
timestamp 1701859473
transform -1 0 10910 0 -1 1830
box -12 -8 32 272
use FILL  FILL_5__2763_
timestamp 1701859473
transform 1 0 6650 0 1 1830
box -12 -8 32 272
use FILL  FILL_5__2764_
timestamp 1701859473
transform -1 0 6910 0 1 1830
box -12 -8 32 272
use FILL  FILL_5__2765_
timestamp 1701859473
transform -1 0 10210 0 1 1830
box -12 -8 32 272
use FILL  FILL_5__2766_
timestamp 1701859473
transform -1 0 10030 0 -1 1830
box -12 -8 32 272
use FILL  FILL_5__2767_
timestamp 1701859473
transform -1 0 10450 0 -1 1830
box -12 -8 32 272
use FILL  FILL_5__2768_
timestamp 1701859473
transform -1 0 10430 0 1 1830
box -12 -8 32 272
use FILL  FILL_5__2769_
timestamp 1701859473
transform -1 0 10890 0 1 2350
box -12 -8 32 272
use FILL  FILL_5__2770_
timestamp 1701859473
transform -1 0 10670 0 -1 1830
box -12 -8 32 272
use FILL  FILL_5__2771_
timestamp 1701859473
transform 1 0 11090 0 1 2350
box -12 -8 32 272
use FILL  FILL_5__2772_
timestamp 1701859473
transform -1 0 10750 0 1 4950
box -12 -8 32 272
use FILL  FILL_5__2773_
timestamp 1701859473
transform 1 0 10490 0 -1 3910
box -12 -8 32 272
use FILL  FILL_5__2774_
timestamp 1701859473
transform -1 0 10790 0 -1 2350
box -12 -8 32 272
use FILL  FILL_5__2775_
timestamp 1701859473
transform -1 0 9150 0 -1 1310
box -12 -8 32 272
use FILL  FILL_5__2776_
timestamp 1701859473
transform 1 0 10690 0 -1 790
box -12 -8 32 272
use FILL  FILL_5__2777_
timestamp 1701859473
transform -1 0 8450 0 -1 270
box -12 -8 32 272
use FILL  FILL_5__2778_
timestamp 1701859473
transform 1 0 10990 0 1 270
box -12 -8 32 272
use FILL  FILL_5__2779_
timestamp 1701859473
transform 1 0 9070 0 -1 1830
box -12 -8 32 272
use FILL  FILL_5__2780_
timestamp 1701859473
transform -1 0 10090 0 1 1310
box -12 -8 32 272
use FILL  FILL_5__2781_
timestamp 1701859473
transform 1 0 10230 0 -1 1310
box -12 -8 32 272
use FILL  FILL_5__2782_
timestamp 1701859473
transform 1 0 8850 0 1 1830
box -12 -8 32 272
use FILL  FILL_5__2783_
timestamp 1701859473
transform 1 0 8410 0 -1 1310
box -12 -8 32 272
use FILL  FILL_5__2784_
timestamp 1701859473
transform 1 0 8650 0 -1 1310
box -12 -8 32 272
use FILL  FILL_5__2785_
timestamp 1701859473
transform 1 0 8870 0 -1 1830
box -12 -8 32 272
use FILL  FILL_5__2786_
timestamp 1701859473
transform -1 0 9350 0 -1 1310
box -12 -8 32 272
use FILL  FILL_5__2787_
timestamp 1701859473
transform -1 0 9550 0 -1 1830
box -12 -8 32 272
use FILL  FILL_5__2788_
timestamp 1701859473
transform 1 0 10230 0 -1 1830
box -12 -8 32 272
use FILL  FILL_5__2789_
timestamp 1701859473
transform 1 0 10310 0 1 1310
box -12 -8 32 272
use FILL  FILL_5__2790_
timestamp 1701859473
transform -1 0 10110 0 -1 2350
box -12 -8 32 272
use FILL  FILL_5__2791_
timestamp 1701859473
transform 1 0 9870 0 -1 2350
box -12 -8 32 272
use FILL  FILL_5__2792_
timestamp 1701859473
transform -1 0 10330 0 -1 2350
box -12 -8 32 272
use FILL  FILL_5__2793_
timestamp 1701859473
transform -1 0 10570 0 -1 2350
box -12 -8 32 272
use FILL  FILL_5__2794_
timestamp 1701859473
transform -1 0 10990 0 -1 2350
box -12 -8 32 272
use FILL  FILL_5__2795_
timestamp 1701859473
transform -1 0 10950 0 -1 2870
box -12 -8 32 272
use FILL  FILL_5__2796_
timestamp 1701859473
transform -1 0 10290 0 -1 2870
box -12 -8 32 272
use FILL  FILL_5__2797_
timestamp 1701859473
transform -1 0 9790 0 -1 1830
box -12 -8 32 272
use FILL  FILL_5__2798_
timestamp 1701859473
transform -1 0 10670 0 1 2350
box -12 -8 32 272
use FILL  FILL_5__2799_
timestamp 1701859473
transform 1 0 10450 0 -1 2870
box -12 -8 32 272
use FILL  FILL_5__2800_
timestamp 1701859473
transform -1 0 10470 0 -1 4430
box -12 -8 32 272
use FILL  FILL_5__2801_
timestamp 1701859473
transform -1 0 9430 0 -1 2870
box -12 -8 32 272
use FILL  FILL_5__2802_
timestamp 1701859473
transform -1 0 7290 0 -1 1830
box -12 -8 32 272
use FILL  FILL_5__2803_
timestamp 1701859473
transform 1 0 8490 0 -1 2870
box -12 -8 32 272
use FILL  FILL_5__2804_
timestamp 1701859473
transform -1 0 9550 0 -1 3390
box -12 -8 32 272
use FILL  FILL_5__2805_
timestamp 1701859473
transform -1 0 9850 0 -1 2870
box -12 -8 32 272
use FILL  FILL_5__2806_
timestamp 1701859473
transform 1 0 9610 0 -1 2870
box -12 -8 32 272
use FILL  FILL_5__2807_
timestamp 1701859473
transform 1 0 8950 0 -1 2350
box -12 -8 32 272
use FILL  FILL_5__2808_
timestamp 1701859473
transform 1 0 8710 0 -1 2350
box -12 -8 32 272
use FILL  FILL_5__2809_
timestamp 1701859473
transform 1 0 10430 0 1 2350
box -12 -8 32 272
use FILL  FILL_5__2810_
timestamp 1701859473
transform -1 0 10210 0 1 2350
box -12 -8 32 272
use FILL  FILL_5__2811_
timestamp 1701859473
transform 1 0 4990 0 -1 4430
box -12 -8 32 272
use FILL  FILL_5__2812_
timestamp 1701859473
transform -1 0 8950 0 1 4950
box -12 -8 32 272
use FILL  FILL_5__2813_
timestamp 1701859473
transform 1 0 9050 0 1 3390
box -12 -8 32 272
use FILL  FILL_5__2814_
timestamp 1701859473
transform -1 0 8870 0 -1 4430
box -12 -8 32 272
use FILL  FILL_5__2815_
timestamp 1701859473
transform -1 0 8650 0 1 3910
box -12 -8 32 272
use FILL  FILL_5__2816_
timestamp 1701859473
transform -1 0 8270 0 1 4950
box -12 -8 32 272
use FILL  FILL_5__2817_
timestamp 1701859473
transform 1 0 8710 0 1 4950
box -12 -8 32 272
use FILL  FILL_5__2818_
timestamp 1701859473
transform 1 0 8410 0 -1 4430
box -12 -8 32 272
use FILL  FILL_5__2819_
timestamp 1701859473
transform 1 0 8610 0 -1 4430
box -12 -8 32 272
use FILL  FILL_5__2820_
timestamp 1701859473
transform -1 0 9570 0 1 2350
box -12 -8 32 272
use FILL  FILL_5__2821_
timestamp 1701859473
transform 1 0 9090 0 1 2350
box -12 -8 32 272
use FILL  FILL_5__2822_
timestamp 1701859473
transform -1 0 9090 0 1 1830
box -12 -8 32 272
use FILL  FILL_5__2823_
timestamp 1701859473
transform -1 0 8870 0 1 2350
box -12 -8 32 272
use FILL  FILL_5__2824_
timestamp 1701859473
transform 1 0 9990 0 -1 3390
box -12 -8 32 272
use FILL  FILL_5__2825_
timestamp 1701859473
transform -1 0 10710 0 -1 3390
box -12 -8 32 272
use FILL  FILL_5__2826_
timestamp 1701859473
transform 1 0 9570 0 1 790
box -12 -8 32 272
use FILL  FILL_5__2827_
timestamp 1701859473
transform -1 0 9310 0 -1 1830
box -12 -8 32 272
use FILL  FILL_5__2828_
timestamp 1701859473
transform 1 0 7030 0 -1 1830
box -12 -8 32 272
use FILL  FILL_5__2829_
timestamp 1701859473
transform -1 0 10050 0 1 2870
box -12 -8 32 272
use FILL  FILL_5__2830_
timestamp 1701859473
transform 1 0 8350 0 -1 3390
box -12 -8 32 272
use FILL  FILL_5__2831_
timestamp 1701859473
transform 1 0 8390 0 1 3910
box -12 -8 32 272
use FILL  FILL_5__2832_
timestamp 1701859473
transform -1 0 9370 0 1 2350
box -12 -8 32 272
use FILL  FILL_5__2833_
timestamp 1701859473
transform -1 0 9310 0 -1 3390
box -12 -8 32 272
use FILL  FILL_5__2834_
timestamp 1701859473
transform -1 0 9070 0 -1 3390
box -12 -8 32 272
use FILL  FILL_5__2835_
timestamp 1701859473
transform -1 0 9370 0 1 790
box -12 -8 32 272
use FILL  FILL_5__2836_
timestamp 1701859473
transform 1 0 8950 0 1 1310
box -12 -8 32 272
use FILL  FILL_5__2837_
timestamp 1701859473
transform -1 0 9630 0 1 1310
box -12 -8 32 272
use FILL  FILL_5__2838_
timestamp 1701859473
transform -1 0 9750 0 1 3390
box -12 -8 32 272
use FILL  FILL_5__2839_
timestamp 1701859473
transform -1 0 9790 0 -1 3390
box -12 -8 32 272
use FILL  FILL_5__2840_
timestamp 1701859473
transform 1 0 9110 0 -1 270
box -12 -8 32 272
use FILL  FILL_5__2841_
timestamp 1701859473
transform -1 0 8910 0 -1 270
box -12 -8 32 272
use FILL  FILL_5__2842_
timestamp 1701859473
transform 1 0 9330 0 -1 270
box -12 -8 32 272
use FILL  FILL_5__2843_
timestamp 1701859473
transform 1 0 9570 0 -1 270
box -12 -8 32 272
use FILL  FILL_5__2844_
timestamp 1701859473
transform 1 0 9370 0 1 270
box -12 -8 32 272
use FILL  FILL_5__2845_
timestamp 1701859473
transform -1 0 10050 0 1 270
box -12 -8 32 272
use FILL  FILL_5__2846_
timestamp 1701859473
transform 1 0 9790 0 1 270
box -12 -8 32 272
use FILL  FILL_5__2847_
timestamp 1701859473
transform -1 0 11190 0 -1 10670
box -12 -8 32 272
use FILL  FILL_5__2848_
timestamp 1701859473
transform -1 0 10670 0 -1 1310
box -12 -8 32 272
use FILL  FILL_5__2849_
timestamp 1701859473
transform -1 0 11010 0 1 1310
box -12 -8 32 272
use FILL  FILL_5__2850_
timestamp 1701859473
transform -1 0 11150 0 -1 1830
box -12 -8 32 272
use FILL  FILL_5__2851_
timestamp 1701859473
transform 1 0 10750 0 -1 3910
box -12 -8 32 272
use FILL  FILL_5__2852_
timestamp 1701859473
transform -1 0 8950 0 1 270
box -12 -8 32 272
use FILL  FILL_5__2853_
timestamp 1701859473
transform -1 0 9170 0 1 270
box -12 -8 32 272
use FILL  FILL_5__2854_
timestamp 1701859473
transform 1 0 10670 0 1 790
box -12 -8 32 272
use FILL  FILL_5__2855_
timestamp 1701859473
transform -1 0 9870 0 1 1310
box -12 -8 32 272
use FILL  FILL_5__2856_
timestamp 1701859473
transform -1 0 10530 0 1 1310
box -12 -8 32 272
use FILL  FILL_5__2857_
timestamp 1701859473
transform -1 0 10770 0 1 1310
box -12 -8 32 272
use FILL  FILL_5__2858_
timestamp 1701859473
transform -1 0 11130 0 1 1830
box -12 -8 32 272
use FILL  FILL_5__2859_
timestamp 1701859473
transform 1 0 10990 0 -1 3910
box -12 -8 32 272
use FILL  FILL_5__2860_
timestamp 1701859473
transform 1 0 10910 0 -1 3390
box -12 -8 32 272
use FILL  FILL_5__2861_
timestamp 1701859473
transform 1 0 9790 0 -1 270
box -12 -8 32 272
use FILL  FILL_5__2862_
timestamp 1701859473
transform 1 0 8650 0 -1 270
box -12 -8 32 272
use FILL  FILL_5__2863_
timestamp 1701859473
transform -1 0 10290 0 1 270
box -12 -8 32 272
use FILL  FILL_5__2864_
timestamp 1701859473
transform 1 0 10530 0 1 270
box -12 -8 32 272
use FILL  FILL_5__2865_
timestamp 1701859473
transform -1 0 10770 0 1 270
box -12 -8 32 272
use FILL  FILL_5__2866_
timestamp 1701859473
transform -1 0 11150 0 -1 790
box -12 -8 32 272
use FILL  FILL_5__2867_
timestamp 1701859473
transform 1 0 11110 0 -1 3390
box -12 -8 32 272
use FILL  FILL_5__2868_
timestamp 1701859473
transform 1 0 11090 0 1 790
box -12 -8 32 272
use FILL  FILL_5__2869_
timestamp 1701859473
transform 1 0 10210 0 1 790
box -12 -8 32 272
use FILL  FILL_5__2870_
timestamp 1701859473
transform -1 0 10430 0 1 790
box -12 -8 32 272
use FILL  FILL_5__2871_
timestamp 1701859473
transform -1 0 10870 0 1 790
box -12 -8 32 272
use FILL  FILL_5__2872_
timestamp 1701859473
transform -1 0 11210 0 1 1310
box -12 -8 32 272
use FILL  FILL_5__2873_
timestamp 1701859473
transform -1 0 9990 0 1 3390
box -12 -8 32 272
use FILL  FILL_5__2874_
timestamp 1701859473
transform -1 0 10230 0 1 3390
box -12 -8 32 272
use FILL  FILL_5__2875_
timestamp 1701859473
transform -1 0 10810 0 -1 4950
box -12 -8 32 272
use FILL  FILL_5__2876_
timestamp 1701859473
transform -1 0 9770 0 1 1830
box -12 -8 32 272
use FILL  FILL_5__2877_
timestamp 1701859473
transform 1 0 9950 0 1 1830
box -12 -8 32 272
use FILL  FILL_5__2878_
timestamp 1701859473
transform 1 0 9770 0 -1 1310
box -12 -8 32 272
use FILL  FILL_5__2879_
timestamp 1701859473
transform -1 0 10010 0 -1 1310
box -12 -8 32 272
use FILL  FILL_5__2880_
timestamp 1701859473
transform 1 0 9510 0 1 1830
box -12 -8 32 272
use FILL  FILL_5__2881_
timestamp 1701859473
transform 1 0 10890 0 -1 790
box -12 -8 32 272
use FILL  FILL_5__2882_
timestamp 1701859473
transform -1 0 9570 0 -1 1310
box -12 -8 32 272
use FILL  FILL_5__2883_
timestamp 1701859473
transform -1 0 10470 0 -1 1310
box -12 -8 32 272
use FILL  FILL_5__2884_
timestamp 1701859473
transform 1 0 11110 0 -1 1310
box -12 -8 32 272
use FILL  FILL_5__2885_
timestamp 1701859473
transform -1 0 10890 0 -1 1310
box -12 -8 32 272
use FILL  FILL_5__2886_
timestamp 1701859473
transform 1 0 10650 0 1 1830
box -12 -8 32 272
use FILL  FILL_5__2887_
timestamp 1701859473
transform 1 0 10210 0 -1 4430
box -12 -8 32 272
use FILL  FILL_5__2888_
timestamp 1701859473
transform -1 0 4030 0 1 5470
box -12 -8 32 272
use FILL  FILL_5__2889_
timestamp 1701859473
transform 1 0 6150 0 1 2350
box -12 -8 32 272
use FILL  FILL_5__2890_
timestamp 1701859473
transform -1 0 8430 0 1 5990
box -12 -8 32 272
use FILL  FILL_5__2891_
timestamp 1701859473
transform -1 0 8230 0 1 5990
box -12 -8 32 272
use FILL  FILL_5__2892_
timestamp 1701859473
transform 1 0 7450 0 -1 5470
box -12 -8 32 272
use FILL  FILL_5__2893_
timestamp 1701859473
transform 1 0 7270 0 1 5470
box -12 -8 32 272
use FILL  FILL_5__2894_
timestamp 1701859473
transform 1 0 6550 0 -1 6510
box -12 -8 32 272
use FILL  FILL_5__2895_
timestamp 1701859473
transform 1 0 6690 0 1 6510
box -12 -8 32 272
use FILL  FILL_5__2896_
timestamp 1701859473
transform -1 0 7950 0 -1 5470
box -12 -8 32 272
use FILL  FILL_5__2897_
timestamp 1701859473
transform 1 0 7750 0 1 5470
box -12 -8 32 272
use FILL  FILL_5__2898_
timestamp 1701859473
transform 1 0 7270 0 -1 6510
box -12 -8 32 272
use FILL  FILL_5__2899_
timestamp 1701859473
transform 1 0 6790 0 -1 6510
box -12 -8 32 272
use FILL  FILL_5__2900_
timestamp 1701859473
transform -1 0 6330 0 -1 6510
box -12 -8 32 272
use FILL  FILL_5__2901_
timestamp 1701859473
transform 1 0 6070 0 -1 6510
box -12 -8 32 272
use FILL  FILL_5__2902_
timestamp 1701859473
transform -1 0 7990 0 1 5990
box -12 -8 32 272
use FILL  FILL_5__2903_
timestamp 1701859473
transform 1 0 7270 0 1 5990
box -12 -8 32 272
use FILL  FILL_5__2904_
timestamp 1701859473
transform 1 0 8390 0 -1 5470
box -12 -8 32 272
use FILL  FILL_5__2905_
timestamp 1701859473
transform 1 0 8410 0 1 5470
box -12 -8 32 272
use FILL  FILL_5__2906_
timestamp 1701859473
transform 1 0 8150 0 -1 5990
box -12 -8 32 272
use FILL  FILL_5__2907_
timestamp 1701859473
transform -1 0 7930 0 -1 5990
box -12 -8 32 272
use FILL  FILL_5__2908_
timestamp 1701859473
transform -1 0 8250 0 -1 4950
box -12 -8 32 272
use FILL  FILL_5__2909_
timestamp 1701859473
transform 1 0 3390 0 -1 4430
box -12 -8 32 272
use FILL  FILL_5__2910_
timestamp 1701859473
transform -1 0 6550 0 -1 4430
box -12 -8 32 272
use FILL  FILL_5__2911_
timestamp 1701859473
transform -1 0 6890 0 1 4430
box -12 -8 32 272
use FILL  FILL_5__2912_
timestamp 1701859473
transform 1 0 8670 0 -1 4950
box -12 -8 32 272
use FILL  FILL_5__2913_
timestamp 1701859473
transform -1 0 6850 0 -1 4950
box -12 -8 32 272
use FILL  FILL_5__2914_
timestamp 1701859473
transform 1 0 7110 0 -1 8070
box -12 -8 32 272
use FILL  FILL_5__2915_
timestamp 1701859473
transform 1 0 7230 0 -1 5990
box -12 -8 32 272
use FILL  FILL_5__2916_
timestamp 1701859473
transform 1 0 6990 0 -1 5990
box -12 -8 32 272
use FILL  FILL_5__2917_
timestamp 1701859473
transform -1 0 6370 0 -1 5990
box -12 -8 32 272
use FILL  FILL_5__2918_
timestamp 1701859473
transform 1 0 6290 0 1 5470
box -12 -8 32 272
use FILL  FILL_5__2919_
timestamp 1701859473
transform 1 0 6210 0 1 4950
box -12 -8 32 272
use FILL  FILL_5__2920_
timestamp 1701859473
transform 1 0 5970 0 1 4950
box -12 -8 32 272
use FILL  FILL_5__2921_
timestamp 1701859473
transform -1 0 7430 0 -1 3910
box -12 -8 32 272
use FILL  FILL_5__2922_
timestamp 1701859473
transform -1 0 7470 0 1 3910
box -12 -8 32 272
use FILL  FILL_5__2923_
timestamp 1701859473
transform -1 0 6790 0 -1 4430
box -12 -8 32 272
use FILL  FILL_5__2924_
timestamp 1701859473
transform 1 0 6410 0 1 4950
box -12 -8 32 272
use FILL  FILL_5__2925_
timestamp 1701859473
transform 1 0 7310 0 1 7550
box -12 -8 32 272
use FILL  FILL_5__2926_
timestamp 1701859473
transform -1 0 7550 0 1 4430
box -12 -8 32 272
use FILL  FILL_5__2927_
timestamp 1701859473
transform 1 0 7330 0 -1 4950
box -12 -8 32 272
use FILL  FILL_5__2928_
timestamp 1701859473
transform 1 0 7070 0 -1 4950
box -12 -8 32 272
use FILL  FILL_5__2929_
timestamp 1701859473
transform -1 0 6650 0 1 4950
box -12 -8 32 272
use FILL  FILL_5__2930_
timestamp 1701859473
transform 1 0 6190 0 1 1830
box -12 -8 32 272
use FILL  FILL_5__2931_
timestamp 1701859473
transform 1 0 7070 0 -1 2870
box -12 -8 32 272
use FILL  FILL_5__2932_
timestamp 1701859473
transform 1 0 5230 0 -1 4430
box -12 -8 32 272
use FILL  FILL_5__2933_
timestamp 1701859473
transform 1 0 5430 0 -1 4430
box -12 -8 32 272
use FILL  FILL_5__2934_
timestamp 1701859473
transform 1 0 5670 0 -1 4430
box -12 -8 32 272
use FILL  FILL_5__2935_
timestamp 1701859473
transform 1 0 6490 0 1 6510
box -12 -8 32 272
use FILL  FILL_5__2936_
timestamp 1701859473
transform 1 0 6370 0 -1 4950
box -12 -8 32 272
use FILL  FILL_5__2937_
timestamp 1701859473
transform 1 0 6590 0 -1 4950
box -12 -8 32 272
use FILL  FILL_5__2938_
timestamp 1701859473
transform 1 0 5070 0 1 4950
box -12 -8 32 272
use FILL  FILL_5__2939_
timestamp 1701859473
transform 1 0 4850 0 1 4950
box -12 -8 32 272
use FILL  FILL_5__2940_
timestamp 1701859473
transform -1 0 5910 0 -1 5470
box -12 -8 32 272
use FILL  FILL_5__2941_
timestamp 1701859473
transform 1 0 5670 0 -1 5470
box -12 -8 32 272
use FILL  FILL_5__2942_
timestamp 1701859473
transform -1 0 9370 0 1 4430
box -12 -8 32 272
use FILL  FILL_5__2943_
timestamp 1701859473
transform 1 0 6330 0 -1 4430
box -12 -8 32 272
use FILL  FILL_5__2944_
timestamp 1701859473
transform -1 0 6350 0 1 3910
box -12 -8 32 272
use FILL  FILL_5__2945_
timestamp 1701859473
transform -1 0 6430 0 1 4430
box -12 -8 32 272
use FILL  FILL_5__2946_
timestamp 1701859473
transform 1 0 6190 0 1 4430
box -12 -8 32 272
use FILL  FILL_5__2947_
timestamp 1701859473
transform -1 0 6590 0 -1 5990
box -12 -8 32 272
use FILL  FILL_5__2948_
timestamp 1701859473
transform 1 0 6130 0 -1 5990
box -12 -8 32 272
use FILL  FILL_5__2949_
timestamp 1701859473
transform -1 0 5950 0 -1 5990
box -12 -8 32 272
use FILL  FILL_5__2950_
timestamp 1701859473
transform 1 0 5810 0 1 5470
box -12 -8 32 272
use FILL  FILL_5__2951_
timestamp 1701859473
transform -1 0 6070 0 1 5470
box -12 -8 32 272
use FILL  FILL_5__2952_
timestamp 1701859473
transform -1 0 6150 0 -1 4950
box -12 -8 32 272
use FILL  FILL_5__2953_
timestamp 1701859473
transform -1 0 4430 0 1 4950
box -12 -8 32 272
use FILL  FILL_5__2954_
timestamp 1701859473
transform -1 0 6690 0 1 4430
box -12 -8 32 272
use FILL  FILL_5__2955_
timestamp 1701859473
transform -1 0 5970 0 1 4430
box -12 -8 32 272
use FILL  FILL_5__2956_
timestamp 1701859473
transform 1 0 5250 0 1 4430
box -12 -8 32 272
use FILL  FILL_5__2957_
timestamp 1701859473
transform 1 0 5190 0 -1 4950
box -12 -8 32 272
use FILL  FILL_5__2958_
timestamp 1701859473
transform -1 0 5510 0 1 4430
box -12 -8 32 272
use FILL  FILL_5__2959_
timestamp 1701859473
transform 1 0 7010 0 -1 5470
box -12 -8 32 272
use FILL  FILL_5__2960_
timestamp 1701859473
transform -1 0 6550 0 1 5470
box -12 -8 32 272
use FILL  FILL_5__2961_
timestamp 1701859473
transform 1 0 6310 0 -1 5470
box -12 -8 32 272
use FILL  FILL_5__2962_
timestamp 1701859473
transform -1 0 6570 0 -1 5470
box -12 -8 32 272
use FILL  FILL_5__2963_
timestamp 1701859473
transform -1 0 6810 0 -1 5470
box -12 -8 32 272
use FILL  FILL_5__2964_
timestamp 1701859473
transform -1 0 5450 0 -1 4950
box -12 -8 32 272
use FILL  FILL_5__2965_
timestamp 1701859473
transform 1 0 4950 0 -1 4950
box -12 -8 32 272
use FILL  FILL_5__2966_
timestamp 1701859473
transform -1 0 6410 0 1 2350
box -12 -8 32 272
use FILL  FILL_5__2967_
timestamp 1701859473
transform 1 0 7670 0 1 3910
box -12 -8 32 272
use FILL  FILL_5__2968_
timestamp 1701859473
transform -1 0 6990 0 -1 3910
box -12 -8 32 272
use FILL  FILL_5__2969_
timestamp 1701859473
transform -1 0 7210 0 -1 3910
box -12 -8 32 272
use FILL  FILL_5__2970_
timestamp 1701859473
transform -1 0 7250 0 1 3910
box -12 -8 32 272
use FILL  FILL_5__2971_
timestamp 1701859473
transform -1 0 6770 0 1 3910
box -12 -8 32 272
use FILL  FILL_5__2972_
timestamp 1701859473
transform 1 0 6990 0 1 3910
box -12 -8 32 272
use FILL  FILL_5__2973_
timestamp 1701859473
transform -1 0 7110 0 1 4430
box -12 -8 32 272
use FILL  FILL_5__2974_
timestamp 1701859473
transform 1 0 7010 0 -1 4430
box -12 -8 32 272
use FILL  FILL_5__2975_
timestamp 1701859473
transform -1 0 7770 0 -1 4430
box -12 -8 32 272
use FILL  FILL_5__2976_
timestamp 1701859473
transform -1 0 7530 0 -1 4430
box -12 -8 32 272
use FILL  FILL_5__2977_
timestamp 1701859473
transform 1 0 7250 0 -1 4430
box -12 -8 32 272
use FILL  FILL_5__2978_
timestamp 1701859473
transform 1 0 7310 0 1 4430
box -12 -8 32 272
use FILL  FILL_5__2979_
timestamp 1701859473
transform -1 0 3650 0 -1 4950
box -12 -8 32 272
use FILL  FILL_5__2980_
timestamp 1701859473
transform -1 0 3030 0 1 7550
box -12 -8 32 272
use FILL  FILL_5__2981_
timestamp 1701859473
transform 1 0 3550 0 1 4950
box -12 -8 32 272
use FILL  FILL_5__2982_
timestamp 1701859473
transform 1 0 9610 0 1 6510
box -12 -8 32 272
use FILL  FILL_5__2983_
timestamp 1701859473
transform 1 0 1930 0 1 4430
box -12 -8 32 272
use FILL  FILL_5__2984_
timestamp 1701859473
transform -1 0 3550 0 -1 3910
box -12 -8 32 272
use FILL  FILL_5__2985_
timestamp 1701859473
transform 1 0 3710 0 1 4430
box -12 -8 32 272
use FILL  FILL_5__2986_
timestamp 1701859473
transform -1 0 5910 0 -1 4430
box -12 -8 32 272
use FILL  FILL_5__2987_
timestamp 1701859473
transform -1 0 5730 0 1 4430
box -12 -8 32 272
use FILL  FILL_5__2988_
timestamp 1701859473
transform 1 0 9390 0 1 6510
box -12 -8 32 272
use FILL  FILL_5__2989_
timestamp 1701859473
transform 1 0 6010 0 1 6510
box -12 -8 32 272
use FILL  FILL_5__2990_
timestamp 1701859473
transform -1 0 6270 0 1 6510
box -12 -8 32 272
use FILL  FILL_5__2991_
timestamp 1701859473
transform 1 0 7170 0 1 6510
box -12 -8 32 272
use FILL  FILL_5__2992_
timestamp 1701859473
transform 1 0 9690 0 1 7030
box -12 -8 32 272
use FILL  FILL_5__2993_
timestamp 1701859473
transform 1 0 9890 0 1 7030
box -12 -8 32 272
use FILL  FILL_5__2994_
timestamp 1701859473
transform -1 0 10810 0 -1 7550
box -12 -8 32 272
use FILL  FILL_5__2995_
timestamp 1701859473
transform -1 0 7610 0 -1 7550
box -12 -8 32 272
use FILL  FILL_5__2996_
timestamp 1701859473
transform 1 0 7510 0 1 7550
box -12 -8 32 272
use FILL  FILL_5__2997_
timestamp 1701859473
transform -1 0 7390 0 -1 7550
box -12 -8 32 272
use FILL  FILL_5__2998_
timestamp 1701859473
transform -1 0 6450 0 -1 7550
box -12 -8 32 272
use FILL  FILL_5__2999_
timestamp 1701859473
transform 1 0 6170 0 1 7550
box -12 -8 32 272
use FILL  FILL_5__3000_
timestamp 1701859473
transform -1 0 6010 0 -1 7550
box -12 -8 32 272
use FILL  FILL_5__3001_
timestamp 1701859473
transform -1 0 5790 0 -1 7550
box -12 -8 32 272
use FILL  FILL_5__3002_
timestamp 1701859473
transform -1 0 6210 0 -1 7550
box -12 -8 32 272
use FILL  FILL_5__3003_
timestamp 1701859473
transform -1 0 6390 0 1 7550
box -12 -8 32 272
use FILL  FILL_5__3004_
timestamp 1701859473
transform 1 0 8190 0 1 7550
box -12 -8 32 272
use FILL  FILL_5__3005_
timestamp 1701859473
transform 1 0 11010 0 -1 7550
box -12 -8 32 272
use FILL  FILL_5__3006_
timestamp 1701859473
transform -1 0 10490 0 1 7550
box -12 -8 32 272
use FILL  FILL_5__3007_
timestamp 1701859473
transform 1 0 7010 0 1 7030
box -12 -8 32 272
use FILL  FILL_5__3008_
timestamp 1701859473
transform -1 0 6570 0 1 7030
box -12 -8 32 272
use FILL  FILL_5__3009_
timestamp 1701859473
transform -1 0 5970 0 -1 7030
box -12 -8 32 272
use FILL  FILL_5__3010_
timestamp 1701859473
transform 1 0 6190 0 -1 7030
box -12 -8 32 272
use FILL  FILL_5__3011_
timestamp 1701859473
transform 1 0 6770 0 1 7030
box -12 -8 32 272
use FILL  FILL_5__3012_
timestamp 1701859473
transform -1 0 7890 0 -1 7030
box -12 -8 32 272
use FILL  FILL_5__3013_
timestamp 1701859473
transform 1 0 8330 0 -1 7030
box -12 -8 32 272
use FILL  FILL_5__3014_
timestamp 1701859473
transform 1 0 10690 0 1 7550
box -12 -8 32 272
use FILL  FILL_5__3015_
timestamp 1701859473
transform -1 0 6410 0 -1 7030
box -12 -8 32 272
use FILL  FILL_5__3016_
timestamp 1701859473
transform -1 0 7290 0 1 7030
box -12 -8 32 272
use FILL  FILL_5__3017_
timestamp 1701859473
transform 1 0 6630 0 -1 7030
box -12 -8 32 272
use FILL  FILL_5__3018_
timestamp 1701859473
transform -1 0 6930 0 -1 7030
box -12 -8 32 272
use FILL  FILL_5__3019_
timestamp 1701859473
transform -1 0 7170 0 -1 7030
box -12 -8 32 272
use FILL  FILL_5__3020_
timestamp 1701859473
transform 1 0 8330 0 1 7030
box -12 -8 32 272
use FILL  FILL_5__3021_
timestamp 1701859473
transform -1 0 9390 0 -1 8070
box -12 -8 32 272
use FILL  FILL_5__3022_
timestamp 1701859473
transform 1 0 9570 0 -1 8070
box -12 -8 32 272
use FILL  FILL_5__3023_
timestamp 1701859473
transform -1 0 5790 0 1 6510
box -12 -8 32 272
use FILL  FILL_5__3024_
timestamp 1701859473
transform 1 0 5530 0 1 6510
box -12 -8 32 272
use FILL  FILL_5__3025_
timestamp 1701859473
transform -1 0 5550 0 -1 6510
box -12 -8 32 272
use FILL  FILL_5__3026_
timestamp 1701859473
transform 1 0 10970 0 -1 5990
box -12 -8 32 272
use FILL  FILL_5__3027_
timestamp 1701859473
transform -1 0 11210 0 -1 5990
box -12 -8 32 272
use FILL  FILL_5__3028_
timestamp 1701859473
transform -1 0 9830 0 -1 8070
box -12 -8 32 272
use FILL  FILL_5__3029_
timestamp 1701859473
transform -1 0 7150 0 -1 7550
box -12 -8 32 272
use FILL  FILL_5__3030_
timestamp 1701859473
transform -1 0 8130 0 -1 7030
box -12 -8 32 272
use FILL  FILL_5__3031_
timestamp 1701859473
transform 1 0 8110 0 1 7030
box -12 -8 32 272
use FILL  FILL_5__3032_
timestamp 1701859473
transform 1 0 7730 0 1 7550
box -12 -8 32 272
use FILL  FILL_5__3033_
timestamp 1701859473
transform -1 0 6810 0 1 8070
box -12 -8 32 272
use FILL  FILL_5__3034_
timestamp 1701859473
transform -1 0 7790 0 -1 8070
box -12 -8 32 272
use FILL  FILL_5__3035_
timestamp 1701859473
transform 1 0 7530 0 -1 8070
box -12 -8 32 272
use FILL  FILL_5__3036_
timestamp 1701859473
transform -1 0 7010 0 1 8070
box -12 -8 32 272
use FILL  FILL_5__3037_
timestamp 1701859473
transform -1 0 6570 0 1 8070
box -12 -8 32 272
use FILL  FILL_5__3038_
timestamp 1701859473
transform -1 0 7190 0 1 8070
box -12 -8 32 272
use FILL  FILL_5__3039_
timestamp 1701859473
transform 1 0 7410 0 1 8070
box -12 -8 32 272
use FILL  FILL_5__3040_
timestamp 1701859473
transform 1 0 9750 0 1 7550
box -12 -8 32 272
use FILL  FILL_5__3041_
timestamp 1701859473
transform -1 0 9610 0 -1 6510
box -12 -8 32 272
use FILL  FILL_5__3042_
timestamp 1701859473
transform 1 0 7310 0 -1 8070
box -12 -8 32 272
use FILL  FILL_5__3043_
timestamp 1701859473
transform -1 0 6630 0 1 7550
box -12 -8 32 272
use FILL  FILL_5__3044_
timestamp 1701859473
transform -1 0 6670 0 -1 7550
box -12 -8 32 272
use FILL  FILL_5__3045_
timestamp 1701859473
transform 1 0 6890 0 -1 7550
box -12 -8 32 272
use FILL  FILL_5__3046_
timestamp 1701859473
transform -1 0 7850 0 1 6510
box -12 -8 32 272
use FILL  FILL_5__3047_
timestamp 1701859473
transform 1 0 9190 0 1 6510
box -12 -8 32 272
use FILL  FILL_5__3048_
timestamp 1701859473
transform 1 0 9810 0 -1 6510
box -12 -8 32 272
use FILL  FILL_5__3049_
timestamp 1701859473
transform -1 0 6890 0 1 7550
box -12 -8 32 272
use FILL  FILL_5__3050_
timestamp 1701859473
transform -1 0 7110 0 1 7550
box -12 -8 32 272
use FILL  FILL_5__3051_
timestamp 1701859473
transform -1 0 7850 0 1 7030
box -12 -8 32 272
use FILL  FILL_5__3052_
timestamp 1701859473
transform 1 0 7550 0 1 7030
box -12 -8 32 272
use FILL  FILL_5__3053_
timestamp 1701859473
transform 1 0 7390 0 -1 7030
box -12 -8 32 272
use FILL  FILL_5__3054_
timestamp 1701859473
transform -1 0 7650 0 -1 7030
box -12 -8 32 272
use FILL  FILL_5__3055_
timestamp 1701859473
transform 1 0 8070 0 1 6510
box -12 -8 32 272
use FILL  FILL_5__3056_
timestamp 1701859473
transform -1 0 9590 0 1 5470
box -12 -8 32 272
use FILL  FILL_5__3057_
timestamp 1701859473
transform -1 0 9350 0 1 5470
box -12 -8 32 272
use FILL  FILL_5__3058_
timestamp 1701859473
transform 1 0 8770 0 -1 7550
box -12 -8 32 272
use FILL  FILL_5__3059_
timestamp 1701859473
transform -1 0 8650 0 -1 5990
box -12 -8 32 272
use FILL  FILL_5__3060_
timestamp 1701859473
transform 1 0 9830 0 1 6510
box -12 -8 32 272
use FILL  FILL_5__3061_
timestamp 1701859473
transform 1 0 10070 0 1 6510
box -12 -8 32 272
use FILL  FILL_5__3062_
timestamp 1701859473
transform -1 0 9690 0 -1 7550
box -12 -8 32 272
use FILL  FILL_5__3063_
timestamp 1701859473
transform 1 0 9430 0 -1 7550
box -12 -8 32 272
use FILL  FILL_5__3064_
timestamp 1701859473
transform -1 0 10390 0 -1 7030
box -12 -8 32 272
use FILL  FILL_5__3065_
timestamp 1701859473
transform -1 0 10630 0 -1 7030
box -12 -8 32 272
use FILL  FILL_5__3066_
timestamp 1701859473
transform -1 0 8550 0 -1 7550
box -12 -8 32 272
use FILL  FILL_5__3067_
timestamp 1701859473
transform 1 0 8290 0 -1 7550
box -12 -8 32 272
use FILL  FILL_5__3068_
timestamp 1701859473
transform 1 0 10250 0 -1 5990
box -12 -8 32 272
use FILL  FILL_5__3069_
timestamp 1701859473
transform 1 0 10490 0 -1 5990
box -12 -8 32 272
use FILL  FILL_5__3070_
timestamp 1701859473
transform 1 0 8950 0 -1 7550
box -12 -8 32 272
use FILL  FILL_5__3071_
timestamp 1701859473
transform -1 0 9210 0 -1 7550
box -12 -8 32 272
use FILL  FILL_5__3072_
timestamp 1701859473
transform -1 0 9830 0 1 5990
box -12 -8 32 272
use FILL  FILL_5__3073_
timestamp 1701859473
transform -1 0 10050 0 1 5990
box -12 -8 32 272
use FILL  FILL_5__3074_
timestamp 1701859473
transform 1 0 8870 0 1 5990
box -12 -8 32 272
use FILL  FILL_5__3075_
timestamp 1701859473
transform 1 0 8870 0 -1 5990
box -12 -8 32 272
use FILL  FILL_5__3076_
timestamp 1701859473
transform 1 0 10770 0 1 6510
box -12 -8 32 272
use FILL  FILL_5__3077_
timestamp 1701859473
transform 1 0 10970 0 1 6510
box -12 -8 32 272
use FILL  FILL_5__3078_
timestamp 1701859473
transform -1 0 8770 0 -1 7030
box -12 -8 32 272
use FILL  FILL_5__3079_
timestamp 1701859473
transform -1 0 8550 0 -1 7030
box -12 -8 32 272
use FILL  FILL_5__3080_
timestamp 1701859473
transform 1 0 11030 0 -1 8590
box -12 -8 32 272
use FILL  FILL_5__3081_
timestamp 1701859473
transform -1 0 11030 0 -1 270
box -12 -8 32 272
use FILL  FILL_5__3082_
timestamp 1701859473
transform 1 0 10130 0 -1 8590
box -12 -8 32 272
use FILL  FILL_5__3083_
timestamp 1701859473
transform -1 0 9910 0 -1 8590
box -12 -8 32 272
use FILL  FILL_5__3084_
timestamp 1701859473
transform -1 0 9090 0 1 7550
box -12 -8 32 272
use FILL  FILL_5__3085_
timestamp 1701859473
transform 1 0 8990 0 1 7030
box -12 -8 32 272
use FILL  FILL_5__3086_
timestamp 1701859473
transform -1 0 10750 0 1 5990
box -12 -8 32 272
use FILL  FILL_5__3087_
timestamp 1701859473
transform 1 0 10950 0 1 5990
box -12 -8 32 272
use FILL  FILL_5__3088_
timestamp 1701859473
transform 1 0 8310 0 1 8070
box -12 -8 32 272
use FILL  FILL_5__3089_
timestamp 1701859473
transform -1 0 8090 0 1 8070
box -12 -8 32 272
use FILL  FILL_5__3090_
timestamp 1701859473
transform -1 0 11190 0 1 4950
box -12 -8 32 272
use FILL  FILL_5__3091_
timestamp 1701859473
transform 1 0 10930 0 1 4950
box -12 -8 32 272
use FILL  FILL_5__3092_
timestamp 1701859473
transform 1 0 8850 0 -1 5470
box -12 -8 32 272
use FILL  FILL_5__3093_
timestamp 1701859473
transform -1 0 9090 0 -1 5470
box -12 -8 32 272
use FILL  FILL_5__3094_
timestamp 1701859473
transform -1 0 10290 0 -1 5470
box -12 -8 32 272
use FILL  FILL_5__3095_
timestamp 1701859473
transform 1 0 10230 0 1 5470
box -12 -8 32 272
use FILL  FILL_5__3096_
timestamp 1701859473
transform 1 0 8970 0 1 6510
box -12 -8 32 272
use FILL  FILL_5__3097_
timestamp 1701859473
transform -1 0 8750 0 1 6510
box -12 -8 32 272
use FILL  FILL_5__3098_
timestamp 1701859473
transform -1 0 10450 0 1 8070
box -12 -8 32 272
use FILL  FILL_5__3099_
timestamp 1701859473
transform -1 0 11210 0 -1 8070
box -12 -8 32 272
use FILL  FILL_5__3100_
timestamp 1701859473
transform 1 0 10210 0 1 8070
box -12 -8 32 272
use FILL  FILL_5__3101_
timestamp 1701859473
transform 1 0 10350 0 -1 8590
box -12 -8 32 272
use FILL  FILL_5__3102_
timestamp 1701859473
transform 1 0 8430 0 -1 8070
box -12 -8 32 272
use FILL  FILL_5__3103_
timestamp 1701859473
transform -1 0 8410 0 1 7550
box -12 -8 32 272
use FILL  FILL_5__3104_
timestamp 1701859473
transform -1 0 11210 0 1 6510
box -12 -8 32 272
use FILL  FILL_5__3105_
timestamp 1701859473
transform -1 0 11010 0 -1 4950
box -12 -8 32 272
use FILL  FILL_5__3106_
timestamp 1701859473
transform 1 0 9430 0 -1 8590
box -12 -8 32 272
use FILL  FILL_5__3107_
timestamp 1701859473
transform -1 0 9670 0 -1 8590
box -12 -8 32 272
use FILL  FILL_5__3108_
timestamp 1701859473
transform 1 0 10030 0 1 5470
box -12 -8 32 272
use FILL  FILL_5__3109_
timestamp 1701859473
transform -1 0 9810 0 1 5470
box -12 -8 32 272
use FILL  FILL_5__3110_
timestamp 1701859473
transform 1 0 8450 0 -1 6510
box -12 -8 32 272
use FILL  FILL_5__3111_
timestamp 1701859473
transform -1 0 8230 0 -1 6510
box -12 -8 32 272
use FILL  FILL_5__3112_
timestamp 1701859473
transform 1 0 570 0 -1 2870
box -12 -8 32 272
use FILL  FILL_5__3113_
timestamp 1701859473
transform 1 0 110 0 -1 2870
box -12 -8 32 272
use FILL  FILL_5__3114_
timestamp 1701859473
transform -1 0 370 0 -1 2870
box -12 -8 32 272
use FILL  FILL_5__3115_
timestamp 1701859473
transform -1 0 1250 0 1 2350
box -12 -8 32 272
use FILL  FILL_5__3116_
timestamp 1701859473
transform 1 0 1010 0 -1 2350
box -12 -8 32 272
use FILL  FILL_5__3117_
timestamp 1701859473
transform 1 0 2090 0 -1 1310
box -12 -8 32 272
use FILL  FILL_5__3118_
timestamp 1701859473
transform -1 0 1470 0 -1 2350
box -12 -8 32 272
use FILL  FILL_5__3119_
timestamp 1701859473
transform -1 0 1230 0 -1 2350
box -12 -8 32 272
use FILL  FILL_5__3120_
timestamp 1701859473
transform -1 0 530 0 1 2350
box -12 -8 32 272
use FILL  FILL_5__3121_
timestamp 1701859473
transform 1 0 310 0 1 2870
box -12 -8 32 272
use FILL  FILL_5__3122_
timestamp 1701859473
transform 1 0 2570 0 -1 3390
box -12 -8 32 272
use FILL  FILL_5__3123_
timestamp 1701859473
transform 1 0 590 0 1 3390
box -12 -8 32 272
use FILL  FILL_5__3124_
timestamp 1701859473
transform -1 0 370 0 1 3390
box -12 -8 32 272
use FILL  FILL_5__3125_
timestamp 1701859473
transform -1 0 790 0 -1 2350
box -12 -8 32 272
use FILL  FILL_5__3126_
timestamp 1701859473
transform -1 0 1490 0 1 2350
box -12 -8 32 272
use FILL  FILL_5__3127_
timestamp 1701859473
transform -1 0 1010 0 1 2350
box -12 -8 32 272
use FILL  FILL_5__3128_
timestamp 1701859473
transform -1 0 1950 0 1 2350
box -12 -8 32 272
use FILL  FILL_5__3129_
timestamp 1701859473
transform -1 0 1710 0 -1 2350
box -12 -8 32 272
use FILL  FILL_5__3130_
timestamp 1701859473
transform -1 0 1730 0 1 2350
box -12 -8 32 272
use FILL  FILL_5__3131_
timestamp 1701859473
transform -1 0 770 0 1 2350
box -12 -8 32 272
use FILL  FILL_5__3132_
timestamp 1701859473
transform 1 0 530 0 1 2870
box -12 -8 32 272
use FILL  FILL_5__3133_
timestamp 1701859473
transform 1 0 590 0 -1 3910
box -12 -8 32 272
use FILL  FILL_5__3134_
timestamp 1701859473
transform -1 0 1270 0 1 3390
box -12 -8 32 272
use FILL  FILL_5__3135_
timestamp 1701859473
transform 1 0 1030 0 1 3390
box -12 -8 32 272
use FILL  FILL_5__3136_
timestamp 1701859473
transform -1 0 610 0 -1 3390
box -12 -8 32 272
use FILL  FILL_5__3137_
timestamp 1701859473
transform 1 0 330 0 -1 3390
box -12 -8 32 272
use FILL  FILL_5__3138_
timestamp 1701859473
transform -1 0 1730 0 1 4430
box -12 -8 32 272
use FILL  FILL_5__3139_
timestamp 1701859473
transform -1 0 1930 0 -1 3390
box -12 -8 32 272
use FILL  FILL_5__3140_
timestamp 1701859473
transform -1 0 350 0 1 3910
box -12 -8 32 272
use FILL  FILL_5__3141_
timestamp 1701859473
transform 1 0 790 0 1 4430
box -12 -8 32 272
use FILL  FILL_5__3142_
timestamp 1701859473
transform 1 0 1030 0 1 4430
box -12 -8 32 272
use FILL  FILL_5__3143_
timestamp 1701859473
transform 1 0 1050 0 -1 4430
box -12 -8 32 272
use FILL  FILL_5__3144_
timestamp 1701859473
transform -1 0 1290 0 -1 4430
box -12 -8 32 272
use FILL  FILL_5__3145_
timestamp 1701859473
transform -1 0 570 0 1 3910
box -12 -8 32 272
use FILL  FILL_5__3146_
timestamp 1701859473
transform -1 0 790 0 1 3910
box -12 -8 32 272
use FILL  FILL_5__3147_
timestamp 1701859473
transform 1 0 570 0 -1 4430
box -12 -8 32 272
use FILL  FILL_5__3148_
timestamp 1701859473
transform -1 0 830 0 -1 4430
box -12 -8 32 272
use FILL  FILL_5__3149_
timestamp 1701859473
transform -1 0 130 0 -1 3910
box -12 -8 32 272
use FILL  FILL_5__3150_
timestamp 1701859473
transform -1 0 990 0 1 3910
box -12 -8 32 272
use FILL  FILL_5__3151_
timestamp 1701859473
transform 1 0 110 0 1 3910
box -12 -8 32 272
use FILL  FILL_5__3152_
timestamp 1701859473
transform 1 0 110 0 -1 4430
box -12 -8 32 272
use FILL  FILL_5__3153_
timestamp 1701859473
transform -1 0 350 0 -1 4430
box -12 -8 32 272
use FILL  FILL_5__3154_
timestamp 1701859473
transform -1 0 850 0 -1 3390
box -12 -8 32 272
use FILL  FILL_5__3155_
timestamp 1701859473
transform -1 0 130 0 1 2870
box -12 -8 32 272
use FILL  FILL_5__3156_
timestamp 1701859473
transform 1 0 110 0 -1 3390
box -12 -8 32 272
use FILL  FILL_5__3157_
timestamp 1701859473
transform -1 0 130 0 1 3390
box -12 -8 32 272
use FILL  FILL_5__3158_
timestamp 1701859473
transform 1 0 110 0 1 4430
box -12 -8 32 272
use FILL  FILL_5__3159_
timestamp 1701859473
transform 1 0 330 0 1 4430
box -12 -8 32 272
use FILL  FILL_5__3160_
timestamp 1701859473
transform -1 0 570 0 1 4430
box -12 -8 32 272
use FILL  FILL_5__3161_
timestamp 1701859473
transform 1 0 4210 0 -1 7030
box -12 -8 32 272
use FILL  FILL_5__3162_
timestamp 1701859473
transform -1 0 4450 0 -1 7030
box -12 -8 32 272
use FILL  FILL_5__3163_
timestamp 1701859473
transform 1 0 4670 0 -1 7030
box -12 -8 32 272
use FILL  FILL_5__3164_
timestamp 1701859473
transform 1 0 4910 0 1 7030
box -12 -8 32 272
use FILL  FILL_5__3165_
timestamp 1701859473
transform 1 0 4170 0 1 7550
box -12 -8 32 272
use FILL  FILL_5__3166_
timestamp 1701859473
transform -1 0 4410 0 1 7550
box -12 -8 32 272
use FILL  FILL_5__3167_
timestamp 1701859473
transform 1 0 4890 0 -1 10150
box -12 -8 32 272
use FILL  FILL_5__3168_
timestamp 1701859473
transform 1 0 5090 0 -1 10150
box -12 -8 32 272
use FILL  FILL_5__3169_
timestamp 1701859473
transform -1 0 3730 0 -1 10670
box -12 -8 32 272
use FILL  FILL_5__3170_
timestamp 1701859473
transform -1 0 3950 0 -1 10670
box -12 -8 32 272
use FILL  FILL_5__3171_
timestamp 1701859473
transform 1 0 4370 0 -1 10670
box -12 -8 32 272
use FILL  FILL_5__3172_
timestamp 1701859473
transform -1 0 4610 0 -1 10670
box -12 -8 32 272
use FILL  FILL_5__3173_
timestamp 1701859473
transform 1 0 4210 0 1 10150
box -12 -8 32 272
use FILL  FILL_5__3174_
timestamp 1701859473
transform -1 0 4450 0 1 10150
box -12 -8 32 272
use FILL  FILL_5__3175_
timestamp 1701859473
transform 1 0 5550 0 1 10150
box -12 -8 32 272
use FILL  FILL_5__3176_
timestamp 1701859473
transform 1 0 5310 0 1 10150
box -12 -8 32 272
use FILL  FILL_5__3177_
timestamp 1701859473
transform -1 0 1790 0 -1 5990
box -12 -8 32 272
use FILL  FILL_5__3178_
timestamp 1701859473
transform 1 0 2230 0 -1 5990
box -12 -8 32 272
use FILL  FILL_5__3179_
timestamp 1701859473
transform -1 0 1510 0 1 6510
box -12 -8 32 272
use FILL  FILL_5__3180_
timestamp 1701859473
transform -1 0 1730 0 1 6510
box -12 -8 32 272
use FILL  FILL_5__3181_
timestamp 1701859473
transform -1 0 590 0 -1 6510
box -12 -8 32 272
use FILL  FILL_5__3182_
timestamp 1701859473
transform -1 0 990 0 -1 6510
box -12 -8 32 272
use FILL  FILL_5__3183_
timestamp 1701859473
transform 1 0 350 0 1 8070
box -12 -8 32 272
use FILL  FILL_5__3184_
timestamp 1701859473
transform -1 0 590 0 1 8070
box -12 -8 32 272
use FILL  FILL_5__3185_
timestamp 1701859473
transform -1 0 130 0 -1 8590
box -12 -8 32 272
use FILL  FILL_5__3186_
timestamp 1701859473
transform -1 0 130 0 1 8070
box -12 -8 32 272
use FILL  FILL_5__3187_
timestamp 1701859473
transform 1 0 750 0 -1 9110
box -12 -8 32 272
use FILL  FILL_5__3188_
timestamp 1701859473
transform 1 0 970 0 -1 9110
box -12 -8 32 272
use FILL  FILL_5__3189_
timestamp 1701859473
transform 1 0 2150 0 -1 9630
box -12 -8 32 272
use FILL  FILL_5__3190_
timestamp 1701859473
transform 1 0 2390 0 1 9110
box -12 -8 32 272
use FILL  FILL_5__3191_
timestamp 1701859473
transform 1 0 1450 0 -1 9110
box -12 -8 32 272
use FILL  FILL_5__3192_
timestamp 1701859473
transform -1 0 1690 0 -1 9110
box -12 -8 32 272
use FILL  FILL_5__3324_
timestamp 1701859473
transform 1 0 5630 0 1 8070
box -12 -8 32 272
use FILL  FILL_5__3325_
timestamp 1701859473
transform -1 0 6350 0 1 8070
box -12 -8 32 272
use FILL  FILL_5__3326_
timestamp 1701859473
transform -1 0 6250 0 -1 8070
box -12 -8 32 272
use FILL  FILL_5__3327_
timestamp 1701859473
transform -1 0 6210 0 -1 8590
box -12 -8 32 272
use FILL  FILL_5__3328_
timestamp 1701859473
transform -1 0 6110 0 1 8070
box -12 -8 32 272
use FILL  FILL_5__3329_
timestamp 1701859473
transform 1 0 5870 0 1 8070
box -12 -8 32 272
use FILL  FILL_5__3330_
timestamp 1701859473
transform -1 0 7050 0 1 8590
box -12 -8 32 272
use FILL  FILL_5__3331_
timestamp 1701859473
transform 1 0 7330 0 -1 8590
box -12 -8 32 272
use FILL  FILL_5__3332_
timestamp 1701859473
transform 1 0 7050 0 -1 8590
box -12 -8 32 272
use FILL  FILL_5__3333_
timestamp 1701859473
transform 1 0 10250 0 1 8590
box -12 -8 32 272
use FILL  FILL_5__3334_
timestamp 1701859473
transform 1 0 9370 0 1 8590
box -12 -8 32 272
use FILL  FILL_5__3335_
timestamp 1701859473
transform 1 0 7910 0 -1 10150
box -12 -8 32 272
use FILL  FILL_5__3336_
timestamp 1701859473
transform -1 0 6750 0 1 9630
box -12 -8 32 272
use FILL  FILL_5__3337_
timestamp 1701859473
transform -1 0 6270 0 1 9630
box -12 -8 32 272
use FILL  FILL_5__3338_
timestamp 1701859473
transform 1 0 7230 0 -1 10150
box -12 -8 32 272
use FILL  FILL_5__3339_
timestamp 1701859473
transform -1 0 8110 0 1 10150
box -12 -8 32 272
use FILL  FILL_5__3340_
timestamp 1701859473
transform 1 0 7870 0 1 10150
box -12 -8 32 272
use FILL  FILL_5__3341_
timestamp 1701859473
transform 1 0 7630 0 1 10150
box -12 -8 32 272
use FILL  FILL_5__3342_
timestamp 1701859473
transform 1 0 6850 0 -1 11190
box -12 -8 32 272
use FILL  FILL_5__3343_
timestamp 1701859473
transform -1 0 7450 0 -1 10150
box -12 -8 32 272
use FILL  FILL_5__3344_
timestamp 1701859473
transform 1 0 7670 0 -1 10150
box -12 -8 32 272
use FILL  FILL_5__3345_
timestamp 1701859473
transform -1 0 9050 0 1 9630
box -12 -8 32 272
use FILL  FILL_5__3346_
timestamp 1701859473
transform 1 0 8570 0 1 10150
box -12 -8 32 272
use FILL  FILL_5__3347_
timestamp 1701859473
transform -1 0 8350 0 1 10150
box -12 -8 32 272
use FILL  FILL_5__3348_
timestamp 1701859473
transform 1 0 9170 0 -1 10670
box -12 -8 32 272
use FILL  FILL_5__3349_
timestamp 1701859473
transform 1 0 7910 0 1 9630
box -12 -8 32 272
use FILL  FILL_5__3350_
timestamp 1701859473
transform 1 0 7610 0 -1 8590
box -12 -8 32 272
use FILL  FILL_5__3351_
timestamp 1701859473
transform -1 0 7790 0 1 8590
box -12 -8 32 272
use FILL  FILL_5__3352_
timestamp 1701859473
transform -1 0 8250 0 -1 9110
box -12 -8 32 272
use FILL  FILL_5__3353_
timestamp 1701859473
transform 1 0 8130 0 -1 10150
box -12 -8 32 272
use FILL  FILL_5__3354_
timestamp 1701859473
transform 1 0 7810 0 -1 10670
box -12 -8 32 272
use FILL  FILL_5__3355_
timestamp 1701859473
transform -1 0 7590 0 -1 10670
box -12 -8 32 272
use FILL  FILL_5__3356_
timestamp 1701859473
transform 1 0 7370 0 -1 10670
box -12 -8 32 272
use FILL  FILL_5__3357_
timestamp 1701859473
transform 1 0 7190 0 1 10670
box -12 -8 32 272
use FILL  FILL_5__3358_
timestamp 1701859473
transform 1 0 7450 0 1 10670
box -12 -8 32 272
use FILL  FILL_5__3359_
timestamp 1701859473
transform 1 0 7690 0 1 10670
box -12 -8 32 272
use FILL  FILL_5__3360_
timestamp 1701859473
transform -1 0 7950 0 1 10670
box -12 -8 32 272
use FILL  FILL_5__3361_
timestamp 1701859473
transform 1 0 8970 0 -1 10670
box -12 -8 32 272
use FILL  FILL_5__3362_
timestamp 1701859473
transform 1 0 8030 0 -1 10670
box -12 -8 32 272
use FILL  FILL_5__3363_
timestamp 1701859473
transform 1 0 8150 0 1 10670
box -12 -8 32 272
use FILL  FILL_5__3364_
timestamp 1701859473
transform 1 0 7990 0 -1 11190
box -12 -8 32 272
use FILL  FILL_5__3365_
timestamp 1701859473
transform -1 0 7530 0 -1 11190
box -12 -8 32 272
use FILL  FILL_5__3366_
timestamp 1701859473
transform 1 0 7050 0 -1 11190
box -12 -8 32 272
use FILL  FILL_5__3367_
timestamp 1701859473
transform 1 0 6930 0 1 10670
box -12 -8 32 272
use FILL  FILL_5__3368_
timestamp 1701859473
transform 1 0 7270 0 -1 11190
box -12 -8 32 272
use FILL  FILL_5__3369_
timestamp 1701859473
transform 1 0 7750 0 -1 11190
box -12 -8 32 272
use FILL  FILL_5__3370_
timestamp 1701859473
transform 1 0 8270 0 -1 10670
box -12 -8 32 272
use FILL  FILL_5__3371_
timestamp 1701859473
transform 1 0 8370 0 1 10670
box -12 -8 32 272
use FILL  FILL_5__3372_
timestamp 1701859473
transform 1 0 9550 0 1 10670
box -12 -8 32 272
use FILL  FILL_5__3373_
timestamp 1701859473
transform -1 0 6650 0 -1 11190
box -12 -8 32 272
use FILL  FILL_5__3374_
timestamp 1701859473
transform 1 0 5750 0 1 10670
box -12 -8 32 272
use FILL  FILL_5__3375_
timestamp 1701859473
transform -1 0 6010 0 1 10670
box -12 -8 32 272
use FILL  FILL_5__3376_
timestamp 1701859473
transform -1 0 6230 0 1 10670
box -12 -8 32 272
use FILL  FILL_5__3377_
timestamp 1701859473
transform 1 0 6470 0 1 10670
box -12 -8 32 272
use FILL  FILL_5__3378_
timestamp 1701859473
transform 1 0 6410 0 -1 11190
box -12 -8 32 272
use FILL  FILL_5__3379_
timestamp 1701859473
transform 1 0 8730 0 -1 10670
box -12 -8 32 272
use FILL  FILL_5__3380_
timestamp 1701859473
transform 1 0 8850 0 1 10670
box -12 -8 32 272
use FILL  FILL_5__3381_
timestamp 1701859473
transform -1 0 6730 0 1 10670
box -12 -8 32 272
use FILL  FILL_5__3382_
timestamp 1701859473
transform 1 0 6190 0 -1 10670
box -12 -8 32 272
use FILL  FILL_5__3383_
timestamp 1701859473
transform -1 0 6450 0 -1 10670
box -12 -8 32 272
use FILL  FILL_5__3384_
timestamp 1701859473
transform -1 0 6890 0 -1 10670
box -12 -8 32 272
use FILL  FILL_5__3385_
timestamp 1701859473
transform 1 0 6650 0 -1 10670
box -12 -8 32 272
use FILL  FILL_5__3386_
timestamp 1701859473
transform 1 0 7130 0 -1 10670
box -12 -8 32 272
use FILL  FILL_5__3387_
timestamp 1701859473
transform 1 0 8490 0 -1 10670
box -12 -8 32 272
use FILL  FILL_5__3388_
timestamp 1701859473
transform 1 0 8610 0 1 10670
box -12 -8 32 272
use FILL  FILL_5__3389_
timestamp 1701859473
transform 1 0 10270 0 -1 10670
box -12 -8 32 272
use FILL  FILL_5__3390_
timestamp 1701859473
transform 1 0 9830 0 -1 10670
box -12 -8 32 272
use FILL  FILL_5__3391_
timestamp 1701859473
transform 1 0 10030 0 -1 10670
box -12 -8 32 272
use FILL  FILL_5__3392_
timestamp 1701859473
transform 1 0 10490 0 -1 10670
box -12 -8 32 272
use FILL  FILL_5__3393_
timestamp 1701859473
transform -1 0 11230 0 -1 10150
box -12 -8 32 272
use FILL  FILL_5__3394_
timestamp 1701859473
transform 1 0 7410 0 1 10150
box -12 -8 32 272
use FILL  FILL_5__3395_
timestamp 1701859473
transform 1 0 6470 0 1 10150
box -12 -8 32 272
use FILL  FILL_5__3396_
timestamp 1701859473
transform -1 0 6730 0 1 10150
box -12 -8 32 272
use FILL  FILL_5__3397_
timestamp 1701859473
transform -1 0 7050 0 -1 10150
box -12 -8 32 272
use FILL  FILL_5__3398_
timestamp 1701859473
transform 1 0 6330 0 -1 10150
box -12 -8 32 272
use FILL  FILL_5__3399_
timestamp 1701859473
transform -1 0 6810 0 -1 10150
box -12 -8 32 272
use FILL  FILL_5__3400_
timestamp 1701859473
transform -1 0 6990 0 1 10150
box -12 -8 32 272
use FILL  FILL_5__3401_
timestamp 1701859473
transform 1 0 7170 0 1 10150
box -12 -8 32 272
use FILL  FILL_5__3402_
timestamp 1701859473
transform -1 0 9110 0 1 10150
box -12 -8 32 272
use FILL  FILL_5__3403_
timestamp 1701859473
transform 1 0 9550 0 1 10150
box -12 -8 32 272
use FILL  FILL_5__3404_
timestamp 1701859473
transform -1 0 5810 0 1 9630
box -12 -8 32 272
use FILL  FILL_5__3405_
timestamp 1701859473
transform -1 0 6090 0 -1 10150
box -12 -8 32 272
use FILL  FILL_5__3406_
timestamp 1701859473
transform 1 0 6450 0 -1 9630
box -12 -8 32 272
use FILL  FILL_5__3407_
timestamp 1701859473
transform -1 0 6670 0 -1 9630
box -12 -8 32 272
use FILL  FILL_5__3408_
timestamp 1701859473
transform 1 0 6930 0 1 9630
box -12 -8 32 272
use FILL  FILL_5__3409_
timestamp 1701859473
transform -1 0 6550 0 -1 10150
box -12 -8 32 272
use FILL  FILL_5__3410_
timestamp 1701859473
transform 1 0 9290 0 -1 10150
box -12 -8 32 272
use FILL  FILL_5__3411_
timestamp 1701859473
transform 1 0 9310 0 1 10150
box -12 -8 32 272
use FILL  FILL_5__3412_
timestamp 1701859473
transform 1 0 10030 0 1 10150
box -12 -8 32 272
use FILL  FILL_5__3413_
timestamp 1701859473
transform -1 0 6050 0 1 9630
box -12 -8 32 272
use FILL  FILL_5__3414_
timestamp 1701859473
transform 1 0 8190 0 1 9110
box -12 -8 32 272
use FILL  FILL_5__3415_
timestamp 1701859473
transform 1 0 6470 0 1 9630
box -12 -8 32 272
use FILL  FILL_5__3416_
timestamp 1701859473
transform 1 0 7310 0 1 8590
box -12 -8 32 272
use FILL  FILL_5__3417_
timestamp 1701859473
transform 1 0 7390 0 -1 9110
box -12 -8 32 272
use FILL  FILL_5__3418_
timestamp 1701859473
transform -1 0 7530 0 -1 9630
box -12 -8 32 272
use FILL  FILL_5__3419_
timestamp 1701859473
transform 1 0 7290 0 -1 9630
box -12 -8 32 272
use FILL  FILL_5__3420_
timestamp 1701859473
transform -1 0 6870 0 -1 9630
box -12 -8 32 272
use FILL  FILL_5__3421_
timestamp 1701859473
transform -1 0 7090 0 -1 9630
box -12 -8 32 272
use FILL  FILL_5__3422_
timestamp 1701859473
transform -1 0 7190 0 1 9630
box -12 -8 32 272
use FILL  FILL_5__3423_
timestamp 1701859473
transform -1 0 8250 0 -1 9630
box -12 -8 32 272
use FILL  FILL_5__3424_
timestamp 1701859473
transform -1 0 7770 0 -1 9630
box -12 -8 32 272
use FILL  FILL_5__3425_
timestamp 1701859473
transform -1 0 7430 0 1 9630
box -12 -8 32 272
use FILL  FILL_5__3426_
timestamp 1701859473
transform -1 0 9070 0 -1 10150
box -12 -8 32 272
use FILL  FILL_5__3427_
timestamp 1701859473
transform 1 0 8830 0 -1 10150
box -12 -8 32 272
use FILL  FILL_5__3428_
timestamp 1701859473
transform 1 0 7510 0 1 8590
box -12 -8 32 272
use FILL  FILL_5__3429_
timestamp 1701859473
transform 1 0 7590 0 -1 9110
box -12 -8 32 272
use FILL  FILL_5__3430_
timestamp 1701859473
transform -1 0 7810 0 -1 9110
box -12 -8 32 272
use FILL  FILL_5__3431_
timestamp 1701859473
transform 1 0 7730 0 1 9110
box -12 -8 32 272
use FILL  FILL_5__3432_
timestamp 1701859473
transform 1 0 7970 0 1 9110
box -12 -8 32 272
use FILL  FILL_5__3433_
timestamp 1701859473
transform -1 0 8010 0 -1 9630
box -12 -8 32 272
use FILL  FILL_5__3434_
timestamp 1701859473
transform 1 0 7650 0 1 9630
box -12 -8 32 272
use FILL  FILL_5__3435_
timestamp 1701859473
transform 1 0 10270 0 1 10150
box -12 -8 32 272
use FILL  FILL_5__3436_
timestamp 1701859473
transform -1 0 10270 0 -1 10150
box -12 -8 32 272
use FILL  FILL_5__3437_
timestamp 1701859473
transform 1 0 10710 0 1 10150
box -12 -8 32 272
use FILL  FILL_5__3438_
timestamp 1701859473
transform 1 0 10490 0 1 10150
box -12 -8 32 272
use FILL  FILL_5__3439_
timestamp 1701859473
transform 1 0 10930 0 1 10150
box -12 -8 32 272
use FILL  FILL_5__3440_
timestamp 1701859473
transform -1 0 10750 0 -1 10150
box -12 -8 32 272
use FILL  FILL_5__3441_
timestamp 1701859473
transform -1 0 10610 0 1 9630
box -12 -8 32 272
use FILL  FILL_5__3442_
timestamp 1701859473
transform -1 0 10490 0 -1 10150
box -12 -8 32 272
use FILL  FILL_5__3443_
timestamp 1701859473
transform -1 0 11050 0 1 9630
box -12 -8 32 272
use FILL  FILL_5__3444_
timestamp 1701859473
transform -1 0 8450 0 -1 9630
box -12 -8 32 272
use FILL  FILL_5__3445_
timestamp 1701859473
transform -1 0 8150 0 1 9630
box -12 -8 32 272
use FILL  FILL_5__3446_
timestamp 1701859473
transform 1 0 8590 0 1 9630
box -12 -8 32 272
use FILL  FILL_5__3447_
timestamp 1701859473
transform 1 0 8370 0 1 9630
box -12 -8 32 272
use FILL  FILL_5__3448_
timestamp 1701859473
transform -1 0 8810 0 1 9630
box -12 -8 32 272
use FILL  FILL_5__3449_
timestamp 1701859473
transform -1 0 9850 0 1 10150
box -12 -8 32 272
use FILL  FILL_5__3450_
timestamp 1701859473
transform -1 0 9810 0 -1 10150
box -12 -8 32 272
use FILL  FILL_5__3451_
timestamp 1701859473
transform 1 0 9530 0 -1 10150
box -12 -8 32 272
use FILL  FILL_5__3452_
timestamp 1701859473
transform -1 0 9270 0 1 9630
box -12 -8 32 272
use FILL  FILL_5__3453_
timestamp 1701859473
transform -1 0 10030 0 -1 10150
box -12 -8 32 272
use FILL  FILL_5__3454_
timestamp 1701859473
transform 1 0 9470 0 1 9630
box -12 -8 32 272
use FILL  FILL_5__3455_
timestamp 1701859473
transform 1 0 9690 0 1 9630
box -12 -8 32 272
use FILL  FILL_5__3456_
timestamp 1701859473
transform -1 0 10390 0 1 9630
box -12 -8 32 272
use FILL  FILL_5__3457_
timestamp 1701859473
transform -1 0 9930 0 1 9630
box -12 -8 32 272
use FILL  FILL_5__3458_
timestamp 1701859473
transform -1 0 10170 0 1 9630
box -12 -8 32 272
use FILL  FILL_5__3459_
timestamp 1701859473
transform -1 0 10310 0 -1 9630
box -12 -8 32 272
use FILL  FILL_5__3460_
timestamp 1701859473
transform 1 0 10970 0 -1 10150
box -12 -8 32 272
use FILL  FILL_5__3461_
timestamp 1701859473
transform -1 0 11210 0 -1 9630
box -12 -8 32 272
use FILL  FILL_5__3462_
timestamp 1701859473
transform -1 0 10750 0 -1 9630
box -12 -8 32 272
use FILL  FILL_5__3463_
timestamp 1701859473
transform 1 0 10430 0 -1 11190
box -12 -8 32 272
use FILL  FILL_5__3464_
timestamp 1701859473
transform 1 0 9770 0 -1 11190
box -12 -8 32 272
use FILL  FILL_5__3465_
timestamp 1701859473
transform 1 0 10010 0 -1 11190
box -12 -8 32 272
use FILL  FILL_5__3466_
timestamp 1701859473
transform 1 0 10190 0 -1 11190
box -12 -8 32 272
use FILL  FILL_5__3467_
timestamp 1701859473
transform -1 0 11170 0 1 10670
box -12 -8 32 272
use FILL  FILL_5__3468_
timestamp 1701859473
transform 1 0 10670 0 1 10670
box -12 -8 32 272
use FILL  FILL_5__3469_
timestamp 1701859473
transform 1 0 9390 0 -1 10670
box -12 -8 32 272
use FILL  FILL_5__3470_
timestamp 1701859473
transform 1 0 9630 0 -1 10670
box -12 -8 32 272
use FILL  FILL_5__3471_
timestamp 1701859473
transform 1 0 9770 0 1 10670
box -12 -8 32 272
use FILL  FILL_5__3472_
timestamp 1701859473
transform -1 0 10030 0 1 10670
box -12 -8 32 272
use FILL  FILL_5__3473_
timestamp 1701859473
transform 1 0 8650 0 -1 11190
box -12 -8 32 272
use FILL  FILL_5__3474_
timestamp 1701859473
transform 1 0 8210 0 -1 11190
box -12 -8 32 272
use FILL  FILL_5__3475_
timestamp 1701859473
transform 1 0 8450 0 -1 11190
box -12 -8 32 272
use FILL  FILL_5__3476_
timestamp 1701859473
transform -1 0 8890 0 -1 11190
box -12 -8 32 272
use FILL  FILL_5__3477_
timestamp 1701859473
transform 1 0 9110 0 -1 11190
box -12 -8 32 272
use FILL  FILL_5__3478_
timestamp 1701859473
transform 1 0 9090 0 1 10670
box -12 -8 32 272
use FILL  FILL_5__3479_
timestamp 1701859473
transform 1 0 8370 0 -1 10150
box -12 -8 32 272
use FILL  FILL_5__3480_
timestamp 1701859473
transform -1 0 8630 0 -1 10150
box -12 -8 32 272
use FILL  FILL_5__3481_
timestamp 1701859473
transform -1 0 8410 0 1 9110
box -12 -8 32 272
use FILL  FILL_5__3482_
timestamp 1701859473
transform -1 0 8630 0 1 9110
box -12 -8 32 272
use FILL  FILL_5__3483_
timestamp 1701859473
transform 1 0 8810 0 1 10150
box -12 -8 32 272
use FILL  FILL_5__3484_
timestamp 1701859473
transform -1 0 10110 0 -1 9630
box -12 -8 32 272
use FILL  FILL_5__3485_
timestamp 1701859473
transform 1 0 11130 0 1 10150
box -12 -8 32 272
use FILL  FILL_5__3486_
timestamp 1701859473
transform 1 0 10470 0 1 9110
box -12 -8 32 272
use FILL  FILL_5__3487_
timestamp 1701859473
transform 1 0 10510 0 -1 9630
box -12 -8 32 272
use FILL  FILL_5__3488_
timestamp 1701859473
transform -1 0 10810 0 1 9630
box -12 -8 32 272
use FILL  FILL_5__3489_
timestamp 1701859473
transform 1 0 10650 0 -1 11190
box -12 -8 32 272
use FILL  FILL_5__3490_
timestamp 1701859473
transform 1 0 11110 0 -1 11190
box -12 -8 32 272
use FILL  FILL_5__3491_
timestamp 1701859473
transform -1 0 10910 0 -1 11190
box -12 -8 32 272
use FILL  FILL_5__3492_
timestamp 1701859473
transform -1 0 10470 0 1 10670
box -12 -8 32 272
use FILL  FILL_5__3493_
timestamp 1701859473
transform -1 0 10250 0 1 10670
box -12 -8 32 272
use FILL  FILL_5__3494_
timestamp 1701859473
transform 1 0 9350 0 1 10670
box -12 -8 32 272
use FILL  FILL_5__3495_
timestamp 1701859473
transform -1 0 9550 0 -1 11190
box -12 -8 32 272
use FILL  FILL_5__3496_
timestamp 1701859473
transform 1 0 9310 0 -1 11190
box -12 -8 32 272
use FILL  FILL_5__3497_
timestamp 1701859473
transform -1 0 9410 0 -1 9630
box -12 -8 32 272
use FILL  FILL_5__3498_
timestamp 1701859473
transform -1 0 8910 0 1 9110
box -12 -8 32 272
use FILL  FILL_5__3499_
timestamp 1701859473
transform 1 0 8430 0 -1 9110
box -12 -8 32 272
use FILL  FILL_5__3500_
timestamp 1701859473
transform 1 0 9810 0 1 9110
box -12 -8 32 272
use FILL  FILL_5__3501_
timestamp 1701859473
transform -1 0 10050 0 1 9110
box -12 -8 32 272
use FILL  FILL_5__3502_
timestamp 1701859473
transform -1 0 8310 0 -1 8590
box -12 -8 32 272
use FILL  FILL_5__3503_
timestamp 1701859473
transform -1 0 8690 0 -1 9630
box -12 -8 32 272
use FILL  FILL_5__3504_
timestamp 1701859473
transform 1 0 8910 0 -1 9630
box -12 -8 32 272
use FILL  FILL_5__3505_
timestamp 1701859473
transform -1 0 9170 0 -1 9630
box -12 -8 32 272
use FILL  FILL_5__3506_
timestamp 1701859473
transform -1 0 8690 0 1 8590
box -12 -8 32 272
use FILL  FILL_5__3507_
timestamp 1701859473
transform 1 0 10770 0 -1 9110
box -12 -8 32 272
use FILL  FILL_5__3508_
timestamp 1701859473
transform 1 0 10530 0 -1 9110
box -12 -8 32 272
use FILL  FILL_5__3509_
timestamp 1701859473
transform 1 0 8470 0 1 8590
box -12 -8 32 272
use FILL  FILL_5__3510_
timestamp 1701859473
transform -1 0 8930 0 1 8590
box -12 -8 32 272
use FILL  FILL_5__3511_
timestamp 1701859473
transform 1 0 9990 0 -1 270
box -12 -8 32 272
use FILL  FILL_5__3512_
timestamp 1701859473
transform 1 0 10990 0 -1 9110
box -12 -8 32 272
use FILL  FILL_5__3513_
timestamp 1701859473
transform 1 0 10970 0 -1 9630
box -12 -8 32 272
use FILL  FILL_5__3514_
timestamp 1701859473
transform 1 0 10930 0 1 10670
box -12 -8 32 272
use FILL  FILL_5__3515_
timestamp 1701859473
transform -1 0 10730 0 -1 10670
box -12 -8 32 272
use FILL  FILL_5__3516_
timestamp 1701859473
transform 1 0 10950 0 -1 10670
box -12 -8 32 272
use FILL  FILL_5__3517_
timestamp 1701859473
transform 1 0 9630 0 -1 9630
box -12 -8 32 272
use FILL  FILL_5__3518_
timestamp 1701859473
transform 1 0 9850 0 -1 9630
box -12 -8 32 272
use FILL  FILL_5__3519_
timestamp 1701859473
transform 1 0 9130 0 1 9110
box -12 -8 32 272
use FILL  FILL_5__3520_
timestamp 1701859473
transform -1 0 9370 0 1 9110
box -12 -8 32 272
use FILL  FILL_5__3521_
timestamp 1701859473
transform 1 0 6610 0 1 8590
box -12 -8 32 272
use FILL  FILL_5__3522_
timestamp 1701859473
transform 1 0 8010 0 -1 9110
box -12 -8 32 272
use FILL  FILL_5__3523_
timestamp 1701859473
transform 1 0 6810 0 1 8590
box -12 -8 32 272
use FILL  FILL_5__3524_
timestamp 1701859473
transform 1 0 7530 0 1 9110
box -12 -8 32 272
use FILL  FILL_5__3525_
timestamp 1701859473
transform 1 0 7070 0 1 9110
box -12 -8 32 272
use FILL  FILL_5__3526_
timestamp 1701859473
transform -1 0 7310 0 1 9110
box -12 -8 32 272
use FILL  FILL_5__3539_
timestamp 1701859473
transform 1 0 11170 0 -1 7030
box -12 -8 32 272
use FILL  FILL_5__3540_
timestamp 1701859473
transform 1 0 4670 0 1 10670
box -12 -8 32 272
use FILL  FILL_5__3541_
timestamp 1701859473
transform -1 0 130 0 1 5990
box -12 -8 32 272
use FILL  FILL_5__3542_
timestamp 1701859473
transform -1 0 130 0 -1 8070
box -12 -8 32 272
use FILL  FILL_5__3543_
timestamp 1701859473
transform -1 0 130 0 1 8590
box -12 -8 32 272
use FILL  FILL_5__3544_
timestamp 1701859473
transform -1 0 130 0 1 9110
box -12 -8 32 272
use FILL  FILL_5__3545_
timestamp 1701859473
transform -1 0 1970 0 -1 11190
box -12 -8 32 272
use FILL  FILL_5__3546_
timestamp 1701859473
transform -1 0 590 0 1 9110
box -12 -8 32 272
use FILL  FILL_5__3547_
timestamp 1701859473
transform 1 0 4710 0 -1 11190
box -12 -8 32 272
use FILL  FILL_5__3548_
timestamp 1701859473
transform 1 0 5310 0 1 10670
box -12 -8 32 272
use FILL  FILL_5__3549_
timestamp 1701859473
transform -1 0 4310 0 -1 11190
box -12 -8 32 272
use FILL  FILL_5__3550_
timestamp 1701859473
transform -1 0 5150 0 -1 11190
box -12 -8 32 272
use FILL  FILL_5__3551_
timestamp 1701859473
transform 1 0 5550 0 -1 11190
box -12 -8 32 272
use FILL  FILL_5__3552_
timestamp 1701859473
transform 1 0 5330 0 -1 11190
box -12 -8 32 272
use FILL  FILL_5__3553_
timestamp 1701859473
transform -1 0 130 0 -1 5990
box -12 -8 32 272
use FILL  FILL_5__3554_
timestamp 1701859473
transform -1 0 330 0 1 7030
box -12 -8 32 272
use FILL  FILL_5__3555_
timestamp 1701859473
transform -1 0 5110 0 1 10670
box -12 -8 32 272
use FILL  FILL_5__3556_
timestamp 1701859473
transform 1 0 6250 0 1 10150
box -12 -8 32 272
use FILL  FILL_5__3557_
timestamp 1701859473
transform -1 0 5790 0 -1 11190
box -12 -8 32 272
use FILL  FILL_5__3558_
timestamp 1701859473
transform 1 0 6190 0 -1 11190
box -12 -8 32 272
use FILL  FILL_5__3559_
timestamp 1701859473
transform -1 0 4850 0 -1 10670
box -12 -8 32 272
use FILL  FILL_5__3560_
timestamp 1701859473
transform 1 0 5530 0 1 10670
box -12 -8 32 272
use FILL  FILL_5__3561_
timestamp 1701859473
transform 1 0 5970 0 -1 11190
box -12 -8 32 272
use FILL  FILL_5__3562_
timestamp 1701859473
transform 1 0 5770 0 1 10150
box -12 -8 32 272
use FILL  FILL_5__3563_
timestamp 1701859473
transform 1 0 5230 0 1 3390
box -12 -8 32 272
use FILL  FILL_5_BUFX2_insert0
timestamp 1701859473
transform 1 0 5850 0 -1 10150
box -12 -8 32 272
use FILL  FILL_5_BUFX2_insert1
timestamp 1701859473
transform 1 0 6610 0 1 2350
box -12 -8 32 272
use FILL  FILL_5_BUFX2_insert2
timestamp 1701859473
transform 1 0 5450 0 -1 1830
box -12 -8 32 272
use FILL  FILL_5_BUFX2_insert3
timestamp 1701859473
transform -1 0 590 0 -1 5470
box -12 -8 32 272
use FILL  FILL_5_BUFX2_insert4
timestamp 1701859473
transform 1 0 3330 0 1 4950
box -12 -8 32 272
use FILL  FILL_5_BUFX2_insert5
timestamp 1701859473
transform 1 0 1390 0 -1 1830
box -12 -8 32 272
use FILL  FILL_5_BUFX2_insert6
timestamp 1701859473
transform -1 0 130 0 -1 11190
box -12 -8 32 272
use FILL  FILL_5_BUFX2_insert7
timestamp 1701859473
transform 1 0 1690 0 1 10670
box -12 -8 32 272
use FILL  FILL_5_BUFX2_insert8
timestamp 1701859473
transform 1 0 1650 0 1 1830
box -12 -8 32 272
use FILL  FILL_5_BUFX2_insert9
timestamp 1701859473
transform 1 0 1950 0 -1 3910
box -12 -8 32 272
use FILL  FILL_5_BUFX2_insert10
timestamp 1701859473
transform 1 0 1770 0 -1 4430
box -12 -8 32 272
use FILL  FILL_5_BUFX2_insert11
timestamp 1701859473
transform -1 0 1750 0 -1 3910
box -12 -8 32 272
use FILL  FILL_5_BUFX2_insert12
timestamp 1701859473
transform -1 0 1530 0 -1 3910
box -12 -8 32 272
use FILL  FILL_5_BUFX2_insert13
timestamp 1701859473
transform -1 0 1430 0 -1 1310
box -12 -8 32 272
use FILL  FILL_5_BUFX2_insert14
timestamp 1701859473
transform -1 0 3670 0 1 3390
box -12 -8 32 272
use FILL  FILL_5_BUFX2_insert15
timestamp 1701859473
transform 1 0 4550 0 -1 5470
box -12 -8 32 272
use FILL  FILL_5_BUFX2_insert16
timestamp 1701859473
transform 1 0 1350 0 -1 4950
box -12 -8 32 272
use FILL  FILL_5_BUFX2_insert17
timestamp 1701859473
transform 1 0 3630 0 1 1310
box -12 -8 32 272
use FILL  FILL_5_BUFX2_insert18
timestamp 1701859473
transform -1 0 9770 0 1 2350
box -12 -8 32 272
use FILL  FILL_5_BUFX2_insert19
timestamp 1701859473
transform -1 0 8510 0 -1 790
box -12 -8 32 272
use FILL  FILL_5_BUFX2_insert20
timestamp 1701859473
transform 1 0 9970 0 1 2350
box -12 -8 32 272
use FILL  FILL_5_BUFX2_insert21
timestamp 1701859473
transform -1 0 7810 0 -1 1310
box -12 -8 32 272
use FILL  FILL_5_BUFX2_insert22
timestamp 1701859473
transform -1 0 3210 0 -1 2870
box -12 -8 32 272
use FILL  FILL_5_BUFX2_insert23
timestamp 1701859473
transform -1 0 2750 0 -1 4950
box -12 -8 32 272
use FILL  FILL_5_BUFX2_insert24
timestamp 1701859473
transform -1 0 3650 0 -1 4430
box -12 -8 32 272
use FILL  FILL_5_BUFX2_insert25
timestamp 1701859473
transform 1 0 4390 0 1 4430
box -12 -8 32 272
use FILL  FILL_5_BUFX2_insert26
timestamp 1701859473
transform 1 0 4210 0 1 2870
box -12 -8 32 272
use FILL  FILL_5_BUFX2_insert27
timestamp 1701859473
transform 1 0 9610 0 1 4950
box -12 -8 32 272
use FILL  FILL_5_BUFX2_insert28
timestamp 1701859473
transform -1 0 7490 0 -1 5990
box -12 -8 32 272
use FILL  FILL_5_BUFX2_insert29
timestamp 1701859473
transform -1 0 1290 0 1 6510
box -12 -8 32 272
use FILL  FILL_5_BUFX2_insert30
timestamp 1701859473
transform -1 0 8790 0 -1 3910
box -12 -8 32 272
use FILL  FILL_5_BUFX2_insert31
timestamp 1701859473
transform -1 0 9570 0 1 3910
box -12 -8 32 272
use FILL  FILL_5_BUFX2_insert32
timestamp 1701859473
transform 1 0 5870 0 -1 3910
box -12 -8 32 272
use FILL  FILL_5_BUFX2_insert33
timestamp 1701859473
transform -1 0 9550 0 -1 4950
box -12 -8 32 272
use FILL  FILL_5_BUFX2_insert34
timestamp 1701859473
transform 1 0 5210 0 1 8590
box -12 -8 32 272
use FILL  FILL_5_BUFX2_insert35
timestamp 1701859473
transform -1 0 5970 0 1 7550
box -12 -8 32 272
use FILL  FILL_5_BUFX2_insert36
timestamp 1701859473
transform -1 0 1210 0 1 8590
box -12 -8 32 272
use FILL  FILL_5_BUFX2_insert37
timestamp 1701859473
transform -1 0 9590 0 1 8590
box -12 -8 32 272
use FILL  FILL_5_BUFX2_insert49
timestamp 1701859473
transform -1 0 3050 0 1 6510
box -12 -8 32 272
use FILL  FILL_5_BUFX2_insert50
timestamp 1701859473
transform 1 0 2350 0 -1 8590
box -12 -8 32 272
use FILL  FILL_5_BUFX2_insert51
timestamp 1701859473
transform 1 0 3210 0 -1 8590
box -12 -8 32 272
use FILL  FILL_5_BUFX2_insert52
timestamp 1701859473
transform 1 0 3390 0 1 5470
box -12 -8 32 272
use FILL  FILL_5_BUFX2_insert53
timestamp 1701859473
transform -1 0 11230 0 1 9110
box -12 -8 32 272
use FILL  FILL_5_BUFX2_insert54
timestamp 1701859473
transform -1 0 9170 0 1 8590
box -12 -8 32 272
use FILL  FILL_5_BUFX2_insert55
timestamp 1701859473
transform -1 0 9610 0 1 9110
box -12 -8 32 272
use FILL  FILL_5_BUFX2_insert56
timestamp 1701859473
transform -1 0 10270 0 1 9110
box -12 -8 32 272
use FILL  FILL_5_BUFX2_insert57
timestamp 1701859473
transform -1 0 11230 0 -1 2350
box -12 -8 32 272
use FILL  FILL_5_BUFX2_insert58
timestamp 1701859473
transform -1 0 8970 0 1 2870
box -12 -8 32 272
use FILL  FILL_5_BUFX2_insert59
timestamp 1701859473
transform -1 0 7550 0 1 1830
box -12 -8 32 272
use FILL  FILL_5_BUFX2_insert60
timestamp 1701859473
transform 1 0 10890 0 1 1830
box -12 -8 32 272
use FILL  FILL_5_BUFX2_insert61
timestamp 1701859473
transform -1 0 11170 0 1 2870
box -12 -8 32 272
use FILL  FILL_5_BUFX2_insert62
timestamp 1701859473
transform 1 0 2210 0 1 3910
box -12 -8 32 272
use FILL  FILL_5_BUFX2_insert63
timestamp 1701859473
transform 1 0 2130 0 1 3390
box -12 -8 32 272
use FILL  FILL_5_BUFX2_insert64
timestamp 1701859473
transform -1 0 1790 0 1 3910
box -12 -8 32 272
use FILL  FILL_5_BUFX2_insert65
timestamp 1701859473
transform -1 0 1730 0 1 3390
box -12 -8 32 272
use FILL  FILL_5_BUFX2_insert66
timestamp 1701859473
transform -1 0 4310 0 1 1310
box -12 -8 32 272
use FILL  FILL_5_BUFX2_insert67
timestamp 1701859473
transform -1 0 3610 0 -1 10150
box -12 -8 32 272
use FILL  FILL_5_BUFX2_insert68
timestamp 1701859473
transform -1 0 7170 0 1 2870
box -12 -8 32 272
use FILL  FILL_5_BUFX2_insert69
timestamp 1701859473
transform -1 0 5650 0 -1 3390
box -12 -8 32 272
use FILL  FILL_5_BUFX2_insert70
timestamp 1701859473
transform -1 0 3670 0 -1 1830
box -12 -8 32 272
use FILL  FILL_5_BUFX2_insert71
timestamp 1701859473
transform -1 0 7310 0 1 2350
box -12 -8 32 272
use FILL  FILL_5_BUFX2_insert72
timestamp 1701859473
transform -1 0 6490 0 1 1310
box -12 -8 32 272
use FILL  FILL_5_BUFX2_insert73
timestamp 1701859473
transform 1 0 3610 0 1 5470
box -12 -8 32 272
use FILL  FILL_5_BUFX2_insert74
timestamp 1701859473
transform 1 0 7570 0 -1 2350
box -12 -8 32 272
use FILL  FILL_5_BUFX2_insert75
timestamp 1701859473
transform 1 0 7590 0 1 2870
box -12 -8 32 272
use FILL  FILL_5_BUFX2_insert76
timestamp 1701859473
transform 1 0 7370 0 1 2870
box -12 -8 32 272
use FILL  FILL_5_BUFX2_insert77
timestamp 1701859473
transform -1 0 3430 0 -1 2870
box -12 -8 32 272
use FILL  FILL_5_BUFX2_insert78
timestamp 1701859473
transform 1 0 1930 0 -1 2870
box -12 -8 32 272
use FILL  FILL_5_BUFX2_insert79
timestamp 1701859473
transform -1 0 2170 0 -1 2870
box -12 -8 32 272
use FILL  FILL_5_BUFX2_insert80
timestamp 1701859473
transform 1 0 2410 0 1 4430
box -12 -8 32 272
use FILL  FILL_5_BUFX2_insert81
timestamp 1701859473
transform -1 0 2010 0 1 3910
box -12 -8 32 272
use FILL  FILL_5_BUFX2_insert82
timestamp 1701859473
transform -1 0 330 0 1 8590
box -12 -8 32 272
use FILL  FILL_5_BUFX2_insert83
timestamp 1701859473
transform 1 0 4210 0 -1 10150
box -12 -8 32 272
use FILL  FILL_5_BUFX2_insert84
timestamp 1701859473
transform 1 0 4170 0 -1 7550
box -12 -8 32 272
use FILL  FILL_5_BUFX2_insert85
timestamp 1701859473
transform -1 0 130 0 -1 6510
box -12 -8 32 272
use FILL  FILL_5_BUFX2_insert86
timestamp 1701859473
transform 1 0 1930 0 -1 10150
box -12 -8 32 272
use FILL  FILL_5_CLKBUF1_insert38
timestamp 1701859473
transform 1 0 2930 0 -1 7550
box -12 -8 32 272
use FILL  FILL_5_CLKBUF1_insert39
timestamp 1701859473
transform -1 0 4730 0 -1 6510
box -12 -8 32 272
use FILL  FILL_5_CLKBUF1_insert40
timestamp 1701859473
transform -1 0 1030 0 -1 4950
box -12 -8 32 272
use FILL  FILL_5_CLKBUF1_insert41
timestamp 1701859473
transform -1 0 10690 0 -1 270
box -12 -8 32 272
use FILL  FILL_5_CLKBUF1_insert42
timestamp 1701859473
transform 1 0 9750 0 -1 4950
box -12 -8 32 272
use FILL  FILL_5_CLKBUF1_insert43
timestamp 1701859473
transform -1 0 11070 0 1 7030
box -12 -8 32 272
use FILL  FILL_5_CLKBUF1_insert44
timestamp 1701859473
transform -1 0 10810 0 1 4430
box -12 -8 32 272
use FILL  FILL_5_CLKBUF1_insert45
timestamp 1701859473
transform 1 0 5730 0 -1 6510
box -12 -8 32 272
use FILL  FILL_5_CLKBUF1_insert46
timestamp 1701859473
transform 1 0 4050 0 1 5990
box -12 -8 32 272
use FILL  FILL_5_CLKBUF1_insert47
timestamp 1701859473
transform -1 0 2170 0 1 7550
box -12 -8 32 272
use FILL  FILL_5_CLKBUF1_insert48
timestamp 1701859473
transform -1 0 10850 0 -1 7030
box -12 -8 32 272
use FILL  FILL_6__1668_
timestamp 1701859473
transform 1 0 6810 0 -1 3390
box -12 -8 32 272
use FILL  FILL_6__1669_
timestamp 1701859473
transform -1 0 6850 0 -1 790
box -12 -8 32 272
use FILL  FILL_6__1670_
timestamp 1701859473
transform 1 0 6630 0 -1 2870
box -12 -8 32 272
use FILL  FILL_6__1671_
timestamp 1701859473
transform -1 0 6430 0 -1 8590
box -12 -8 32 272
use FILL  FILL_6__1672_
timestamp 1701859473
transform 1 0 5990 0 -1 10670
box -12 -8 32 272
use FILL  FILL_6__1673_
timestamp 1701859473
transform 1 0 6390 0 1 8590
box -12 -8 32 272
use FILL  FILL_6__1674_
timestamp 1701859473
transform -1 0 6470 0 -1 9110
box -12 -8 32 272
use FILL  FILL_6__1675_
timestamp 1701859473
transform 1 0 130 0 -1 5470
box -12 -8 32 272
use FILL  FILL_6__1676_
timestamp 1701859473
transform -1 0 370 0 -1 5470
box -12 -8 32 272
use FILL  FILL_6__1677_
timestamp 1701859473
transform -1 0 610 0 1 5470
box -12 -8 32 272
use FILL  FILL_6__1678_
timestamp 1701859473
transform 1 0 130 0 -1 10670
box -12 -8 32 272
use FILL  FILL_6__1679_
timestamp 1701859473
transform -1 0 350 0 -1 11190
box -12 -8 32 272
use FILL  FILL_6__1680_
timestamp 1701859473
transform 1 0 330 0 -1 10670
box -12 -8 32 272
use FILL  FILL_6__1681_
timestamp 1701859473
transform -1 0 150 0 -1 7030
box -12 -8 32 272
use FILL  FILL_6__1682_
timestamp 1701859473
transform -1 0 150 0 1 7030
box -12 -8 32 272
use FILL  FILL_6__1683_
timestamp 1701859473
transform 1 0 130 0 1 6510
box -12 -8 32 272
use FILL  FILL_6__1684_
timestamp 1701859473
transform 1 0 1010 0 -1 11190
box -12 -8 32 272
use FILL  FILL_6__1685_
timestamp 1701859473
transform -1 0 1270 0 -1 11190
box -12 -8 32 272
use FILL  FILL_6__1686_
timestamp 1701859473
transform -1 0 1070 0 1 10670
box -12 -8 32 272
use FILL  FILL_6__1687_
timestamp 1701859473
transform 1 0 1490 0 -1 11190
box -12 -8 32 272
use FILL  FILL_6__1688_
timestamp 1701859473
transform -1 0 1750 0 -1 11190
box -12 -8 32 272
use FILL  FILL_6__1689_
timestamp 1701859473
transform -1 0 2010 0 1 10150
box -12 -8 32 272
use FILL  FILL_6__1690_
timestamp 1701859473
transform 1 0 2170 0 1 9110
box -12 -8 32 272
use FILL  FILL_6__1691_
timestamp 1701859473
transform -1 0 2190 0 -1 9110
box -12 -8 32 272
use FILL  FILL_6__1692_
timestamp 1701859473
transform 1 0 130 0 1 790
box -12 -8 32 272
use FILL  FILL_6__1693_
timestamp 1701859473
transform 1 0 130 0 -1 1310
box -12 -8 32 272
use FILL  FILL_6__1694_
timestamp 1701859473
transform 1 0 550 0 -1 270
box -12 -8 32 272
use FILL  FILL_6__1695_
timestamp 1701859473
transform -1 0 770 0 -1 270
box -12 -8 32 272
use FILL  FILL_6__1696_
timestamp 1701859473
transform 1 0 1190 0 1 2870
box -12 -8 32 272
use FILL  FILL_6__1697_
timestamp 1701859473
transform -1 0 2850 0 -1 2870
box -12 -8 32 272
use FILL  FILL_6__1698_
timestamp 1701859473
transform -1 0 1950 0 1 3390
box -12 -8 32 272
use FILL  FILL_6__1699_
timestamp 1701859473
transform 1 0 3870 0 1 3390
box -12 -8 32 272
use FILL  FILL_6__1700_
timestamp 1701859473
transform -1 0 2670 0 -1 3910
box -12 -8 32 272
use FILL  FILL_6__1701_
timestamp 1701859473
transform -1 0 1210 0 1 270
box -12 -8 32 272
use FILL  FILL_6__1702_
timestamp 1701859473
transform 1 0 970 0 1 270
box -12 -8 32 272
use FILL  FILL_6__1703_
timestamp 1701859473
transform -1 0 1450 0 1 1830
box -12 -8 32 272
use FILL  FILL_6__1704_
timestamp 1701859473
transform -1 0 9210 0 1 2870
box -12 -8 32 272
use FILL  FILL_6__1705_
timestamp 1701859473
transform 1 0 9830 0 -1 790
box -12 -8 32 272
use FILL  FILL_6__1706_
timestamp 1701859473
transform -1 0 8050 0 -1 4950
box -12 -8 32 272
use FILL  FILL_6__1707_
timestamp 1701859473
transform 1 0 8490 0 -1 4950
box -12 -8 32 272
use FILL  FILL_6__1708_
timestamp 1701859473
transform 1 0 5110 0 -1 5990
box -12 -8 32 272
use FILL  FILL_6__1709_
timestamp 1701859473
transform -1 0 11210 0 1 5990
box -12 -8 32 272
use FILL  FILL_6__1710_
timestamp 1701859473
transform 1 0 5490 0 -1 5470
box -12 -8 32 272
use FILL  FILL_6__1711_
timestamp 1701859473
transform -1 0 5330 0 -1 5990
box -12 -8 32 272
use FILL  FILL_6__1712_
timestamp 1701859473
transform -1 0 5150 0 1 5470
box -12 -8 32 272
use FILL  FILL_6__1713_
timestamp 1701859473
transform 1 0 8010 0 1 4430
box -12 -8 32 272
use FILL  FILL_6__1714_
timestamp 1701859473
transform 1 0 7810 0 1 4950
box -12 -8 32 272
use FILL  FILL_6__1715_
timestamp 1701859473
transform -1 0 8050 0 1 4950
box -12 -8 32 272
use FILL  FILL_6__1716_
timestamp 1701859473
transform -1 0 8270 0 1 4430
box -12 -8 32 272
use FILL  FILL_6__1717_
timestamp 1701859473
transform -1 0 8050 0 1 1310
box -12 -8 32 272
use FILL  FILL_6__1718_
timestamp 1701859473
transform -1 0 5990 0 1 5990
box -12 -8 32 272
use FILL  FILL_6__1719_
timestamp 1701859473
transform -1 0 6850 0 -1 5990
box -12 -8 32 272
use FILL  FILL_6__1720_
timestamp 1701859473
transform -1 0 6830 0 1 5470
box -12 -8 32 272
use FILL  FILL_6__1721_
timestamp 1701859473
transform -1 0 7070 0 1 5470
box -12 -8 32 272
use FILL  FILL_6__1722_
timestamp 1701859473
transform -1 0 7770 0 1 4430
box -12 -8 32 272
use FILL  FILL_6__1723_
timestamp 1701859473
transform 1 0 7990 0 1 1830
box -12 -8 32 272
use FILL  FILL_6__1724_
timestamp 1701859473
transform -1 0 8030 0 -1 1310
box -12 -8 32 272
use FILL  FILL_6__1725_
timestamp 1701859473
transform 1 0 6630 0 1 5990
box -12 -8 32 272
use FILL  FILL_6__1726_
timestamp 1701859473
transform 1 0 6830 0 1 5990
box -12 -8 32 272
use FILL  FILL_6__1727_
timestamp 1701859473
transform -1 0 7070 0 1 5990
box -12 -8 32 272
use FILL  FILL_6__1728_
timestamp 1701859473
transform 1 0 7770 0 1 5990
box -12 -8 32 272
use FILL  FILL_6__1729_
timestamp 1701859473
transform -1 0 7710 0 -1 5990
box -12 -8 32 272
use FILL  FILL_6__1730_
timestamp 1701859473
transform -1 0 8190 0 1 3390
box -12 -8 32 272
use FILL  FILL_6__1731_
timestamp 1701859473
transform -1 0 8050 0 -1 270
box -12 -8 32 272
use FILL  FILL_6__1732_
timestamp 1701859473
transform -1 0 8010 0 1 5470
box -12 -8 32 272
use FILL  FILL_6__1733_
timestamp 1701859473
transform -1 0 8230 0 1 5470
box -12 -8 32 272
use FILL  FILL_6__1734_
timestamp 1701859473
transform 1 0 8190 0 -1 5470
box -12 -8 32 272
use FILL  FILL_6__1735_
timestamp 1701859473
transform 1 0 8650 0 -1 5470
box -12 -8 32 272
use FILL  FILL_6__1736_
timestamp 1701859473
transform 1 0 8490 0 1 4950
box -12 -8 32 272
use FILL  FILL_6__1737_
timestamp 1701859473
transform -1 0 8570 0 -1 3910
box -12 -8 32 272
use FILL  FILL_6__1738_
timestamp 1701859473
transform 1 0 8970 0 1 790
box -12 -8 32 272
use FILL  FILL_6__1739_
timestamp 1701859473
transform -1 0 9190 0 -1 790
box -12 -8 32 272
use FILL  FILL_6__1740_
timestamp 1701859473
transform 1 0 6550 0 1 270
box -12 -8 32 272
use FILL  FILL_6__1741_
timestamp 1701859473
transform 1 0 6450 0 1 790
box -12 -8 32 272
use FILL  FILL_6__1742_
timestamp 1701859473
transform -1 0 6390 0 -1 790
box -12 -8 32 272
use FILL  FILL_6__1743_
timestamp 1701859473
transform -1 0 2390 0 -1 3390
box -12 -8 32 272
use FILL  FILL_6__1744_
timestamp 1701859473
transform 1 0 370 0 -1 4950
box -12 -8 32 272
use FILL  FILL_6__1745_
timestamp 1701859473
transform 1 0 2190 0 -1 3910
box -12 -8 32 272
use FILL  FILL_6__1746_
timestamp 1701859473
transform -1 0 5210 0 -1 3390
box -12 -8 32 272
use FILL  FILL_6__1747_
timestamp 1701859473
transform -1 0 370 0 -1 270
box -12 -8 32 272
use FILL  FILL_6__1748_
timestamp 1701859473
transform -1 0 570 0 1 270
box -12 -8 32 272
use FILL  FILL_6__1749_
timestamp 1701859473
transform -1 0 1010 0 1 1310
box -12 -8 32 272
use FILL  FILL_6__1750_
timestamp 1701859473
transform -1 0 1230 0 1 1310
box -12 -8 32 272
use FILL  FILL_6__1751_
timestamp 1701859473
transform -1 0 4590 0 -1 2870
box -12 -8 32 272
use FILL  FILL_6__1752_
timestamp 1701859473
transform 1 0 4790 0 -1 2870
box -12 -8 32 272
use FILL  FILL_6__1753_
timestamp 1701859473
transform -1 0 4410 0 1 790
box -12 -8 32 272
use FILL  FILL_6__1754_
timestamp 1701859473
transform 1 0 350 0 -1 790
box -12 -8 32 272
use FILL  FILL_6__1755_
timestamp 1701859473
transform -1 0 570 0 -1 790
box -12 -8 32 272
use FILL  FILL_6__1756_
timestamp 1701859473
transform -1 0 150 0 -1 270
box -12 -8 32 272
use FILL  FILL_6__1757_
timestamp 1701859473
transform 1 0 750 0 -1 790
box -12 -8 32 272
use FILL  FILL_6__1758_
timestamp 1701859473
transform 1 0 130 0 1 2350
box -12 -8 32 272
use FILL  FILL_6__1759_
timestamp 1701859473
transform -1 0 2630 0 -1 2870
box -12 -8 32 272
use FILL  FILL_6__1760_
timestamp 1701859473
transform 1 0 3010 0 -1 2870
box -12 -8 32 272
use FILL  FILL_6__1761_
timestamp 1701859473
transform -1 0 3330 0 -1 3390
box -12 -8 32 272
use FILL  FILL_6__1762_
timestamp 1701859473
transform -1 0 150 0 1 270
box -12 -8 32 272
use FILL  FILL_6__1763_
timestamp 1701859473
transform 1 0 130 0 -1 790
box -12 -8 32 272
use FILL  FILL_6__1764_
timestamp 1701859473
transform 1 0 570 0 1 1310
box -12 -8 32 272
use FILL  FILL_6__1765_
timestamp 1701859473
transform 1 0 1430 0 1 1310
box -12 -8 32 272
use FILL  FILL_6__1766_
timestamp 1701859473
transform -1 0 3230 0 -1 1830
box -12 -8 32 272
use FILL  FILL_6__1767_
timestamp 1701859473
transform 1 0 1530 0 -1 4430
box -12 -8 32 272
use FILL  FILL_6__1768_
timestamp 1701859473
transform 1 0 350 0 -1 1310
box -12 -8 32 272
use FILL  FILL_6__1769_
timestamp 1701859473
transform -1 0 570 0 1 1830
box -12 -8 32 272
use FILL  FILL_6__1770_
timestamp 1701859473
transform 1 0 2170 0 -1 3390
box -12 -8 32 272
use FILL  FILL_6__1771_
timestamp 1701859473
transform -1 0 2430 0 -1 3910
box -12 -8 32 272
use FILL  FILL_6__1772_
timestamp 1701859473
transform -1 0 3090 0 -1 3910
box -12 -8 32 272
use FILL  FILL_6__1773_
timestamp 1701859473
transform 1 0 3990 0 1 2870
box -12 -8 32 272
use FILL  FILL_6__1774_
timestamp 1701859473
transform -1 0 5370 0 -1 2350
box -12 -8 32 272
use FILL  FILL_6__1775_
timestamp 1701859473
transform 1 0 330 0 1 790
box -12 -8 32 272
use FILL  FILL_6__1776_
timestamp 1701859473
transform -1 0 370 0 1 1310
box -12 -8 32 272
use FILL  FILL_6__1777_
timestamp 1701859473
transform 1 0 790 0 -1 1830
box -12 -8 32 272
use FILL  FILL_6__1778_
timestamp 1701859473
transform -1 0 4510 0 1 5470
box -12 -8 32 272
use FILL  FILL_6__1779_
timestamp 1701859473
transform -1 0 6150 0 -1 5470
box -12 -8 32 272
use FILL  FILL_6__1780_
timestamp 1701859473
transform 1 0 4870 0 1 2870
box -12 -8 32 272
use FILL  FILL_6__1781_
timestamp 1701859473
transform 1 0 4450 0 1 2870
box -12 -8 32 272
use FILL  FILL_6__1782_
timestamp 1701859473
transform -1 0 150 0 1 1310
box -12 -8 32 272
use FILL  FILL_6__1783_
timestamp 1701859473
transform -1 0 1430 0 1 2870
box -12 -8 32 272
use FILL  FILL_6__1784_
timestamp 1701859473
transform -1 0 5130 0 1 2870
box -12 -8 32 272
use FILL  FILL_6__1785_
timestamp 1701859473
transform 1 0 5050 0 -1 2870
box -12 -8 32 272
use FILL  FILL_6__1786_
timestamp 1701859473
transform -1 0 5130 0 -1 2350
box -12 -8 32 272
use FILL  FILL_6__1787_
timestamp 1701859473
transform 1 0 5110 0 1 2350
box -12 -8 32 272
use FILL  FILL_6__1788_
timestamp 1701859473
transform -1 0 4910 0 -1 2350
box -12 -8 32 272
use FILL  FILL_6__1789_
timestamp 1701859473
transform 1 0 130 0 1 1830
box -12 -8 32 272
use FILL  FILL_6__1790_
timestamp 1701859473
transform -1 0 370 0 -1 2350
box -12 -8 32 272
use FILL  FILL_6__1791_
timestamp 1701859473
transform -1 0 2170 0 -1 2350
box -12 -8 32 272
use FILL  FILL_6__1792_
timestamp 1701859473
transform -1 0 3550 0 -1 2350
box -12 -8 32 272
use FILL  FILL_6__1793_
timestamp 1701859473
transform -1 0 4650 0 1 1830
box -12 -8 32 272
use FILL  FILL_6__1794_
timestamp 1701859473
transform 1 0 970 0 1 1830
box -12 -8 32 272
use FILL  FILL_6__1795_
timestamp 1701859473
transform -1 0 2230 0 1 2350
box -12 -8 32 272
use FILL  FILL_6__1796_
timestamp 1701859473
transform -1 0 1850 0 -1 1830
box -12 -8 32 272
use FILL  FILL_6__1797_
timestamp 1701859473
transform 1 0 2070 0 -1 1830
box -12 -8 32 272
use FILL  FILL_6__1798_
timestamp 1701859473
transform 1 0 990 0 -1 1310
box -12 -8 32 272
use FILL  FILL_6__1799_
timestamp 1701859473
transform 1 0 3810 0 1 3910
box -12 -8 32 272
use FILL  FILL_6__1800_
timestamp 1701859473
transform 1 0 3490 0 1 1830
box -12 -8 32 272
use FILL  FILL_6__1801_
timestamp 1701859473
transform -1 0 1230 0 1 1830
box -12 -8 32 272
use FILL  FILL_6__1802_
timestamp 1701859473
transform -1 0 3770 0 1 2350
box -12 -8 32 272
use FILL  FILL_6__1803_
timestamp 1701859473
transform -1 0 3990 0 1 2350
box -12 -8 32 272
use FILL  FILL_6__1804_
timestamp 1701859473
transform -1 0 4230 0 1 2350
box -12 -8 32 272
use FILL  FILL_6__1805_
timestamp 1701859473
transform 1 0 5530 0 1 2350
box -12 -8 32 272
use FILL  FILL_6__1806_
timestamp 1701859473
transform -1 0 4930 0 1 2350
box -12 -8 32 272
use FILL  FILL_6__1807_
timestamp 1701859473
transform -1 0 5330 0 1 2350
box -12 -8 32 272
use FILL  FILL_6__1808_
timestamp 1701859473
transform 1 0 4850 0 1 1830
box -12 -8 32 272
use FILL  FILL_6__1809_
timestamp 1701859473
transform -1 0 7210 0 -1 270
box -12 -8 32 272
use FILL  FILL_6__1810_
timestamp 1701859473
transform -1 0 7190 0 1 1310
box -12 -8 32 272
use FILL  FILL_6__1811_
timestamp 1701859473
transform 1 0 7530 0 -1 1830
box -12 -8 32 272
use FILL  FILL_6__1812_
timestamp 1701859473
transform -1 0 7610 0 -1 1310
box -12 -8 32 272
use FILL  FILL_6__1813_
timestamp 1701859473
transform 1 0 9190 0 1 790
box -12 -8 32 272
use FILL  FILL_6__1814_
timestamp 1701859473
transform -1 0 8230 0 -1 1830
box -12 -8 32 272
use FILL  FILL_6__1815_
timestamp 1701859473
transform 1 0 8430 0 1 2350
box -12 -8 32 272
use FILL  FILL_6__1816_
timestamp 1701859473
transform -1 0 9710 0 -1 2350
box -12 -8 32 272
use FILL  FILL_6__1817_
timestamp 1701859473
transform -1 0 9430 0 1 1310
box -12 -8 32 272
use FILL  FILL_6__1818_
timestamp 1701859473
transform -1 0 9630 0 1 270
box -12 -8 32 272
use FILL  FILL_6__1819_
timestamp 1701859473
transform -1 0 8450 0 -1 1830
box -12 -8 32 272
use FILL  FILL_6__1820_
timestamp 1701859473
transform -1 0 8530 0 1 1310
box -12 -8 32 272
use FILL  FILL_6__1821_
timestamp 1701859473
transform -1 0 4970 0 1 1310
box -12 -8 32 272
use FILL  FILL_6__1822_
timestamp 1701859473
transform -1 0 4770 0 -1 790
box -12 -8 32 272
use FILL  FILL_6__1823_
timestamp 1701859473
transform -1 0 4310 0 -1 790
box -12 -8 32 272
use FILL  FILL_6__1824_
timestamp 1701859473
transform 1 0 4690 0 1 2350
box -12 -8 32 272
use FILL  FILL_6__1825_
timestamp 1701859473
transform 1 0 5750 0 1 1830
box -12 -8 32 272
use FILL  FILL_6__1826_
timestamp 1701859473
transform 1 0 8250 0 -1 270
box -12 -8 32 272
use FILL  FILL_6__1827_
timestamp 1701859473
transform 1 0 9390 0 -1 790
box -12 -8 32 272
use FILL  FILL_6__1828_
timestamp 1701859473
transform 1 0 8550 0 1 270
box -12 -8 32 272
use FILL  FILL_6__1829_
timestamp 1701859473
transform 1 0 5850 0 1 270
box -12 -8 32 272
use FILL  FILL_6__1830_
timestamp 1701859473
transform 1 0 3290 0 1 4430
box -12 -8 32 272
use FILL  FILL_6__1831_
timestamp 1701859473
transform -1 0 8070 0 -1 790
box -12 -8 32 272
use FILL  FILL_6__1832_
timestamp 1701859473
transform 1 0 6570 0 -1 790
box -12 -8 32 272
use FILL  FILL_6__1833_
timestamp 1701859473
transform -1 0 770 0 1 270
box -12 -8 32 272
use FILL  FILL_6__1834_
timestamp 1701859473
transform 1 0 1210 0 -1 1310
box -12 -8 32 272
use FILL  FILL_6__1835_
timestamp 1701859473
transform -1 0 2590 0 -1 1310
box -12 -8 32 272
use FILL  FILL_6__1836_
timestamp 1701859473
transform 1 0 1150 0 1 790
box -12 -8 32 272
use FILL  FILL_6__1837_
timestamp 1701859473
transform -1 0 2550 0 1 790
box -12 -8 32 272
use FILL  FILL_6__1838_
timestamp 1701859473
transform 1 0 2290 0 1 790
box -12 -8 32 272
use FILL  FILL_6__1839_
timestamp 1701859473
transform -1 0 350 0 1 270
box -12 -8 32 272
use FILL  FILL_6__1840_
timestamp 1701859473
transform -1 0 990 0 1 2870
box -12 -8 32 272
use FILL  FILL_6__1841_
timestamp 1701859473
transform 1 0 3770 0 1 2870
box -12 -8 32 272
use FILL  FILL_6__1842_
timestamp 1701859473
transform -1 0 3030 0 -1 1830
box -12 -8 32 272
use FILL  FILL_6__1843_
timestamp 1701859473
transform -1 0 3990 0 -1 2350
box -12 -8 32 272
use FILL  FILL_6__1844_
timestamp 1701859473
transform 1 0 3890 0 -1 2870
box -12 -8 32 272
use FILL  FILL_6__1845_
timestamp 1701859473
transform -1 0 1830 0 -1 4950
box -12 -8 32 272
use FILL  FILL_6__1846_
timestamp 1701859473
transform 1 0 4190 0 1 4430
box -12 -8 32 272
use FILL  FILL_6__1847_
timestamp 1701859473
transform 1 0 3510 0 1 4430
box -12 -8 32 272
use FILL  FILL_6__1848_
timestamp 1701859473
transform 1 0 3950 0 1 4430
box -12 -8 32 272
use FILL  FILL_6__1849_
timestamp 1701859473
transform -1 0 4150 0 -1 2870
box -12 -8 32 272
use FILL  FILL_6__1850_
timestamp 1701859473
transform -1 0 970 0 1 790
box -12 -8 32 272
use FILL  FILL_6__1851_
timestamp 1701859473
transform 1 0 1630 0 -1 1830
box -12 -8 32 272
use FILL  FILL_6__1852_
timestamp 1701859473
transform -1 0 2450 0 1 2350
box -12 -8 32 272
use FILL  FILL_6__1853_
timestamp 1701859473
transform 1 0 130 0 -1 2350
box -12 -8 32 272
use FILL  FILL_6__1854_
timestamp 1701859473
transform 1 0 2370 0 -1 2350
box -12 -8 32 272
use FILL  FILL_6__1855_
timestamp 1701859473
transform -1 0 2630 0 -1 2350
box -12 -8 32 272
use FILL  FILL_6__1856_
timestamp 1701859473
transform 1 0 1530 0 -1 790
box -12 -8 32 272
use FILL  FILL_6__1857_
timestamp 1701859473
transform -1 0 2730 0 -1 790
box -12 -8 32 272
use FILL  FILL_6__1858_
timestamp 1701859473
transform 1 0 2470 0 -1 790
box -12 -8 32 272
use FILL  FILL_6__1859_
timestamp 1701859473
transform 1 0 2250 0 -1 790
box -12 -8 32 272
use FILL  FILL_6__1860_
timestamp 1701859473
transform -1 0 1790 0 -1 790
box -12 -8 32 272
use FILL  FILL_6__1861_
timestamp 1701859473
transform -1 0 2030 0 -1 790
box -12 -8 32 272
use FILL  FILL_6__1862_
timestamp 1701859473
transform -1 0 2110 0 1 270
box -12 -8 32 272
use FILL  FILL_6__1863_
timestamp 1701859473
transform 1 0 2330 0 1 270
box -12 -8 32 272
use FILL  FILL_6__1864_
timestamp 1701859473
transform 1 0 3570 0 1 270
box -12 -8 32 272
use FILL  FILL_6__1865_
timestamp 1701859473
transform 1 0 7370 0 -1 1310
box -12 -8 32 272
use FILL  FILL_6__1866_
timestamp 1701859473
transform 1 0 3730 0 -1 1310
box -12 -8 32 272
use FILL  FILL_6__1867_
timestamp 1701859473
transform 1 0 1190 0 -1 1830
box -12 -8 32 272
use FILL  FILL_6__1868_
timestamp 1701859473
transform 1 0 1630 0 1 1310
box -12 -8 32 272
use FILL  FILL_6__1869_
timestamp 1701859473
transform 1 0 2050 0 1 1310
box -12 -8 32 272
use FILL  FILL_6__1870_
timestamp 1701859473
transform -1 0 1670 0 -1 1310
box -12 -8 32 272
use FILL  FILL_6__1871_
timestamp 1701859473
transform -1 0 2790 0 -1 1310
box -12 -8 32 272
use FILL  FILL_6__1872_
timestamp 1701859473
transform -1 0 570 0 1 790
box -12 -8 32 272
use FILL  FILL_6__1873_
timestamp 1701859473
transform 1 0 750 0 1 790
box -12 -8 32 272
use FILL  FILL_6__1874_
timestamp 1701859473
transform -1 0 1390 0 1 790
box -12 -8 32 272
use FILL  FILL_6__1875_
timestamp 1701859473
transform 1 0 970 0 -1 790
box -12 -8 32 272
use FILL  FILL_6__1876_
timestamp 1701859473
transform 1 0 1290 0 -1 790
box -12 -8 32 272
use FILL  FILL_6__1877_
timestamp 1701859473
transform 1 0 2230 0 1 4950
box -12 -8 32 272
use FILL  FILL_6__1878_
timestamp 1701859473
transform 1 0 570 0 -1 1310
box -12 -8 32 272
use FILL  FILL_6__1879_
timestamp 1701859473
transform 1 0 790 0 1 1310
box -12 -8 32 272
use FILL  FILL_6__1880_
timestamp 1701859473
transform -1 0 2050 0 -1 4950
box -12 -8 32 272
use FILL  FILL_6__1881_
timestamp 1701859473
transform -1 0 2290 0 -1 4950
box -12 -8 32 272
use FILL  FILL_6__1882_
timestamp 1701859473
transform 1 0 1610 0 -1 3390
box -12 -8 32 272
use FILL  FILL_6__1883_
timestamp 1701859473
transform 1 0 1090 0 -1 3390
box -12 -8 32 272
use FILL  FILL_6__1884_
timestamp 1701859473
transform -1 0 4110 0 1 3390
box -12 -8 32 272
use FILL  FILL_6__1885_
timestamp 1701859473
transform -1 0 3830 0 -1 3390
box -12 -8 32 272
use FILL  FILL_6__1886_
timestamp 1701859473
transform 1 0 3570 0 -1 3390
box -12 -8 32 272
use FILL  FILL_6__1887_
timestamp 1701859473
transform -1 0 3550 0 1 2870
box -12 -8 32 272
use FILL  FILL_6__1888_
timestamp 1701859473
transform -1 0 2590 0 1 270
box -12 -8 32 272
use FILL  FILL_6__1889_
timestamp 1701859473
transform 1 0 1730 0 -1 2870
box -12 -8 32 272
use FILL  FILL_6__1890_
timestamp 1701859473
transform -1 0 370 0 -1 1830
box -12 -8 32 272
use FILL  FILL_6__1891_
timestamp 1701859473
transform 1 0 130 0 -1 1830
box -12 -8 32 272
use FILL  FILL_6__1892_
timestamp 1701859473
transform 1 0 4970 0 -1 3390
box -12 -8 32 272
use FILL  FILL_6__1893_
timestamp 1701859473
transform 1 0 3970 0 1 1830
box -12 -8 32 272
use FILL  FILL_6__1894_
timestamp 1701859473
transform 1 0 4170 0 1 1830
box -12 -8 32 272
use FILL  FILL_6__1895_
timestamp 1701859473
transform -1 0 1910 0 1 1830
box -12 -8 32 272
use FILL  FILL_6__1896_
timestamp 1701859473
transform 1 0 1930 0 -1 2350
box -12 -8 32 272
use FILL  FILL_6__1897_
timestamp 1701859473
transform 1 0 3550 0 1 2350
box -12 -8 32 272
use FILL  FILL_6__1898_
timestamp 1701859473
transform 1 0 3330 0 1 2350
box -12 -8 32 272
use FILL  FILL_6__1899_
timestamp 1701859473
transform -1 0 3310 0 -1 2350
box -12 -8 32 272
use FILL  FILL_6__1900_
timestamp 1701859473
transform -1 0 4150 0 -1 1830
box -12 -8 32 272
use FILL  FILL_6__1901_
timestamp 1701859473
transform -1 0 790 0 1 1830
box -12 -8 32 272
use FILL  FILL_6__1902_
timestamp 1701859473
transform 1 0 5090 0 1 1830
box -12 -8 32 272
use FILL  FILL_6__1903_
timestamp 1701859473
transform 1 0 3410 0 1 1310
box -12 -8 32 272
use FILL  FILL_6__1904_
timestamp 1701859473
transform -1 0 3510 0 -1 1310
box -12 -8 32 272
use FILL  FILL_6__1905_
timestamp 1701859473
transform 1 0 3050 0 1 270
box -12 -8 32 272
use FILL  FILL_6__1906_
timestamp 1701859473
transform 1 0 330 0 1 2350
box -12 -8 32 272
use FILL  FILL_6__1907_
timestamp 1701859473
transform -1 0 3090 0 -1 2350
box -12 -8 32 272
use FILL  FILL_6__1908_
timestamp 1701859473
transform 1 0 6510 0 -1 2350
box -12 -8 32 272
use FILL  FILL_6__1909_
timestamp 1701859473
transform -1 0 6110 0 -1 2350
box -12 -8 32 272
use FILL  FILL_6__1910_
timestamp 1701859473
transform -1 0 5610 0 -1 2350
box -12 -8 32 272
use FILL  FILL_6__1911_
timestamp 1701859473
transform -1 0 770 0 1 2870
box -12 -8 32 272
use FILL  FILL_6__1912_
timestamp 1701859473
transform -1 0 3370 0 1 3910
box -12 -8 32 272
use FILL  FILL_6__1913_
timestamp 1701859473
transform -1 0 1090 0 -1 2870
box -12 -8 32 272
use FILL  FILL_6__1914_
timestamp 1701859473
transform -1 0 1530 0 1 3390
box -12 -8 32 272
use FILL  FILL_6__1915_
timestamp 1701859473
transform 1 0 2610 0 1 3390
box -12 -8 32 272
use FILL  FILL_6__1916_
timestamp 1701859473
transform -1 0 3470 0 1 3390
box -12 -8 32 272
use FILL  FILL_6__1917_
timestamp 1701859473
transform -1 0 4750 0 -1 3390
box -12 -8 32 272
use FILL  FILL_6__1918_
timestamp 1701859473
transform 1 0 1790 0 1 4950
box -12 -8 32 272
use FILL  FILL_6__1919_
timestamp 1701859473
transform -1 0 1310 0 -1 2870
box -12 -8 32 272
use FILL  FILL_6__1920_
timestamp 1701859473
transform -1 0 5090 0 1 4430
box -12 -8 32 272
use FILL  FILL_6__1921_
timestamp 1701859473
transform 1 0 4850 0 1 4430
box -12 -8 32 272
use FILL  FILL_6__1922_
timestamp 1701859473
transform -1 0 4650 0 1 4430
box -12 -8 32 272
use FILL  FILL_6__1923_
timestamp 1701859473
transform 1 0 4510 0 -1 3390
box -12 -8 32 272
use FILL  FILL_6__1924_
timestamp 1701859473
transform 1 0 2010 0 1 4950
box -12 -8 32 272
use FILL  FILL_6__1925_
timestamp 1701859473
transform 1 0 6150 0 -1 4430
box -12 -8 32 272
use FILL  FILL_6__1926_
timestamp 1701859473
transform 1 0 770 0 -1 1310
box -12 -8 32 272
use FILL  FILL_6__1927_
timestamp 1701859473
transform 1 0 3010 0 -1 1310
box -12 -8 32 272
use FILL  FILL_6__1928_
timestamp 1701859473
transform -1 0 3270 0 -1 1310
box -12 -8 32 272
use FILL  FILL_6__1929_
timestamp 1701859473
transform 1 0 3450 0 1 790
box -12 -8 32 272
use FILL  FILL_6__1930_
timestamp 1701859473
transform 1 0 3270 0 1 270
box -12 -8 32 272
use FILL  FILL_6__1931_
timestamp 1701859473
transform 1 0 3870 0 1 270
box -12 -8 32 272
use FILL  FILL_6__1932_
timestamp 1701859473
transform -1 0 4110 0 1 270
box -12 -8 32 272
use FILL  FILL_6__1933_
timestamp 1701859473
transform -1 0 1910 0 1 270
box -12 -8 32 272
use FILL  FILL_6__1934_
timestamp 1701859473
transform -1 0 5530 0 1 790
box -12 -8 32 272
use FILL  FILL_6__1935_
timestamp 1701859473
transform 1 0 5650 0 -1 270
box -12 -8 32 272
use FILL  FILL_6__1936_
timestamp 1701859473
transform -1 0 8410 0 1 3390
box -12 -8 32 272
use FILL  FILL_6__1937_
timestamp 1701859473
transform -1 0 7630 0 -1 270
box -12 -8 32 272
use FILL  FILL_6__1938_
timestamp 1701859473
transform -1 0 7830 0 -1 270
box -12 -8 32 272
use FILL  FILL_6__1939_
timestamp 1701859473
transform -1 0 6750 0 -1 270
box -12 -8 32 272
use FILL  FILL_6__1940_
timestamp 1701859473
transform -1 0 5870 0 -1 270
box -12 -8 32 272
use FILL  FILL_6__1941_
timestamp 1701859473
transform 1 0 5890 0 -1 790
box -12 -8 32 272
use FILL  FILL_6__1942_
timestamp 1701859473
transform 1 0 4870 0 -1 1310
box -12 -8 32 272
use FILL  FILL_6__1943_
timestamp 1701859473
transform 1 0 8130 0 1 270
box -12 -8 32 272
use FILL  FILL_6__1944_
timestamp 1701859473
transform -1 0 8370 0 1 270
box -12 -8 32 272
use FILL  FILL_6__1945_
timestamp 1701859473
transform 1 0 7910 0 1 270
box -12 -8 32 272
use FILL  FILL_6__1946_
timestamp 1701859473
transform -1 0 6110 0 1 270
box -12 -8 32 272
use FILL  FILL_6__1947_
timestamp 1701859473
transform -1 0 6130 0 -1 790
box -12 -8 32 272
use FILL  FILL_6__1948_
timestamp 1701859473
transform 1 0 5410 0 -1 790
box -12 -8 32 272
use FILL  FILL_6__1949_
timestamp 1701859473
transform 1 0 4650 0 -1 1310
box -12 -8 32 272
use FILL  FILL_6__1950_
timestamp 1701859473
transform -1 0 8290 0 -1 790
box -12 -8 32 272
use FILL  FILL_6__1951_
timestamp 1701859473
transform 1 0 570 0 -1 2350
box -12 -8 32 272
use FILL  FILL_6__1952_
timestamp 1701859473
transform -1 0 5750 0 1 2350
box -12 -8 32 272
use FILL  FILL_6__1953_
timestamp 1701859473
transform 1 0 5850 0 -1 2350
box -12 -8 32 272
use FILL  FILL_6__1954_
timestamp 1701859473
transform 1 0 8230 0 -1 1310
box -12 -8 32 272
use FILL  FILL_6__1955_
timestamp 1701859473
transform -1 0 8770 0 1 1310
box -12 -8 32 272
use FILL  FILL_6__1956_
timestamp 1701859473
transform -1 0 6310 0 -1 1310
box -12 -8 32 272
use FILL  FILL_6__1957_
timestamp 1701859473
transform -1 0 6070 0 -1 1310
box -12 -8 32 272
use FILL  FILL_6__1958_
timestamp 1701859473
transform 1 0 5330 0 -1 1310
box -12 -8 32 272
use FILL  FILL_6__1959_
timestamp 1701859473
transform 1 0 5770 0 -1 2870
box -12 -8 32 272
use FILL  FILL_6__1960_
timestamp 1701859473
transform -1 0 6210 0 -1 2870
box -12 -8 32 272
use FILL  FILL_6__1961_
timestamp 1701859473
transform -1 0 4470 0 1 2350
box -12 -8 32 272
use FILL  FILL_6__1962_
timestamp 1701859473
transform 1 0 5930 0 1 2350
box -12 -8 32 272
use FILL  FILL_6__1963_
timestamp 1701859473
transform 1 0 5390 0 1 1310
box -12 -8 32 272
use FILL  FILL_6__1964_
timestamp 1701859473
transform 1 0 9210 0 1 1310
box -12 -8 32 272
use FILL  FILL_6__1965_
timestamp 1701859473
transform 1 0 7610 0 1 790
box -12 -8 32 272
use FILL  FILL_6__1966_
timestamp 1701859473
transform -1 0 7730 0 1 270
box -12 -8 32 272
use FILL  FILL_6__1967_
timestamp 1701859473
transform -1 0 6790 0 1 270
box -12 -8 32 272
use FILL  FILL_6__1968_
timestamp 1701859473
transform 1 0 5570 0 -1 1310
box -12 -8 32 272
use FILL  FILL_6__1969_
timestamp 1701859473
transform 1 0 5770 0 1 2870
box -12 -8 32 272
use FILL  FILL_6__1970_
timestamp 1701859473
transform 1 0 5410 0 -1 3390
box -12 -8 32 272
use FILL  FILL_6__1971_
timestamp 1701859473
transform 1 0 5850 0 1 3910
box -12 -8 32 272
use FILL  FILL_6__1972_
timestamp 1701859473
transform 1 0 5790 0 1 4950
box -12 -8 32 272
use FILL  FILL_6__1973_
timestamp 1701859473
transform -1 0 6130 0 -1 3910
box -12 -8 32 272
use FILL  FILL_6__1974_
timestamp 1701859473
transform 1 0 6310 0 -1 3910
box -12 -8 32 272
use FILL  FILL_6__1975_
timestamp 1701859473
transform -1 0 6110 0 1 3910
box -12 -8 32 272
use FILL  FILL_6__1976_
timestamp 1701859473
transform -1 0 6570 0 -1 3910
box -12 -8 32 272
use FILL  FILL_6__1977_
timestamp 1701859473
transform 1 0 6890 0 1 2870
box -12 -8 32 272
use FILL  FILL_6__1978_
timestamp 1701859473
transform -1 0 6430 0 -1 2870
box -12 -8 32 272
use FILL  FILL_6__1979_
timestamp 1701859473
transform 1 0 6470 0 1 2870
box -12 -8 32 272
use FILL  FILL_6__1980_
timestamp 1701859473
transform 1 0 6670 0 1 2870
box -12 -8 32 272
use FILL  FILL_6__1981_
timestamp 1701859473
transform 1 0 6250 0 1 2870
box -12 -8 32 272
use FILL  FILL_6__1982_
timestamp 1701859473
transform -1 0 5710 0 -1 1830
box -12 -8 32 272
use FILL  FILL_6__1983_
timestamp 1701859473
transform -1 0 4810 0 -1 270
box -12 -8 32 272
use FILL  FILL_6__1984_
timestamp 1701859473
transform -1 0 6510 0 -1 1310
box -12 -8 32 272
use FILL  FILL_6__1985_
timestamp 1701859473
transform 1 0 5070 0 -1 1310
box -12 -8 32 272
use FILL  FILL_6__1986_
timestamp 1701859473
transform 1 0 8270 0 1 790
box -12 -8 32 272
use FILL  FILL_6__1987_
timestamp 1701859473
transform 1 0 6950 0 1 1310
box -12 -8 32 272
use FILL  FILL_6__1988_
timestamp 1701859473
transform -1 0 7410 0 1 1310
box -12 -8 32 272
use FILL  FILL_6__1989_
timestamp 1701859473
transform 1 0 2770 0 -1 5470
box -12 -8 32 272
use FILL  FILL_6__1990_
timestamp 1701859473
transform 1 0 2090 0 1 1830
box -12 -8 32 272
use FILL  FILL_6__1991_
timestamp 1701859473
transform -1 0 2810 0 1 1830
box -12 -8 32 272
use FILL  FILL_6__1992_
timestamp 1701859473
transform -1 0 4210 0 -1 2350
box -12 -8 32 272
use FILL  FILL_6__1993_
timestamp 1701859473
transform -1 0 4450 0 -1 2350
box -12 -8 32 272
use FILL  FILL_6__1994_
timestamp 1701859473
transform 1 0 2550 0 1 1830
box -12 -8 32 272
use FILL  FILL_6__1995_
timestamp 1701859473
transform 1 0 3030 0 1 1830
box -12 -8 32 272
use FILL  FILL_6__1996_
timestamp 1701859473
transform -1 0 6710 0 1 790
box -12 -8 32 272
use FILL  FILL_6__1997_
timestamp 1701859473
transform -1 0 5050 0 1 790
box -12 -8 32 272
use FILL  FILL_6__1998_
timestamp 1701859473
transform 1 0 4310 0 1 270
box -12 -8 32 272
use FILL  FILL_6__1999_
timestamp 1701859473
transform -1 0 3910 0 -1 270
box -12 -8 32 272
use FILL  FILL_6__2000_
timestamp 1701859473
transform -1 0 4590 0 -1 270
box -12 -8 32 272
use FILL  FILL_6__2001_
timestamp 1701859473
transform -1 0 5970 0 -1 2870
box -12 -8 32 272
use FILL  FILL_6__2002_
timestamp 1701859473
transform -1 0 1910 0 1 2870
box -12 -8 32 272
use FILL  FILL_6__2003_
timestamp 1701859473
transform 1 0 1410 0 -1 3390
box -12 -8 32 272
use FILL  FILL_6__2004_
timestamp 1701859473
transform 1 0 2830 0 -1 3390
box -12 -8 32 272
use FILL  FILL_6__2005_
timestamp 1701859473
transform -1 0 3110 0 1 2870
box -12 -8 32 272
use FILL  FILL_6__2006_
timestamp 1701859473
transform 1 0 2850 0 1 2870
box -12 -8 32 272
use FILL  FILL_6__2007_
timestamp 1701859473
transform 1 0 6870 0 -1 2870
box -12 -8 32 272
use FILL  FILL_6__2008_
timestamp 1701859473
transform 1 0 550 0 -1 1830
box -12 -8 32 272
use FILL  FILL_6__2009_
timestamp 1701859473
transform -1 0 4070 0 -1 3390
box -12 -8 32 272
use FILL  FILL_6__2010_
timestamp 1701859473
transform -1 0 4370 0 -1 2870
box -12 -8 32 272
use FILL  FILL_6__2011_
timestamp 1701859473
transform -1 0 2110 0 1 790
box -12 -8 32 272
use FILL  FILL_6__2012_
timestamp 1701859473
transform 1 0 1610 0 1 790
box -12 -8 32 272
use FILL  FILL_6__2013_
timestamp 1701859473
transform -1 0 1870 0 1 790
box -12 -8 32 272
use FILL  FILL_6__2014_
timestamp 1701859473
transform 1 0 4530 0 1 1310
box -12 -8 32 272
use FILL  FILL_6__2015_
timestamp 1701859473
transform 1 0 3250 0 1 1830
box -12 -8 32 272
use FILL  FILL_6__2016_
timestamp 1701859473
transform -1 0 3750 0 1 1830
box -12 -8 32 272
use FILL  FILL_6__2017_
timestamp 1701859473
transform -1 0 5270 0 -1 1830
box -12 -8 32 272
use FILL  FILL_6__2018_
timestamp 1701859473
transform 1 0 5030 0 -1 1830
box -12 -8 32 272
use FILL  FILL_6__2019_
timestamp 1701859473
transform -1 0 5550 0 -1 2870
box -12 -8 32 272
use FILL  FILL_6__2020_
timestamp 1701859473
transform -1 0 5310 0 -1 2870
box -12 -8 32 272
use FILL  FILL_6__2021_
timestamp 1701859473
transform -1 0 6950 0 -1 1310
box -12 -8 32 272
use FILL  FILL_6__2022_
timestamp 1701859473
transform -1 0 7190 0 1 790
box -12 -8 32 272
use FILL  FILL_6__2023_
timestamp 1701859473
transform 1 0 8230 0 1 1830
box -12 -8 32 272
use FILL  FILL_6__2024_
timestamp 1701859473
transform -1 0 8450 0 1 1830
box -12 -8 32 272
use FILL  FILL_6__2025_
timestamp 1701859473
transform 1 0 9610 0 -1 790
box -12 -8 32 272
use FILL  FILL_6__2026_
timestamp 1701859473
transform -1 0 8750 0 1 790
box -12 -8 32 272
use FILL  FILL_6__2027_
timestamp 1701859473
transform -1 0 6950 0 1 790
box -12 -8 32 272
use FILL  FILL_6__2028_
timestamp 1701859473
transform 1 0 7050 0 -1 790
box -12 -8 32 272
use FILL  FILL_6__2029_
timestamp 1701859473
transform 1 0 7490 0 1 270
box -12 -8 32 272
use FILL  FILL_6__2030_
timestamp 1701859473
transform -1 0 7170 0 -1 1310
box -12 -8 32 272
use FILL  FILL_6__2031_
timestamp 1701859473
transform 1 0 7490 0 -1 790
box -12 -8 32 272
use FILL  FILL_6__2032_
timestamp 1701859473
transform -1 0 8790 0 1 270
box -12 -8 32 272
use FILL  FILL_6__2033_
timestamp 1701859473
transform 1 0 8270 0 1 1310
box -12 -8 32 272
use FILL  FILL_6__2034_
timestamp 1701859473
transform -1 0 8950 0 -1 1310
box -12 -8 32 272
use FILL  FILL_6__2035_
timestamp 1701859473
transform -1 0 8530 0 1 790
box -12 -8 32 272
use FILL  FILL_6__2036_
timestamp 1701859473
transform -1 0 8690 0 -1 1830
box -12 -8 32 272
use FILL  FILL_6__2037_
timestamp 1701859473
transform -1 0 8750 0 -1 790
box -12 -8 32 272
use FILL  FILL_6__2038_
timestamp 1701859473
transform 1 0 8050 0 1 790
box -12 -8 32 272
use FILL  FILL_6__2039_
timestamp 1701859473
transform 1 0 7830 0 1 790
box -12 -8 32 272
use FILL  FILL_6__2040_
timestamp 1701859473
transform -1 0 7750 0 -1 790
box -12 -8 32 272
use FILL  FILL_6__2041_
timestamp 1701859473
transform -1 0 6970 0 -1 270
box -12 -8 32 272
use FILL  FILL_6__2042_
timestamp 1701859473
transform 1 0 8950 0 -1 790
box -12 -8 32 272
use FILL  FILL_6__2043_
timestamp 1701859473
transform 1 0 7270 0 1 270
box -12 -8 32 272
use FILL  FILL_6__2044_
timestamp 1701859473
transform 1 0 7010 0 1 270
box -12 -8 32 272
use FILL  FILL_6__2045_
timestamp 1701859473
transform -1 0 6330 0 1 270
box -12 -8 32 272
use FILL  FILL_6__2046_
timestamp 1701859473
transform 1 0 6510 0 -1 270
box -12 -8 32 272
use FILL  FILL_6__2047_
timestamp 1701859473
transform -1 0 6290 0 -1 270
box -12 -8 32 272
use FILL  FILL_6__2048_
timestamp 1701859473
transform -1 0 6090 0 -1 270
box -12 -8 32 272
use FILL  FILL_6__2049_
timestamp 1701859473
transform -1 0 7270 0 -1 790
box -12 -8 32 272
use FILL  FILL_6__2050_
timestamp 1701859473
transform 1 0 1510 0 -1 2870
box -12 -8 32 272
use FILL  FILL_6__2051_
timestamp 1701859473
transform 1 0 6310 0 -1 2350
box -12 -8 32 272
use FILL  FILL_6__2052_
timestamp 1701859473
transform -1 0 6210 0 1 790
box -12 -8 32 272
use FILL  FILL_6__2053_
timestamp 1701859473
transform -1 0 4430 0 1 1830
box -12 -8 32 272
use FILL  FILL_6__2054_
timestamp 1701859473
transform 1 0 2930 0 1 1310
box -12 -8 32 272
use FILL  FILL_6__2055_
timestamp 1701859473
transform -1 0 3190 0 1 1310
box -12 -8 32 272
use FILL  FILL_6__2056_
timestamp 1701859473
transform -1 0 1910 0 -1 1310
box -12 -8 32 272
use FILL  FILL_6__2057_
timestamp 1701859473
transform 1 0 2770 0 1 790
box -12 -8 32 272
use FILL  FILL_6__2058_
timestamp 1701859473
transform 1 0 3690 0 1 790
box -12 -8 32 272
use FILL  FILL_6__2059_
timestamp 1701859473
transform 1 0 3930 0 1 790
box -12 -8 32 272
use FILL  FILL_6__2060_
timestamp 1701859473
transform -1 0 4170 0 1 790
box -12 -8 32 272
use FILL  FILL_6__2061_
timestamp 1701859473
transform -1 0 3030 0 -1 270
box -12 -8 32 272
use FILL  FILL_6__2062_
timestamp 1701859473
transform 1 0 2810 0 1 270
box -12 -8 32 272
use FILL  FILL_6__2063_
timestamp 1701859473
transform 1 0 3190 0 -1 270
box -12 -8 32 272
use FILL  FILL_6__2064_
timestamp 1701859473
transform 1 0 3430 0 -1 270
box -12 -8 32 272
use FILL  FILL_6__2065_
timestamp 1701859473
transform -1 0 3670 0 -1 270
box -12 -8 32 272
use FILL  FILL_6__2066_
timestamp 1701859473
transform -1 0 5450 0 -1 270
box -12 -8 32 272
use FILL  FILL_6__2067_
timestamp 1701859473
transform 1 0 7390 0 1 790
box -12 -8 32 272
use FILL  FILL_6__2068_
timestamp 1701859473
transform 1 0 5950 0 1 790
box -12 -8 32 272
use FILL  FILL_6__2069_
timestamp 1701859473
transform 1 0 3430 0 -1 1830
box -12 -8 32 272
use FILL  FILL_6__2070_
timestamp 1701859473
transform -1 0 3910 0 -1 1830
box -12 -8 32 272
use FILL  FILL_6__2071_
timestamp 1701859473
transform -1 0 5750 0 1 790
box -12 -8 32 272
use FILL  FILL_6__2072_
timestamp 1701859473
transform -1 0 7810 0 1 1310
box -12 -8 32 272
use FILL  FILL_6__2073_
timestamp 1701859473
transform 1 0 6690 0 1 1310
box -12 -8 32 272
use FILL  FILL_6__2074_
timestamp 1701859473
transform 1 0 1830 0 1 1310
box -12 -8 32 272
use FILL  FILL_6__2075_
timestamp 1701859473
transform -1 0 2310 0 1 1310
box -12 -8 32 272
use FILL  FILL_6__2076_
timestamp 1701859473
transform -1 0 2350 0 -1 1310
box -12 -8 32 272
use FILL  FILL_6__2077_
timestamp 1701859473
transform 1 0 4210 0 -1 1310
box -12 -8 32 272
use FILL  FILL_6__2078_
timestamp 1701859473
transform -1 0 2350 0 1 1830
box -12 -8 32 272
use FILL  FILL_6__2079_
timestamp 1701859473
transform -1 0 990 0 -1 1830
box -12 -8 32 272
use FILL  FILL_6__2080_
timestamp 1701859473
transform 1 0 2310 0 -1 1830
box -12 -8 32 272
use FILL  FILL_6__2081_
timestamp 1701859473
transform 1 0 2550 0 -1 1830
box -12 -8 32 272
use FILL  FILL_6__2082_
timestamp 1701859473
transform -1 0 2770 0 -1 1830
box -12 -8 32 272
use FILL  FILL_6__2083_
timestamp 1701859473
transform 1 0 4450 0 -1 1310
box -12 -8 32 272
use FILL  FILL_6__2084_
timestamp 1701859473
transform -1 0 5290 0 1 790
box -12 -8 32 272
use FILL  FILL_6__2085_
timestamp 1701859473
transform -1 0 5130 0 -1 270
box -12 -8 32 272
use FILL  FILL_6__2086_
timestamp 1701859473
transform -1 0 4350 0 -1 270
box -12 -8 32 272
use FILL  FILL_6__2087_
timestamp 1701859473
transform -1 0 4830 0 1 790
box -12 -8 32 272
use FILL  FILL_6__2088_
timestamp 1701859473
transform -1 0 5670 0 1 270
box -12 -8 32 272
use FILL  FILL_6__2089_
timestamp 1701859473
transform 1 0 5430 0 1 270
box -12 -8 32 272
use FILL  FILL_6__2090_
timestamp 1701859473
transform -1 0 5010 0 -1 790
box -12 -8 32 272
use FILL  FILL_6__2091_
timestamp 1701859473
transform 1 0 3230 0 1 790
box -12 -8 32 272
use FILL  FILL_6__2092_
timestamp 1701859473
transform 1 0 2790 0 -1 270
box -12 -8 32 272
use FILL  FILL_6__2093_
timestamp 1701859473
transform -1 0 2950 0 -1 790
box -12 -8 32 272
use FILL  FILL_6__2094_
timestamp 1701859473
transform 1 0 2350 0 -1 270
box -12 -8 32 272
use FILL  FILL_6__2095_
timestamp 1701859473
transform 1 0 2550 0 -1 270
box -12 -8 32 272
use FILL  FILL_6__2096_
timestamp 1701859473
transform -1 0 5010 0 1 270
box -12 -8 32 272
use FILL  FILL_6__2097_
timestamp 1701859473
transform -1 0 5230 0 1 270
box -12 -8 32 272
use FILL  FILL_6__2098_
timestamp 1701859473
transform 1 0 4770 0 1 270
box -12 -8 32 272
use FILL  FILL_6__2099_
timestamp 1701859473
transform 1 0 4090 0 -1 270
box -12 -8 32 272
use FILL  FILL_6__2100_
timestamp 1701859473
transform -1 0 5950 0 -1 1830
box -12 -8 32 272
use FILL  FILL_6__2101_
timestamp 1701859473
transform -1 0 5870 0 1 1310
box -12 -8 32 272
use FILL  FILL_6__2102_
timestamp 1701859473
transform -1 0 6270 0 1 1310
box -12 -8 32 272
use FILL  FILL_6__2103_
timestamp 1701859473
transform 1 0 5830 0 -1 1310
box -12 -8 32 272
use FILL  FILL_6__2104_
timestamp 1701859473
transform -1 0 6070 0 1 1310
box -12 -8 32 272
use FILL  FILL_6__2105_
timestamp 1701859473
transform -1 0 4370 0 -1 1830
box -12 -8 32 272
use FILL  FILL_6__2106_
timestamp 1701859473
transform 1 0 4050 0 -1 790
box -12 -8 32 272
use FILL  FILL_6__2107_
timestamp 1701859473
transform -1 0 3630 0 -1 790
box -12 -8 32 272
use FILL  FILL_6__2108_
timestamp 1701859473
transform 1 0 2990 0 1 790
box -12 -8 32 272
use FILL  FILL_6__2109_
timestamp 1701859473
transform -1 0 3410 0 -1 790
box -12 -8 32 272
use FILL  FILL_6__2110_
timestamp 1701859473
transform 1 0 3170 0 -1 790
box -12 -8 32 272
use FILL  FILL_6__2111_
timestamp 1701859473
transform -1 0 3850 0 -1 790
box -12 -8 32 272
use FILL  FILL_6__2112_
timestamp 1701859473
transform -1 0 5210 0 -1 790
box -12 -8 32 272
use FILL  FILL_6__2113_
timestamp 1701859473
transform -1 0 5190 0 1 1310
box -12 -8 32 272
use FILL  FILL_6__2114_
timestamp 1701859473
transform -1 0 5630 0 1 1310
box -12 -8 32 272
use FILL  FILL_6__2115_
timestamp 1701859473
transform -1 0 5670 0 -1 790
box -12 -8 32 272
use FILL  FILL_6__2116_
timestamp 1701859473
transform 1 0 2490 0 1 1310
box -12 -8 32 272
use FILL  FILL_6__2117_
timestamp 1701859473
transform 1 0 2690 0 1 1310
box -12 -8 32 272
use FILL  FILL_6__2118_
timestamp 1701859473
transform 1 0 3870 0 1 1310
box -12 -8 32 272
use FILL  FILL_6__2119_
timestamp 1701859473
transform -1 0 4130 0 1 1310
box -12 -8 32 272
use FILL  FILL_6__2120_
timestamp 1701859473
transform 1 0 3990 0 -1 1310
box -12 -8 32 272
use FILL  FILL_6__2121_
timestamp 1701859473
transform -1 0 4570 0 1 270
box -12 -8 32 272
use FILL  FILL_6__2122_
timestamp 1701859473
transform -1 0 2910 0 1 2350
box -12 -8 32 272
use FILL  FILL_6__2123_
timestamp 1701859473
transform 1 0 2850 0 -1 2350
box -12 -8 32 272
use FILL  FILL_6__2124_
timestamp 1701859473
transform -1 0 3750 0 -1 2350
box -12 -8 32 272
use FILL  FILL_6__2125_
timestamp 1701859473
transform 1 0 5870 0 -1 3390
box -12 -8 32 272
use FILL  FILL_6__2126_
timestamp 1701859473
transform 1 0 5550 0 1 2870
box -12 -8 32 272
use FILL  FILL_6__2127_
timestamp 1701859473
transform -1 0 6030 0 1 2870
box -12 -8 32 272
use FILL  FILL_6__2128_
timestamp 1701859473
transform 1 0 4650 0 1 2870
box -12 -8 32 272
use FILL  FILL_6__2129_
timestamp 1701859473
transform 1 0 5330 0 1 2870
box -12 -8 32 272
use FILL  FILL_6__2130_
timestamp 1701859473
transform -1 0 4690 0 -1 2350
box -12 -8 32 272
use FILL  FILL_6__2131_
timestamp 1701859473
transform 1 0 4730 0 1 1310
box -12 -8 32 272
use FILL  FILL_6__2132_
timestamp 1701859473
transform -1 0 4610 0 1 790
box -12 -8 32 272
use FILL  FILL_6__2133_
timestamp 1701859473
transform 1 0 4530 0 -1 790
box -12 -8 32 272
use FILL  FILL_6__2134_
timestamp 1701859473
transform 1 0 3650 0 -1 2870
box -12 -8 32 272
use FILL  FILL_6__2135_
timestamp 1701859473
transform 1 0 4270 0 -1 3390
box -12 -8 32 272
use FILL  FILL_6__2136_
timestamp 1701859473
transform -1 0 2810 0 1 3390
box -12 -8 32 272
use FILL  FILL_6__2137_
timestamp 1701859473
transform 1 0 2370 0 1 3390
box -12 -8 32 272
use FILL  FILL_6__2138_
timestamp 1701859473
transform 1 0 3170 0 -1 4430
box -12 -8 32 272
use FILL  FILL_6__2139_
timestamp 1701859473
transform -1 0 2950 0 -1 4430
box -12 -8 32 272
use FILL  FILL_6__2140_
timestamp 1701859473
transform 1 0 2870 0 1 4430
box -12 -8 32 272
use FILL  FILL_6__2141_
timestamp 1701859473
transform -1 0 3110 0 1 4430
box -12 -8 32 272
use FILL  FILL_6__2142_
timestamp 1701859473
transform 1 0 2990 0 1 3390
box -12 -8 32 272
use FILL  FILL_6__2143_
timestamp 1701859473
transform -1 0 7490 0 -1 3390
box -12 -8 32 272
use FILL  FILL_6__2144_
timestamp 1701859473
transform 1 0 2130 0 1 2870
box -12 -8 32 272
use FILL  FILL_6__2145_
timestamp 1701859473
transform -1 0 10110 0 -1 2870
box -12 -8 32 272
use FILL  FILL_6__2146_
timestamp 1701859473
transform -1 0 7690 0 -1 3390
box -12 -8 32 272
use FILL  FILL_6__2147_
timestamp 1701859473
transform 1 0 7650 0 -1 3910
box -12 -8 32 272
use FILL  FILL_6__2148_
timestamp 1701859473
transform 1 0 7490 0 1 3390
box -12 -8 32 272
use FILL  FILL_6__2149_
timestamp 1701859473
transform 1 0 7690 0 1 3390
box -12 -8 32 272
use FILL  FILL_6__2150_
timestamp 1701859473
transform -1 0 7950 0 1 3390
box -12 -8 32 272
use FILL  FILL_6__2151_
timestamp 1701859473
transform 1 0 7230 0 -1 3390
box -12 -8 32 272
use FILL  FILL_6__2152_
timestamp 1701859473
transform 1 0 6990 0 -1 3390
box -12 -8 32 272
use FILL  FILL_6__2153_
timestamp 1701859473
transform -1 0 6130 0 -1 3390
box -12 -8 32 272
use FILL  FILL_6__2154_
timestamp 1701859473
transform 1 0 2890 0 -1 7030
box -12 -8 32 272
use FILL  FILL_6__2155_
timestamp 1701859473
transform 1 0 6450 0 1 5990
box -12 -8 32 272
use FILL  FILL_6__2156_
timestamp 1701859473
transform -1 0 4670 0 1 3910
box -12 -8 32 272
use FILL  FILL_6__2157_
timestamp 1701859473
transform -1 0 4810 0 -1 4430
box -12 -8 32 272
use FILL  FILL_6__2158_
timestamp 1701859473
transform -1 0 2670 0 1 2350
box -12 -8 32 272
use FILL  FILL_6__2159_
timestamp 1701859473
transform 1 0 3570 0 1 3910
box -12 -8 32 272
use FILL  FILL_6__2160_
timestamp 1701859473
transform -1 0 3890 0 -1 4430
box -12 -8 32 272
use FILL  FILL_6__2161_
timestamp 1701859473
transform -1 0 4030 0 1 3910
box -12 -8 32 272
use FILL  FILL_6__2162_
timestamp 1701859473
transform -1 0 4470 0 1 3910
box -12 -8 32 272
use FILL  FILL_6__2163_
timestamp 1701859473
transform 1 0 3790 0 -1 3910
box -12 -8 32 272
use FILL  FILL_6__2164_
timestamp 1701859473
transform -1 0 610 0 -1 4950
box -12 -8 32 272
use FILL  FILL_6__2165_
timestamp 1701859473
transform -1 0 3310 0 -1 3910
box -12 -8 32 272
use FILL  FILL_6__2166_
timestamp 1701859473
transform 1 0 4010 0 -1 3910
box -12 -8 32 272
use FILL  FILL_6__2167_
timestamp 1701859473
transform 1 0 4210 0 1 3910
box -12 -8 32 272
use FILL  FILL_6__2168_
timestamp 1701859473
transform 1 0 3130 0 1 3910
box -12 -8 32 272
use FILL  FILL_6__2169_
timestamp 1701859473
transform 1 0 2490 0 -1 4430
box -12 -8 32 272
use FILL  FILL_6__2170_
timestamp 1701859473
transform -1 0 2750 0 -1 4430
box -12 -8 32 272
use FILL  FILL_6__2171_
timestamp 1701859473
transform 1 0 4090 0 -1 4430
box -12 -8 32 272
use FILL  FILL_6__2172_
timestamp 1701859473
transform 1 0 4330 0 -1 4430
box -12 -8 32 272
use FILL  FILL_6__2173_
timestamp 1701859473
transform -1 0 4570 0 -1 4430
box -12 -8 32 272
use FILL  FILL_6__2174_
timestamp 1701859473
transform 1 0 6070 0 1 7030
box -12 -8 32 272
use FILL  FILL_6__2175_
timestamp 1701859473
transform -1 0 2570 0 1 8070
box -12 -8 32 272
use FILL  FILL_6__2176_
timestamp 1701859473
transform -1 0 6490 0 -1 8070
box -12 -8 32 272
use FILL  FILL_6__2177_
timestamp 1701859473
transform 1 0 5010 0 1 8070
box -12 -8 32 272
use FILL  FILL_6__2178_
timestamp 1701859473
transform -1 0 4190 0 -1 8590
box -12 -8 32 272
use FILL  FILL_6__2179_
timestamp 1701859473
transform -1 0 6010 0 -1 8070
box -12 -8 32 272
use FILL  FILL_6__2180_
timestamp 1701859473
transform -1 0 3030 0 -1 9630
box -12 -8 32 272
use FILL  FILL_6__2181_
timestamp 1701859473
transform 1 0 5090 0 1 7550
box -12 -8 32 272
use FILL  FILL_6__2182_
timestamp 1701859473
transform 1 0 5610 0 -1 10150
box -12 -8 32 272
use FILL  FILL_6__2183_
timestamp 1701859473
transform -1 0 3590 0 1 10150
box -12 -8 32 272
use FILL  FILL_6__2184_
timestamp 1701859473
transform 1 0 4410 0 1 8070
box -12 -8 32 272
use FILL  FILL_6__2185_
timestamp 1701859473
transform 1 0 6010 0 1 10150
box -12 -8 32 272
use FILL  FILL_6__2186_
timestamp 1701859473
transform 1 0 3570 0 1 10670
box -12 -8 32 272
use FILL  FILL_6__2187_
timestamp 1701859473
transform -1 0 5490 0 -1 10670
box -12 -8 32 272
use FILL  FILL_6__2188_
timestamp 1701859473
transform 1 0 2170 0 -1 10670
box -12 -8 32 272
use FILL  FILL_6__2189_
timestamp 1701859473
transform 1 0 5730 0 -1 10670
box -12 -8 32 272
use FILL  FILL_6__2190_
timestamp 1701859473
transform -1 0 2890 0 1 10150
box -12 -8 32 272
use FILL  FILL_6__2191_
timestamp 1701859473
transform -1 0 5370 0 -1 10150
box -12 -8 32 272
use FILL  FILL_6__2192_
timestamp 1701859473
transform -1 0 11170 0 1 3910
box -12 -8 32 272
use FILL  FILL_6__2193_
timestamp 1701859473
transform 1 0 1290 0 -1 3910
box -12 -8 32 272
use FILL  FILL_6__2194_
timestamp 1701859473
transform 1 0 1090 0 -1 3910
box -12 -8 32 272
use FILL  FILL_6__2195_
timestamp 1701859473
transform 1 0 2670 0 1 3910
box -12 -8 32 272
use FILL  FILL_6__2196_
timestamp 1701859473
transform 1 0 2910 0 1 3910
box -12 -8 32 272
use FILL  FILL_6__2197_
timestamp 1701859473
transform 1 0 5390 0 1 3910
box -12 -8 32 272
use FILL  FILL_6__2198_
timestamp 1701859473
transform 1 0 330 0 1 1830
box -12 -8 32 272
use FILL  FILL_6__2199_
timestamp 1701859473
transform -1 0 2890 0 -1 3910
box -12 -8 32 272
use FILL  FILL_6__2200_
timestamp 1701859473
transform 1 0 5410 0 -1 3910
box -12 -8 32 272
use FILL  FILL_6__2201_
timestamp 1701859473
transform -1 0 5650 0 1 3910
box -12 -8 32 272
use FILL  FILL_6__2202_
timestamp 1701859473
transform -1 0 8230 0 -1 4430
box -12 -8 32 272
use FILL  FILL_6__2203_
timestamp 1701859473
transform -1 0 4950 0 -1 3910
box -12 -8 32 272
use FILL  FILL_6__2204_
timestamp 1701859473
transform 1 0 5170 0 -1 3910
box -12 -8 32 272
use FILL  FILL_6__2205_
timestamp 1701859473
transform -1 0 9030 0 -1 3910
box -12 -8 32 272
use FILL  FILL_6__2206_
timestamp 1701859473
transform 1 0 9110 0 1 3910
box -12 -8 32 272
use FILL  FILL_6__2207_
timestamp 1701859473
transform 1 0 9570 0 -1 3910
box -12 -8 32 272
use FILL  FILL_6__2208_
timestamp 1701859473
transform -1 0 9830 0 -1 3910
box -12 -8 32 272
use FILL  FILL_6__2209_
timestamp 1701859473
transform -1 0 9630 0 1 4430
box -12 -8 32 272
use FILL  FILL_6__2210_
timestamp 1701859473
transform -1 0 10630 0 -1 4950
box -12 -8 32 272
use FILL  FILL_6__2211_
timestamp 1701859473
transform 1 0 9330 0 -1 3910
box -12 -8 32 272
use FILL  FILL_6__2212_
timestamp 1701859473
transform -1 0 8910 0 1 3910
box -12 -8 32 272
use FILL  FILL_6__2213_
timestamp 1701859473
transform -1 0 9350 0 1 3910
box -12 -8 32 272
use FILL  FILL_6__2214_
timestamp 1701859473
transform -1 0 9550 0 -1 4430
box -12 -8 32 272
use FILL  FILL_6__2215_
timestamp 1701859473
transform 1 0 9750 0 -1 4430
box -12 -8 32 272
use FILL  FILL_6__2216_
timestamp 1701859473
transform -1 0 9510 0 -1 7030
box -12 -8 32 272
use FILL  FILL_6__2217_
timestamp 1701859473
transform 1 0 9290 0 -1 4430
box -12 -8 32 272
use FILL  FILL_6__2218_
timestamp 1701859473
transform -1 0 9810 0 1 3910
box -12 -8 32 272
use FILL  FILL_6__2219_
timestamp 1701859473
transform 1 0 9990 0 1 3910
box -12 -8 32 272
use FILL  FILL_6__2220_
timestamp 1701859473
transform 1 0 10370 0 -1 4950
box -12 -8 32 272
use FILL  FILL_6__2221_
timestamp 1701859473
transform -1 0 9750 0 -1 7030
box -12 -8 32 272
use FILL  FILL_6__2222_
timestamp 1701859473
transform 1 0 10110 0 1 4430
box -12 -8 32 272
use FILL  FILL_6__2223_
timestamp 1701859473
transform -1 0 10010 0 -1 4430
box -12 -8 32 272
use FILL  FILL_6__2224_
timestamp 1701859473
transform -1 0 9870 0 1 4430
box -12 -8 32 272
use FILL  FILL_6__2225_
timestamp 1701859473
transform 1 0 10110 0 -1 4950
box -12 -8 32 272
use FILL  FILL_6__2226_
timestamp 1701859473
transform 1 0 8990 0 -1 7030
box -12 -8 32 272
use FILL  FILL_6__2227_
timestamp 1701859473
transform -1 0 9270 0 -1 7030
box -12 -8 32 272
use FILL  FILL_6__2228_
timestamp 1701859473
transform -1 0 5810 0 -1 7030
box -12 -8 32 272
use FILL  FILL_6__2229_
timestamp 1701859473
transform 1 0 4370 0 1 3390
box -12 -8 32 272
use FILL  FILL_6__2230_
timestamp 1701859473
transform -1 0 4470 0 -1 3910
box -12 -8 32 272
use FILL  FILL_6__2231_
timestamp 1701859473
transform -1 0 4250 0 -1 3910
box -12 -8 32 272
use FILL  FILL_6__2232_
timestamp 1701859473
transform 1 0 1650 0 1 2870
box -12 -8 32 272
use FILL  FILL_6__2233_
timestamp 1701859473
transform 1 0 2370 0 1 2870
box -12 -8 32 272
use FILL  FILL_6__2234_
timestamp 1701859473
transform -1 0 2630 0 1 2870
box -12 -8 32 272
use FILL  FILL_6__2235_
timestamp 1701859473
transform 1 0 6390 0 1 3390
box -12 -8 32 272
use FILL  FILL_6__2236_
timestamp 1701859473
transform -1 0 5670 0 -1 3910
box -12 -8 32 272
use FILL  FILL_6__2237_
timestamp 1701859473
transform -1 0 4710 0 -1 3910
box -12 -8 32 272
use FILL  FILL_6__2238_
timestamp 1701859473
transform 1 0 4770 0 -1 4950
box -12 -8 32 272
use FILL  FILL_6__2239_
timestamp 1701859473
transform 1 0 2890 0 1 4950
box -12 -8 32 272
use FILL  FILL_6__2240_
timestamp 1701859473
transform 1 0 2450 0 1 3910
box -12 -8 32 272
use FILL  FILL_6__2241_
timestamp 1701859473
transform -1 0 2470 0 1 4950
box -12 -8 32 272
use FILL  FILL_6__2242_
timestamp 1701859473
transform 1 0 2510 0 -1 4950
box -12 -8 32 272
use FILL  FILL_6__2243_
timestamp 1701859473
transform 1 0 2690 0 1 4950
box -12 -8 32 272
use FILL  FILL_6__2244_
timestamp 1701859473
transform 1 0 3110 0 1 4950
box -12 -8 32 272
use FILL  FILL_6__2245_
timestamp 1701859473
transform 1 0 2950 0 1 5990
box -12 -8 32 272
use FILL  FILL_6__2246_
timestamp 1701859473
transform 1 0 2970 0 -1 4950
box -12 -8 32 272
use FILL  FILL_6__2247_
timestamp 1701859473
transform -1 0 3090 0 -1 6510
box -12 -8 32 272
use FILL  FILL_6__2248_
timestamp 1701859473
transform 1 0 3550 0 -1 7030
box -12 -8 32 272
use FILL  FILL_6__2249_
timestamp 1701859473
transform 1 0 6330 0 1 7030
box -12 -8 32 272
use FILL  FILL_6__2250_
timestamp 1701859473
transform -1 0 10630 0 -1 7550
box -12 -8 32 272
use FILL  FILL_6__2251_
timestamp 1701859473
transform -1 0 10690 0 1 8070
box -12 -8 32 272
use FILL  FILL_6__2252_
timestamp 1701859473
transform -1 0 10990 0 -1 8070
box -12 -8 32 272
use FILL  FILL_6__2253_
timestamp 1701859473
transform -1 0 10750 0 -1 8070
box -12 -8 32 272
use FILL  FILL_6__2254_
timestamp 1701859473
transform 1 0 5450 0 1 8070
box -12 -8 32 272
use FILL  FILL_6__2255_
timestamp 1701859473
transform 1 0 3070 0 1 7030
box -12 -8 32 272
use FILL  FILL_6__2256_
timestamp 1701859473
transform -1 0 5190 0 1 7030
box -12 -8 32 272
use FILL  FILL_6__2257_
timestamp 1701859473
transform 1 0 5130 0 -1 7550
box -12 -8 32 272
use FILL  FILL_6__2258_
timestamp 1701859473
transform 1 0 5770 0 -1 8590
box -12 -8 32 272
use FILL  FILL_6__2259_
timestamp 1701859473
transform 1 0 10390 0 -1 7550
box -12 -8 32 272
use FILL  FILL_6__2260_
timestamp 1701859473
transform 1 0 9970 0 1 8070
box -12 -8 32 272
use FILL  FILL_6__2261_
timestamp 1701859473
transform -1 0 10270 0 1 7550
box -12 -8 32 272
use FILL  FILL_6__2262_
timestamp 1701859473
transform -1 0 10030 0 1 7550
box -12 -8 32 272
use FILL  FILL_6__2263_
timestamp 1701859473
transform 1 0 5530 0 1 7550
box -12 -8 32 272
use FILL  FILL_6__2264_
timestamp 1701859473
transform 1 0 1690 0 -1 6510
box -12 -8 32 272
use FILL  FILL_6__2265_
timestamp 1701859473
transform 1 0 1870 0 -1 6510
box -12 -8 32 272
use FILL  FILL_6__2266_
timestamp 1701859473
transform 1 0 3970 0 1 6510
box -12 -8 32 272
use FILL  FILL_6__2267_
timestamp 1701859473
transform -1 0 3730 0 -1 7550
box -12 -8 32 272
use FILL  FILL_6__2268_
timestamp 1701859473
transform 1 0 4410 0 -1 7550
box -12 -8 32 272
use FILL  FILL_6__2269_
timestamp 1701859473
transform 1 0 5730 0 1 7550
box -12 -8 32 272
use FILL  FILL_6__2270_
timestamp 1701859473
transform 1 0 8650 0 1 7550
box -12 -8 32 272
use FILL  FILL_6__2271_
timestamp 1701859473
transform -1 0 8930 0 -1 8070
box -12 -8 32 272
use FILL  FILL_6__2272_
timestamp 1701859473
transform -1 0 9190 0 -1 8070
box -12 -8 32 272
use FILL  FILL_6__2273_
timestamp 1701859473
transform -1 0 8690 0 -1 8070
box -12 -8 32 272
use FILL  FILL_6__2274_
timestamp 1701859473
transform -1 0 6050 0 -1 9630
box -12 -8 32 272
use FILL  FILL_6__2275_
timestamp 1701859473
transform -1 0 2350 0 1 8070
box -12 -8 32 272
use FILL  FILL_6__2276_
timestamp 1701859473
transform -1 0 3230 0 1 8070
box -12 -8 32 272
use FILL  FILL_6__2277_
timestamp 1701859473
transform -1 0 3710 0 -1 8590
box -12 -8 32 272
use FILL  FILL_6__2278_
timestamp 1701859473
transform 1 0 6610 0 1 9110
box -12 -8 32 272
use FILL  FILL_6__2279_
timestamp 1701859473
transform -1 0 10310 0 1 5990
box -12 -8 32 272
use FILL  FILL_6__2280_
timestamp 1701859473
transform 1 0 10490 0 1 5990
box -12 -8 32 272
use FILL  FILL_6__2281_
timestamp 1701859473
transform -1 0 10770 0 -1 5990
box -12 -8 32 272
use FILL  FILL_6__2282_
timestamp 1701859473
transform -1 0 10550 0 -1 6510
box -12 -8 32 272
use FILL  FILL_6__2283_
timestamp 1701859473
transform 1 0 6010 0 -1 8590
box -12 -8 32 272
use FILL  FILL_6__2284_
timestamp 1701859473
transform -1 0 2130 0 1 8070
box -12 -8 32 272
use FILL  FILL_6__2285_
timestamp 1701859473
transform -1 0 4190 0 1 8070
box -12 -8 32 272
use FILL  FILL_6__2286_
timestamp 1701859473
transform 1 0 5090 0 -1 8590
box -12 -8 32 272
use FILL  FILL_6__2287_
timestamp 1701859473
transform -1 0 6170 0 1 8590
box -12 -8 32 272
use FILL  FILL_6__2288_
timestamp 1701859473
transform -1 0 8890 0 1 7550
box -12 -8 32 272
use FILL  FILL_6__2289_
timestamp 1701859473
transform 1 0 8550 0 1 8070
box -12 -8 32 272
use FILL  FILL_6__2290_
timestamp 1701859473
transform -1 0 10050 0 -1 8070
box -12 -8 32 272
use FILL  FILL_6__2291_
timestamp 1701859473
transform -1 0 8830 0 1 8070
box -12 -8 32 272
use FILL  FILL_6__2292_
timestamp 1701859473
transform -1 0 6270 0 -1 9110
box -12 -8 32 272
use FILL  FILL_6__2293_
timestamp 1701859473
transform -1 0 2590 0 -1 8590
box -12 -8 32 272
use FILL  FILL_6__2294_
timestamp 1701859473
transform -1 0 4070 0 1 8590
box -12 -8 32 272
use FILL  FILL_6__2295_
timestamp 1701859473
transform 1 0 4990 0 1 8590
box -12 -8 32 272
use FILL  FILL_6__2296_
timestamp 1701859473
transform 1 0 6710 0 -1 9110
box -12 -8 32 272
use FILL  FILL_6__2297_
timestamp 1701859473
transform -1 0 9610 0 -1 5990
box -12 -8 32 272
use FILL  FILL_6__2298_
timestamp 1701859473
transform -1 0 10050 0 -1 5470
box -12 -8 32 272
use FILL  FILL_6__2299_
timestamp 1701859473
transform -1 0 9390 0 -1 6510
box -12 -8 32 272
use FILL  FILL_6__2300_
timestamp 1701859473
transform 1 0 9590 0 1 5990
box -12 -8 32 272
use FILL  FILL_6__2301_
timestamp 1701859473
transform 1 0 5630 0 1 9630
box -12 -8 32 272
use FILL  FILL_6__2302_
timestamp 1701859473
transform -1 0 3530 0 -1 9110
box -12 -8 32 272
use FILL  FILL_6__2303_
timestamp 1701859473
transform 1 0 2650 0 1 9110
box -12 -8 32 272
use FILL  FILL_6__2304_
timestamp 1701859473
transform 1 0 2850 0 -1 9110
box -12 -8 32 272
use FILL  FILL_6__2305_
timestamp 1701859473
transform -1 0 3830 0 1 8590
box -12 -8 32 272
use FILL  FILL_6__2306_
timestamp 1701859473
transform 1 0 4510 0 1 8590
box -12 -8 32 272
use FILL  FILL_6__2307_
timestamp 1701859473
transform 1 0 6370 0 1 9110
box -12 -8 32 272
use FILL  FILL_6__2308_
timestamp 1701859473
transform -1 0 8950 0 -1 6510
box -12 -8 32 272
use FILL  FILL_6__2309_
timestamp 1701859473
transform -1 0 8650 0 1 5990
box -12 -8 32 272
use FILL  FILL_6__2310_
timestamp 1701859473
transform -1 0 9150 0 -1 6510
box -12 -8 32 272
use FILL  FILL_6__2311_
timestamp 1701859473
transform -1 0 8710 0 -1 6510
box -12 -8 32 272
use FILL  FILL_6__2312_
timestamp 1701859473
transform -1 0 5610 0 -1 9630
box -12 -8 32 272
use FILL  FILL_6__2313_
timestamp 1701859473
transform -1 0 1890 0 1 8590
box -12 -8 32 272
use FILL  FILL_6__2314_
timestamp 1701859473
transform 1 0 1490 0 -1 8590
box -12 -8 32 272
use FILL  FILL_6__2315_
timestamp 1701859473
transform 1 0 1930 0 -1 8590
box -12 -8 32 272
use FILL  FILL_6__2316_
timestamp 1701859473
transform -1 0 4290 0 1 8590
box -12 -8 32 272
use FILL  FILL_6__2317_
timestamp 1701859473
transform 1 0 4750 0 1 8590
box -12 -8 32 272
use FILL  FILL_6__2318_
timestamp 1701859473
transform 1 0 6850 0 1 9110
box -12 -8 32 272
use FILL  FILL_6__2319_
timestamp 1701859473
transform -1 0 11170 0 1 4430
box -12 -8 32 272
use FILL  FILL_6__2320_
timestamp 1701859473
transform 1 0 5150 0 1 3910
box -12 -8 32 272
use FILL  FILL_6__2321_
timestamp 1701859473
transform 1 0 6570 0 1 3910
box -12 -8 32 272
use FILL  FILL_6__2322_
timestamp 1701859473
transform -1 0 7950 0 1 3910
box -12 -8 32 272
use FILL  FILL_6__2323_
timestamp 1701859473
transform 1 0 7990 0 -1 4430
box -12 -8 32 272
use FILL  FILL_6__2324_
timestamp 1701859473
transform -1 0 11210 0 -1 2870
box -12 -8 32 272
use FILL  FILL_6__2325_
timestamp 1701859473
transform -1 0 8190 0 1 3910
box -12 -8 32 272
use FILL  FILL_6__2326_
timestamp 1701859473
transform -1 0 3230 0 -1 4950
box -12 -8 32 272
use FILL  FILL_6__2327_
timestamp 1701859473
transform -1 0 3430 0 -1 4950
box -12 -8 32 272
use FILL  FILL_6__2328_
timestamp 1701859473
transform 1 0 3910 0 -1 5470
box -12 -8 32 272
use FILL  FILL_6__2329_
timestamp 1701859473
transform 1 0 3670 0 -1 5470
box -12 -8 32 272
use FILL  FILL_6__2330_
timestamp 1701859473
transform 1 0 3810 0 1 4950
box -12 -8 32 272
use FILL  FILL_6__2331_
timestamp 1701859473
transform 1 0 4890 0 1 3910
box -12 -8 32 272
use FILL  FILL_6__2332_
timestamp 1701859473
transform -1 0 4230 0 1 4950
box -12 -8 32 272
use FILL  FILL_6__2333_
timestamp 1701859473
transform -1 0 11190 0 -1 4430
box -12 -8 32 272
use FILL  FILL_6__2334_
timestamp 1701859473
transform 1 0 9070 0 -1 4430
box -12 -8 32 272
use FILL  FILL_6__2335_
timestamp 1701859473
transform 1 0 5250 0 -1 5470
box -12 -8 32 272
use FILL  FILL_6__2336_
timestamp 1701859473
transform -1 0 5110 0 1 5990
box -12 -8 32 272
use FILL  FILL_6__2337_
timestamp 1701859473
transform 1 0 4610 0 1 3390
box -12 -8 32 272
use FILL  FILL_6__2338_
timestamp 1701859473
transform 1 0 3210 0 1 3390
box -12 -8 32 272
use FILL  FILL_6__2339_
timestamp 1701859473
transform 1 0 4790 0 1 3390
box -12 -8 32 272
use FILL  FILL_6__2340_
timestamp 1701859473
transform 1 0 5030 0 1 3390
box -12 -8 32 272
use FILL  FILL_6__2341_
timestamp 1701859473
transform -1 0 610 0 1 5990
box -12 -8 32 272
use FILL  FILL_6__2342_
timestamp 1701859473
transform 1 0 2710 0 1 5470
box -12 -8 32 272
use FILL  FILL_6__2343_
timestamp 1701859473
transform -1 0 4650 0 1 6510
box -12 -8 32 272
use FILL  FILL_6__2344_
timestamp 1701859473
transform -1 0 4930 0 1 5470
box -12 -8 32 272
use FILL  FILL_6__2345_
timestamp 1701859473
transform -1 0 4730 0 1 5470
box -12 -8 32 272
use FILL  FILL_6__2346_
timestamp 1701859473
transform -1 0 4890 0 -1 5990
box -12 -8 32 272
use FILL  FILL_6__2347_
timestamp 1701859473
transform -1 0 5750 0 -1 5990
box -12 -8 32 272
use FILL  FILL_6__2348_
timestamp 1701859473
transform 1 0 5310 0 -1 6510
box -12 -8 32 272
use FILL  FILL_6__2349_
timestamp 1701859473
transform -1 0 5090 0 -1 6510
box -12 -8 32 272
use FILL  FILL_6__2350_
timestamp 1701859473
transform -1 0 4510 0 -1 6510
box -12 -8 32 272
use FILL  FILL_6__2351_
timestamp 1701859473
transform 1 0 5650 0 1 7030
box -12 -8 32 272
use FILL  FILL_6__2352_
timestamp 1701859473
transform -1 0 5870 0 1 7030
box -12 -8 32 272
use FILL  FILL_6__2353_
timestamp 1701859473
transform -1 0 810 0 1 7030
box -12 -8 32 272
use FILL  FILL_6__2354_
timestamp 1701859473
transform 1 0 5510 0 -1 5990
box -12 -8 32 272
use FILL  FILL_6__2355_
timestamp 1701859473
transform 1 0 5410 0 1 7030
box -12 -8 32 272
use FILL  FILL_6__2356_
timestamp 1701859473
transform -1 0 4910 0 -1 7550
box -12 -8 32 272
use FILL  FILL_6__2357_
timestamp 1701859473
transform 1 0 4770 0 1 8070
box -12 -8 32 272
use FILL  FILL_6__2358_
timestamp 1701859473
transform 1 0 5250 0 1 8070
box -12 -8 32 272
use FILL  FILL_6__2359_
timestamp 1701859473
transform -1 0 5570 0 -1 8590
box -12 -8 32 272
use FILL  FILL_6__2360_
timestamp 1701859473
transform -1 0 810 0 -1 6510
box -12 -8 32 272
use FILL  FILL_6__2361_
timestamp 1701859473
transform -1 0 5310 0 1 5990
box -12 -8 32 272
use FILL  FILL_6__2362_
timestamp 1701859473
transform 1 0 5310 0 1 6510
box -12 -8 32 272
use FILL  FILL_6__2363_
timestamp 1701859473
transform 1 0 5330 0 -1 7030
box -12 -8 32 272
use FILL  FILL_6__2364_
timestamp 1701859473
transform 1 0 5330 0 -1 8070
box -12 -8 32 272
use FILL  FILL_6__2365_
timestamp 1701859473
transform 1 0 5570 0 -1 8070
box -12 -8 32 272
use FILL  FILL_6__2366_
timestamp 1701859473
transform -1 0 5790 0 -1 8070
box -12 -8 32 272
use FILL  FILL_6__2367_
timestamp 1701859473
transform 1 0 2750 0 -1 7550
box -12 -8 32 272
use FILL  FILL_6__2368_
timestamp 1701859473
transform -1 0 5590 0 -1 7030
box -12 -8 32 272
use FILL  FILL_6__2369_
timestamp 1701859473
transform 1 0 5290 0 1 7550
box -12 -8 32 272
use FILL  FILL_6__2370_
timestamp 1701859473
transform -1 0 5330 0 -1 8590
box -12 -8 32 272
use FILL  FILL_6__2371_
timestamp 1701859473
transform 1 0 6010 0 -1 9110
box -12 -8 32 272
use FILL  FILL_6__2372_
timestamp 1701859473
transform 1 0 6170 0 1 9110
box -12 -8 32 272
use FILL  FILL_6__2373_
timestamp 1701859473
transform -1 0 6250 0 -1 9630
box -12 -8 32 272
use FILL  FILL_6__2374_
timestamp 1701859473
transform 1 0 130 0 -1 9110
box -12 -8 32 272
use FILL  FILL_6__2375_
timestamp 1701859473
transform -1 0 4270 0 1 5470
box -12 -8 32 272
use FILL  FILL_6__2376_
timestamp 1701859473
transform 1 0 4610 0 -1 5990
box -12 -8 32 272
use FILL  FILL_6__2377_
timestamp 1701859473
transform -1 0 4030 0 -1 6510
box -12 -8 32 272
use FILL  FILL_6__2378_
timestamp 1701859473
transform 1 0 3770 0 -1 6510
box -12 -8 32 272
use FILL  FILL_6__2379_
timestamp 1701859473
transform -1 0 5090 0 1 6510
box -12 -8 32 272
use FILL  FILL_6__2380_
timestamp 1701859473
transform -1 0 4870 0 -1 8590
box -12 -8 32 272
use FILL  FILL_6__2381_
timestamp 1701859473
transform 1 0 3930 0 -1 8590
box -12 -8 32 272
use FILL  FILL_6__2382_
timestamp 1701859473
transform -1 0 4630 0 -1 8590
box -12 -8 32 272
use FILL  FILL_6__2383_
timestamp 1701859473
transform -1 0 5710 0 1 8590
box -12 -8 32 272
use FILL  FILL_6__2384_
timestamp 1701859473
transform -1 0 5930 0 1 8590
box -12 -8 32 272
use FILL  FILL_6__2385_
timestamp 1701859473
transform 1 0 1310 0 -1 10150
box -12 -8 32 272
use FILL  FILL_6__2386_
timestamp 1701859473
transform 1 0 5570 0 -1 7550
box -12 -8 32 272
use FILL  FILL_6__2387_
timestamp 1701859473
transform 1 0 5550 0 -1 9110
box -12 -8 32 272
use FILL  FILL_6__2388_
timestamp 1701859473
transform -1 0 5350 0 -1 9110
box -12 -8 32 272
use FILL  FILL_6__2389_
timestamp 1701859473
transform -1 0 5130 0 -1 9630
box -12 -8 32 272
use FILL  FILL_6__2390_
timestamp 1701859473
transform 1 0 5190 0 1 9630
box -12 -8 32 272
use FILL  FILL_6__2391_
timestamp 1701859473
transform -1 0 5410 0 1 9630
box -12 -8 32 272
use FILL  FILL_6__2392_
timestamp 1701859473
transform 1 0 1510 0 -1 10150
box -12 -8 32 272
use FILL  FILL_6__2393_
timestamp 1701859473
transform -1 0 5370 0 -1 7550
box -12 -8 32 272
use FILL  FILL_6__2394_
timestamp 1701859473
transform 1 0 5450 0 1 8590
box -12 -8 32 272
use FILL  FILL_6__2395_
timestamp 1701859473
transform -1 0 5810 0 -1 9110
box -12 -8 32 272
use FILL  FILL_6__2396_
timestamp 1701859473
transform 1 0 5730 0 1 9110
box -12 -8 32 272
use FILL  FILL_6__2397_
timestamp 1701859473
transform 1 0 5970 0 1 9110
box -12 -8 32 272
use FILL  FILL_6__2398_
timestamp 1701859473
transform 1 0 5790 0 -1 9630
box -12 -8 32 272
use FILL  FILL_6__2399_
timestamp 1701859473
transform -1 0 3230 0 -1 5470
box -12 -8 32 272
use FILL  FILL_6__2400_
timestamp 1701859473
transform -1 0 3410 0 1 5990
box -12 -8 32 272
use FILL  FILL_6__2401_
timestamp 1701859473
transform 1 0 3330 0 -1 6510
box -12 -8 32 272
use FILL  FILL_6__2402_
timestamp 1701859473
transform -1 0 2270 0 -1 4430
box -12 -8 32 272
use FILL  FILL_6__2403_
timestamp 1701859473
transform -1 0 2670 0 1 4430
box -12 -8 32 272
use FILL  FILL_6__2404_
timestamp 1701859473
transform -1 0 2990 0 -1 5470
box -12 -8 32 272
use FILL  FILL_6__2405_
timestamp 1701859473
transform 1 0 2370 0 -1 2870
box -12 -8 32 272
use FILL  FILL_6__2406_
timestamp 1701859473
transform 1 0 3070 0 -1 3390
box -12 -8 32 272
use FILL  FILL_6__2407_
timestamp 1701859473
transform -1 0 3210 0 1 5470
box -12 -8 32 272
use FILL  FILL_6__2408_
timestamp 1701859473
transform 1 0 830 0 -1 2870
box -12 -8 32 272
use FILL  FILL_6__2409_
timestamp 1701859473
transform 1 0 850 0 -1 3910
box -12 -8 32 272
use FILL  FILL_6__2410_
timestamp 1701859473
transform 1 0 1250 0 1 4430
box -12 -8 32 272
use FILL  FILL_6__2411_
timestamp 1701859473
transform -1 0 810 0 -1 4950
box -12 -8 32 272
use FILL  FILL_6__2412_
timestamp 1701859473
transform 1 0 2490 0 -1 5990
box -12 -8 32 272
use FILL  FILL_6__2413_
timestamp 1701859473
transform 1 0 2950 0 1 5470
box -12 -8 32 272
use FILL  FILL_6__2414_
timestamp 1701859473
transform 1 0 4110 0 -1 5470
box -12 -8 32 272
use FILL  FILL_6__2415_
timestamp 1701859473
transform -1 0 4050 0 1 7030
box -12 -8 32 272
use FILL  FILL_6__2416_
timestamp 1701859473
transform 1 0 4010 0 1 4950
box -12 -8 32 272
use FILL  FILL_6__2417_
timestamp 1701859473
transform 1 0 4350 0 -1 5470
box -12 -8 32 272
use FILL  FILL_6__2418_
timestamp 1701859473
transform -1 0 1610 0 -1 4950
box -12 -8 32 272
use FILL  FILL_6__2419_
timestamp 1701859473
transform 1 0 2190 0 1 4430
box -12 -8 32 272
use FILL  FILL_6__2420_
timestamp 1701859473
transform 1 0 3850 0 1 5990
box -12 -8 32 272
use FILL  FILL_6__2421_
timestamp 1701859473
transform -1 0 3630 0 1 5990
box -12 -8 32 272
use FILL  FILL_6__2422_
timestamp 1701859473
transform -1 0 3510 0 -1 5990
box -12 -8 32 272
use FILL  FILL_6__2423_
timestamp 1701859473
transform -1 0 3730 0 -1 5990
box -12 -8 32 272
use FILL  FILL_6__2424_
timestamp 1701859473
transform 1 0 3270 0 -1 5990
box -12 -8 32 272
use FILL  FILL_6__2425_
timestamp 1701859473
transform 1 0 4410 0 1 5990
box -12 -8 32 272
use FILL  FILL_6__2426_
timestamp 1701859473
transform 1 0 4010 0 -1 7030
box -12 -8 32 272
use FILL  FILL_6__2427_
timestamp 1701859473
transform 1 0 4830 0 1 5990
box -12 -8 32 272
use FILL  FILL_6__2428_
timestamp 1701859473
transform 1 0 4590 0 1 5990
box -12 -8 32 272
use FILL  FILL_6__2429_
timestamp 1701859473
transform -1 0 4270 0 -1 6510
box -12 -8 32 272
use FILL  FILL_6__2430_
timestamp 1701859473
transform 1 0 4830 0 1 6510
box -12 -8 32 272
use FILL  FILL_6__2431_
timestamp 1701859473
transform -1 0 4930 0 -1 7030
box -12 -8 32 272
use FILL  FILL_6__2432_
timestamp 1701859473
transform 1 0 5150 0 -1 7030
box -12 -8 32 272
use FILL  FILL_6__2433_
timestamp 1701859473
transform -1 0 4410 0 -1 8070
box -12 -8 32 272
use FILL  FILL_6__2434_
timestamp 1701859473
transform 1 0 4890 0 1 7550
box -12 -8 32 272
use FILL  FILL_6__2435_
timestamp 1701859473
transform 1 0 4230 0 1 7030
box -12 -8 32 272
use FILL  FILL_6__2436_
timestamp 1701859473
transform -1 0 4670 0 -1 7550
box -12 -8 32 272
use FILL  FILL_6__2437_
timestamp 1701859473
transform -1 0 4650 0 -1 8070
box -12 -8 32 272
use FILL  FILL_6__2438_
timestamp 1701859473
transform -1 0 4890 0 -1 8070
box -12 -8 32 272
use FILL  FILL_6__2439_
timestamp 1701859473
transform -1 0 5130 0 -1 8070
box -12 -8 32 272
use FILL  FILL_6__2440_
timestamp 1701859473
transform 1 0 4670 0 1 10150
box -12 -8 32 272
use FILL  FILL_6__2441_
timestamp 1701859473
transform 1 0 3950 0 -1 7550
box -12 -8 32 272
use FILL  FILL_6__2442_
timestamp 1701859473
transform -1 0 4170 0 -1 8070
box -12 -8 32 272
use FILL  FILL_6__2443_
timestamp 1701859473
transform -1 0 3950 0 1 8070
box -12 -8 32 272
use FILL  FILL_6__2444_
timestamp 1701859473
transform 1 0 3690 0 1 8070
box -12 -8 32 272
use FILL  FILL_6__2445_
timestamp 1701859473
transform -1 0 4670 0 1 7550
box -12 -8 32 272
use FILL  FILL_6__2446_
timestamp 1701859473
transform 1 0 4590 0 1 8070
box -12 -8 32 272
use FILL  FILL_6__2447_
timestamp 1701859473
transform 1 0 4330 0 1 9110
box -12 -8 32 272
use FILL  FILL_6__2448_
timestamp 1701859473
transform 1 0 4990 0 1 9110
box -12 -8 32 272
use FILL  FILL_6__2449_
timestamp 1701859473
transform 1 0 5250 0 1 9110
box -12 -8 32 272
use FILL  FILL_6__2450_
timestamp 1701859473
transform 1 0 5490 0 1 9110
box -12 -8 32 272
use FILL  FILL_6__2451_
timestamp 1701859473
transform -1 0 5370 0 -1 9630
box -12 -8 32 272
use FILL  FILL_6__2452_
timestamp 1701859473
transform -1 0 5290 0 -1 10670
box -12 -8 32 272
use FILL  FILL_6__2453_
timestamp 1701859473
transform 1 0 3830 0 -1 10150
box -12 -8 32 272
use FILL  FILL_6__2454_
timestamp 1701859473
transform 1 0 3950 0 1 7550
box -12 -8 32 272
use FILL  FILL_6__2455_
timestamp 1701859473
transform 1 0 3910 0 -1 8070
box -12 -8 32 272
use FILL  FILL_6__2456_
timestamp 1701859473
transform -1 0 3690 0 -1 8070
box -12 -8 32 272
use FILL  FILL_6__2457_
timestamp 1701859473
transform 1 0 3450 0 1 8070
box -12 -8 32 272
use FILL  FILL_6__2458_
timestamp 1701859473
transform -1 0 4390 0 -1 8590
box -12 -8 32 272
use FILL  FILL_6__2459_
timestamp 1701859473
transform -1 0 4550 0 -1 11190
box -12 -8 32 272
use FILL  FILL_6__2460_
timestamp 1701859473
transform 1 0 4190 0 -1 10670
box -12 -8 32 272
use FILL  FILL_6__2461_
timestamp 1701859473
transform 1 0 4370 0 -1 9110
box -12 -8 32 272
use FILL  FILL_6__2462_
timestamp 1701859473
transform -1 0 4630 0 -1 9110
box -12 -8 32 272
use FILL  FILL_6__2463_
timestamp 1701859473
transform -1 0 4870 0 -1 9110
box -12 -8 32 272
use FILL  FILL_6__2464_
timestamp 1701859473
transform -1 0 5110 0 -1 9110
box -12 -8 32 272
use FILL  FILL_6__2465_
timestamp 1701859473
transform -1 0 4970 0 -1 11190
box -12 -8 32 272
use FILL  FILL_6__2466_
timestamp 1701859473
transform -1 0 4050 0 -1 10150
box -12 -8 32 272
use FILL  FILL_6__2467_
timestamp 1701859473
transform -1 0 4150 0 -1 9630
box -12 -8 32 272
use FILL  FILL_6__2468_
timestamp 1701859473
transform -1 0 4410 0 -1 9630
box -12 -8 32 272
use FILL  FILL_6__2469_
timestamp 1701859473
transform -1 0 4270 0 1 9630
box -12 -8 32 272
use FILL  FILL_6__2470_
timestamp 1701859473
transform -1 0 4510 0 1 9630
box -12 -8 32 272
use FILL  FILL_6__2471_
timestamp 1701859473
transform -1 0 5090 0 -1 10670
box -12 -8 32 272
use FILL  FILL_6__2472_
timestamp 1701859473
transform 1 0 4050 0 1 9630
box -12 -8 32 272
use FILL  FILL_6__2473_
timestamp 1701859473
transform 1 0 4610 0 -1 9630
box -12 -8 32 272
use FILL  FILL_6__2474_
timestamp 1701859473
transform -1 0 4890 0 -1 9630
box -12 -8 32 272
use FILL  FILL_6__2475_
timestamp 1701859473
transform 1 0 4730 0 1 9630
box -12 -8 32 272
use FILL  FILL_6__2476_
timestamp 1701859473
transform -1 0 4970 0 1 9630
box -12 -8 32 272
use FILL  FILL_6__2477_
timestamp 1701859473
transform 1 0 4910 0 1 10670
box -12 -8 32 272
use FILL  FILL_6__2478_
timestamp 1701859473
transform 1 0 3150 0 1 5990
box -12 -8 32 272
use FILL  FILL_6__2479_
timestamp 1701859473
transform -1 0 2710 0 1 5990
box -12 -8 32 272
use FILL  FILL_6__2480_
timestamp 1701859473
transform -1 0 2730 0 -1 5990
box -12 -8 32 272
use FILL  FILL_6__2481_
timestamp 1701859473
transform -1 0 2970 0 -1 5990
box -12 -8 32 272
use FILL  FILL_6__2482_
timestamp 1701859473
transform 1 0 1550 0 -1 5990
box -12 -8 32 272
use FILL  FILL_6__2483_
timestamp 1701859473
transform 1 0 2370 0 1 6510
box -12 -8 32 272
use FILL  FILL_6__2484_
timestamp 1701859473
transform -1 0 1990 0 1 6510
box -12 -8 32 272
use FILL  FILL_6__2485_
timestamp 1701859473
transform -1 0 2190 0 1 6510
box -12 -8 32 272
use FILL  FILL_6__2486_
timestamp 1701859473
transform 1 0 2390 0 -1 7030
box -12 -8 32 272
use FILL  FILL_6__2487_
timestamp 1701859473
transform 1 0 2150 0 -1 7030
box -12 -8 32 272
use FILL  FILL_6__2488_
timestamp 1701859473
transform -1 0 1950 0 -1 7030
box -12 -8 32 272
use FILL  FILL_6__2489_
timestamp 1701859473
transform 1 0 1450 0 -1 7030
box -12 -8 32 272
use FILL  FILL_6__2490_
timestamp 1701859473
transform -1 0 1050 0 1 5470
box -12 -8 32 272
use FILL  FILL_6__2491_
timestamp 1701859473
transform 1 0 1250 0 1 5470
box -12 -8 32 272
use FILL  FILL_6__2492_
timestamp 1701859473
transform -1 0 2110 0 -1 6510
box -12 -8 32 272
use FILL  FILL_6__2493_
timestamp 1701859473
transform 1 0 1990 0 1 5990
box -12 -8 32 272
use FILL  FILL_6__2494_
timestamp 1701859473
transform -1 0 1550 0 1 5990
box -12 -8 32 272
use FILL  FILL_6__2495_
timestamp 1701859473
transform 1 0 1290 0 1 5990
box -12 -8 32 272
use FILL  FILL_6__2496_
timestamp 1701859473
transform 1 0 1690 0 -1 7030
box -12 -8 32 272
use FILL  FILL_6__2497_
timestamp 1701859473
transform -1 0 1890 0 -1 7550
box -12 -8 32 272
use FILL  FILL_6__2498_
timestamp 1701859473
transform 1 0 830 0 1 8070
box -12 -8 32 272
use FILL  FILL_6__2499_
timestamp 1701859473
transform 1 0 2510 0 1 7550
box -12 -8 32 272
use FILL  FILL_6__2500_
timestamp 1701859473
transform 1 0 1930 0 1 7550
box -12 -8 32 272
use FILL  FILL_6__2501_
timestamp 1701859473
transform 1 0 1710 0 1 7550
box -12 -8 32 272
use FILL  FILL_6__2502_
timestamp 1701859473
transform -1 0 1250 0 1 7550
box -12 -8 32 272
use FILL  FILL_6__2503_
timestamp 1701859473
transform -1 0 1490 0 1 8070
box -12 -8 32 272
use FILL  FILL_6__2504_
timestamp 1701859473
transform -1 0 1910 0 1 8070
box -12 -8 32 272
use FILL  FILL_6__2505_
timestamp 1701859473
transform 1 0 1250 0 1 8070
box -12 -8 32 272
use FILL  FILL_6__2506_
timestamp 1701859473
transform -1 0 1770 0 -1 8070
box -12 -8 32 272
use FILL  FILL_6__2507_
timestamp 1701859473
transform 1 0 1510 0 -1 8070
box -12 -8 32 272
use FILL  FILL_6__2508_
timestamp 1701859473
transform 1 0 1030 0 1 8070
box -12 -8 32 272
use FILL  FILL_6__2509_
timestamp 1701859473
transform 1 0 590 0 -1 8590
box -12 -8 32 272
use FILL  FILL_6__2510_
timestamp 1701859473
transform -1 0 1530 0 1 9110
box -12 -8 32 272
use FILL  FILL_6__2511_
timestamp 1701859473
transform -1 0 1470 0 -1 9630
box -12 -8 32 272
use FILL  FILL_6__2512_
timestamp 1701859473
transform 1 0 1030 0 -1 9630
box -12 -8 32 272
use FILL  FILL_6__2513_
timestamp 1701859473
transform -1 0 1030 0 1 8590
box -12 -8 32 272
use FILL  FILL_6__2514_
timestamp 1701859473
transform 1 0 2110 0 -1 8590
box -12 -8 32 272
use FILL  FILL_6__2515_
timestamp 1701859473
transform 1 0 1230 0 -1 9110
box -12 -8 32 272
use FILL  FILL_6__2516_
timestamp 1701859473
transform -1 0 1070 0 1 9110
box -12 -8 32 272
use FILL  FILL_6__2517_
timestamp 1701859473
transform -1 0 830 0 1 9110
box -12 -8 32 272
use FILL  FILL_6__2518_
timestamp 1701859473
transform 1 0 1690 0 -1 9630
box -12 -8 32 272
use FILL  FILL_6__2519_
timestamp 1701859473
transform 1 0 1790 0 1 9630
box -12 -8 32 272
use FILL  FILL_6__2520_
timestamp 1701859473
transform -1 0 2630 0 -1 9110
box -12 -8 32 272
use FILL  FILL_6__2521_
timestamp 1701859473
transform 1 0 2370 0 -1 9110
box -12 -8 32 272
use FILL  FILL_6__2522_
timestamp 1701859473
transform -1 0 1990 0 1 9630
box -12 -8 32 272
use FILL  FILL_6__2523_
timestamp 1701859473
transform -1 0 2210 0 1 9630
box -12 -8 32 272
use FILL  FILL_6__2524_
timestamp 1701859473
transform -1 0 1950 0 -1 9110
box -12 -8 32 272
use FILL  FILL_6__2525_
timestamp 1701859473
transform 1 0 830 0 -1 8590
box -12 -8 32 272
use FILL  FILL_6__2526_
timestamp 1701859473
transform -1 0 1730 0 -1 8590
box -12 -8 32 272
use FILL  FILL_6__2527_
timestamp 1701859473
transform -1 0 1270 0 -1 8590
box -12 -8 32 272
use FILL  FILL_6__2528_
timestamp 1701859473
transform -1 0 1050 0 -1 8590
box -12 -8 32 272
use FILL  FILL_6__2529_
timestamp 1701859473
transform -1 0 1290 0 1 9110
box -12 -8 32 272
use FILL  FILL_6__2530_
timestamp 1701859473
transform -1 0 7550 0 -1 6510
box -12 -8 32 272
use FILL  FILL_6__2531_
timestamp 1701859473
transform 1 0 7970 0 1 7550
box -12 -8 32 272
use FILL  FILL_6__2532_
timestamp 1701859473
transform -1 0 9870 0 1 2870
box -12 -8 32 272
use FILL  FILL_6__2533_
timestamp 1701859473
transform -1 0 8950 0 1 4430
box -12 -8 32 272
use FILL  FILL_6__2534_
timestamp 1701859473
transform -1 0 9350 0 -1 5470
box -12 -8 32 272
use FILL  FILL_6__2535_
timestamp 1701859473
transform 1 0 130 0 -1 4950
box -12 -8 32 272
use FILL  FILL_6__2536_
timestamp 1701859473
transform 1 0 690 0 1 4950
box -12 -8 32 272
use FILL  FILL_6__2537_
timestamp 1701859473
transform 1 0 830 0 1 3390
box -12 -8 32 272
use FILL  FILL_6__2538_
timestamp 1701859473
transform -1 0 390 0 -1 3910
box -12 -8 32 272
use FILL  FILL_6__2539_
timestamp 1701859473
transform -1 0 150 0 1 4950
box -12 -8 32 272
use FILL  FILL_6__2540_
timestamp 1701859473
transform 1 0 3090 0 1 2350
box -12 -8 32 272
use FILL  FILL_6__2541_
timestamp 1701859473
transform -1 0 3350 0 1 2870
box -12 -8 32 272
use FILL  FILL_6__2542_
timestamp 1701859473
transform -1 0 2350 0 -1 6510
box -12 -8 32 272
use FILL  FILL_6__2543_
timestamp 1701859473
transform 1 0 910 0 1 4950
box -12 -8 32 272
use FILL  FILL_6__2544_
timestamp 1701859473
transform 1 0 1470 0 1 4430
box -12 -8 32 272
use FILL  FILL_6__2545_
timestamp 1701859473
transform 1 0 1330 0 -1 5470
box -12 -8 32 272
use FILL  FILL_6__2546_
timestamp 1701859473
transform -1 0 2070 0 -1 5470
box -12 -8 32 272
use FILL  FILL_6__2547_
timestamp 1701859473
transform 1 0 2010 0 -1 4430
box -12 -8 32 272
use FILL  FILL_6__2548_
timestamp 1701859473
transform 1 0 1130 0 1 4950
box -12 -8 32 272
use FILL  FILL_6__2549_
timestamp 1701859473
transform 1 0 1350 0 1 4950
box -12 -8 32 272
use FILL  FILL_6__2550_
timestamp 1701859473
transform -1 0 1830 0 -1 5470
box -12 -8 32 272
use FILL  FILL_6__2551_
timestamp 1701859473
transform 1 0 2610 0 -1 9630
box -12 -8 32 272
use FILL  FILL_6__2552_
timestamp 1701859473
transform 1 0 3450 0 -1 5470
box -12 -8 32 272
use FILL  FILL_6__2553_
timestamp 1701859473
transform -1 0 2830 0 -1 6510
box -12 -8 32 272
use FILL  FILL_6__2554_
timestamp 1701859473
transform -1 0 3290 0 1 6510
box -12 -8 32 272
use FILL  FILL_6__2555_
timestamp 1701859473
transform -1 0 3530 0 1 6510
box -12 -8 32 272
use FILL  FILL_6__2556_
timestamp 1701859473
transform -1 0 2850 0 1 6510
box -12 -8 32 272
use FILL  FILL_6__2557_
timestamp 1701859473
transform 1 0 2550 0 -1 6510
box -12 -8 32 272
use FILL  FILL_6__2558_
timestamp 1701859473
transform 1 0 3290 0 -1 7550
box -12 -8 32 272
use FILL  FILL_6__2559_
timestamp 1701859473
transform 1 0 3490 0 -1 7550
box -12 -8 32 272
use FILL  FILL_6__2560_
timestamp 1701859473
transform -1 0 3550 0 1 7030
box -12 -8 32 272
use FILL  FILL_6__2561_
timestamp 1701859473
transform -1 0 1570 0 1 4950
box -12 -8 32 272
use FILL  FILL_6__2562_
timestamp 1701859473
transform 1 0 3290 0 1 7030
box -12 -8 32 272
use FILL  FILL_6__2563_
timestamp 1701859473
transform 1 0 3850 0 1 5470
box -12 -8 32 272
use FILL  FILL_6__2564_
timestamp 1701859473
transform -1 0 3730 0 1 6510
box -12 -8 32 272
use FILL  FILL_6__2565_
timestamp 1701859473
transform 1 0 3790 0 1 7030
box -12 -8 32 272
use FILL  FILL_6__2566_
timestamp 1701859473
transform 1 0 3250 0 1 7550
box -12 -8 32 272
use FILL  FILL_6__2567_
timestamp 1701859473
transform 1 0 3210 0 -1 8070
box -12 -8 32 272
use FILL  FILL_6__2568_
timestamp 1701859473
transform -1 0 3030 0 -1 8590
box -12 -8 32 272
use FILL  FILL_6__2569_
timestamp 1701859473
transform 1 0 2790 0 -1 8590
box -12 -8 32 272
use FILL  FILL_6__2570_
timestamp 1701859473
transform 1 0 2970 0 -1 8070
box -12 -8 32 272
use FILL  FILL_6__2571_
timestamp 1701859473
transform -1 0 3930 0 -1 9630
box -12 -8 32 272
use FILL  FILL_6__2572_
timestamp 1701859473
transform -1 0 3950 0 -1 5990
box -12 -8 32 272
use FILL  FILL_6__2573_
timestamp 1701859473
transform -1 0 3810 0 -1 7030
box -12 -8 32 272
use FILL  FILL_6__2574_
timestamp 1701859473
transform 1 0 3530 0 -1 6510
box -12 -8 32 272
use FILL  FILL_6__2575_
timestamp 1701859473
transform 1 0 3430 0 -1 8070
box -12 -8 32 272
use FILL  FILL_6__2576_
timestamp 1701859473
transform -1 0 3470 0 -1 8590
box -12 -8 32 272
use FILL  FILL_6__2577_
timestamp 1701859473
transform 1 0 3350 0 1 9110
box -12 -8 32 272
use FILL  FILL_6__2578_
timestamp 1701859473
transform 1 0 3850 0 1 9110
box -12 -8 32 272
use FILL  FILL_6__2579_
timestamp 1701859473
transform -1 0 2830 0 -1 9630
box -12 -8 32 272
use FILL  FILL_6__2580_
timestamp 1701859473
transform -1 0 4190 0 -1 9110
box -12 -8 32 272
use FILL  FILL_6__2581_
timestamp 1701859473
transform -1 0 4110 0 1 9110
box -12 -8 32 272
use FILL  FILL_6__2582_
timestamp 1701859473
transform 1 0 3610 0 1 9110
box -12 -8 32 272
use FILL  FILL_6__2583_
timestamp 1701859473
transform 1 0 3110 0 1 9110
box -12 -8 32 272
use FILL  FILL_6__2584_
timestamp 1701859473
transform 1 0 2870 0 1 9110
box -12 -8 32 272
use FILL  FILL_6__2585_
timestamp 1701859473
transform 1 0 3970 0 -1 9110
box -12 -8 32 272
use FILL  FILL_6__2586_
timestamp 1701859473
transform 1 0 3130 0 1 9630
box -12 -8 32 272
use FILL  FILL_6__2587_
timestamp 1701859473
transform 1 0 3710 0 -1 9110
box -12 -8 32 272
use FILL  FILL_6__2588_
timestamp 1701859473
transform 1 0 3310 0 1 8590
box -12 -8 32 272
use FILL  FILL_6__2589_
timestamp 1701859473
transform 1 0 3150 0 -1 10150
box -12 -8 32 272
use FILL  FILL_6__2590_
timestamp 1701859473
transform 1 0 2890 0 -1 10150
box -12 -8 32 272
use FILL  FILL_6__2591_
timestamp 1701859473
transform -1 0 3650 0 -1 11190
box -12 -8 32 272
use FILL  FILL_6__2592_
timestamp 1701859473
transform -1 0 3710 0 -1 9630
box -12 -8 32 272
use FILL  FILL_6__2593_
timestamp 1701859473
transform -1 0 3230 0 -1 9630
box -12 -8 32 272
use FILL  FILL_6__2594_
timestamp 1701859473
transform -1 0 3390 0 -1 10150
box -12 -8 32 272
use FILL  FILL_6__2595_
timestamp 1701859473
transform 1 0 3110 0 -1 11190
box -12 -8 32 272
use FILL  FILL_6__2596_
timestamp 1701859473
transform 1 0 3390 0 -1 11190
box -12 -8 32 272
use FILL  FILL_6__2597_
timestamp 1701859473
transform 1 0 2850 0 -1 10670
box -12 -8 32 272
use FILL  FILL_6__2598_
timestamp 1701859473
transform -1 0 3590 0 1 9630
box -12 -8 32 272
use FILL  FILL_6__2599_
timestamp 1701859473
transform -1 0 3370 0 1 9630
box -12 -8 32 272
use FILL  FILL_6__2600_
timestamp 1701859473
transform -1 0 3090 0 1 10150
box -12 -8 32 272
use FILL  FILL_6__2601_
timestamp 1701859473
transform 1 0 3050 0 -1 10670
box -12 -8 32 272
use FILL  FILL_6__2602_
timestamp 1701859473
transform -1 0 3310 0 -1 10670
box -12 -8 32 272
use FILL  FILL_6__2603_
timestamp 1701859473
transform 1 0 3510 0 -1 10670
box -12 -8 32 272
use FILL  FILL_6__2604_
timestamp 1701859473
transform 1 0 3310 0 1 10150
box -12 -8 32 272
use FILL  FILL_6__2605_
timestamp 1701859473
transform 1 0 2430 0 1 10670
box -12 -8 32 272
use FILL  FILL_6__2606_
timestamp 1701859473
transform 1 0 2630 0 1 10670
box -12 -8 32 272
use FILL  FILL_6__2607_
timestamp 1701859473
transform -1 0 2870 0 1 10670
box -12 -8 32 272
use FILL  FILL_6__2608_
timestamp 1701859473
transform -1 0 3830 0 1 9630
box -12 -8 32 272
use FILL  FILL_6__2609_
timestamp 1701859473
transform -1 0 2450 0 1 9630
box -12 -8 32 272
use FILL  FILL_6__2610_
timestamp 1701859473
transform -1 0 2670 0 -1 10150
box -12 -8 32 272
use FILL  FILL_6__2611_
timestamp 1701859473
transform -1 0 2390 0 -1 10670
box -12 -8 32 272
use FILL  FILL_6__2612_
timestamp 1701859473
transform 1 0 2610 0 -1 10670
box -12 -8 32 272
use FILL  FILL_6__2613_
timestamp 1701859473
transform 1 0 1930 0 1 10670
box -12 -8 32 272
use FILL  FILL_6__2614_
timestamp 1701859473
transform 1 0 1930 0 -1 10670
box -12 -8 32 272
use FILL  FILL_6__2615_
timestamp 1701859473
transform -1 0 2450 0 -1 11190
box -12 -8 32 272
use FILL  FILL_6__2616_
timestamp 1701859473
transform -1 0 3470 0 -1 9630
box -12 -8 32 272
use FILL  FILL_6__2617_
timestamp 1701859473
transform 1 0 2370 0 -1 9630
box -12 -8 32 272
use FILL  FILL_6__2618_
timestamp 1701859473
transform -1 0 2650 0 1 10150
box -12 -8 32 272
use FILL  FILL_6__2619_
timestamp 1701859473
transform 1 0 2150 0 1 10670
box -12 -8 32 272
use FILL  FILL_6__2620_
timestamp 1701859473
transform 1 0 2190 0 -1 11190
box -12 -8 32 272
use FILL  FILL_6__2621_
timestamp 1701859473
transform -1 0 1470 0 1 5470
box -12 -8 32 272
use FILL  FILL_6__2622_
timestamp 1701859473
transform -1 0 1310 0 -1 5990
box -12 -8 32 272
use FILL  FILL_6__2623_
timestamp 1701859473
transform 1 0 2530 0 -1 5470
box -12 -8 32 272
use FILL  FILL_6__2624_
timestamp 1701859473
transform -1 0 2490 0 1 5470
box -12 -8 32 272
use FILL  FILL_6__2625_
timestamp 1701859473
transform 1 0 2290 0 -1 5470
box -12 -8 32 272
use FILL  FILL_6__2626_
timestamp 1701859473
transform -1 0 1030 0 -1 5470
box -12 -8 32 272
use FILL  FILL_6__2627_
timestamp 1701859473
transform -1 0 1550 0 1 3910
box -12 -8 32 272
use FILL  FILL_6__2628_
timestamp 1701859473
transform 1 0 1230 0 1 3910
box -12 -8 32 272
use FILL  FILL_6__2629_
timestamp 1701859473
transform -1 0 830 0 -1 5470
box -12 -8 32 272
use FILL  FILL_6__2630_
timestamp 1701859473
transform 1 0 810 0 -1 5990
box -12 -8 32 272
use FILL  FILL_6__2631_
timestamp 1701859473
transform -1 0 810 0 1 5990
box -12 -8 32 272
use FILL  FILL_6__2632_
timestamp 1701859473
transform 1 0 2190 0 1 10150
box -12 -8 32 272
use FILL  FILL_6__2633_
timestamp 1701859473
transform -1 0 2430 0 1 10150
box -12 -8 32 272
use FILL  FILL_6__2634_
timestamp 1701859473
transform 1 0 2390 0 -1 10150
box -12 -8 32 272
use FILL  FILL_6__2635_
timestamp 1701859473
transform 1 0 2170 0 -1 10150
box -12 -8 32 272
use FILL  FILL_6__2636_
timestamp 1701859473
transform -1 0 810 0 -1 10150
box -12 -8 32 272
use FILL  FILL_6__2637_
timestamp 1701859473
transform -1 0 610 0 1 6510
box -12 -8 32 272
use FILL  FILL_6__2638_
timestamp 1701859473
transform -1 0 390 0 1 6510
box -12 -8 32 272
use FILL  FILL_6__2639_
timestamp 1701859473
transform -1 0 370 0 -1 6510
box -12 -8 32 272
use FILL  FILL_6__2640_
timestamp 1701859473
transform -1 0 370 0 1 5990
box -12 -8 32 272
use FILL  FILL_6__2641_
timestamp 1701859473
transform 1 0 130 0 -1 7550
box -12 -8 32 272
use FILL  FILL_6__2642_
timestamp 1701859473
transform -1 0 470 0 1 4950
box -12 -8 32 272
use FILL  FILL_6__2643_
timestamp 1701859473
transform -1 0 2610 0 1 6510
box -12 -8 32 272
use FILL  FILL_6__2644_
timestamp 1701859473
transform 1 0 2650 0 -1 7030
box -12 -8 32 272
use FILL  FILL_6__2645_
timestamp 1701859473
transform 1 0 2830 0 1 7030
box -12 -8 32 272
use FILL  FILL_6__2646_
timestamp 1701859473
transform 1 0 2130 0 1 7030
box -12 -8 32 272
use FILL  FILL_6__2647_
timestamp 1701859473
transform 1 0 810 0 1 7550
box -12 -8 32 272
use FILL  FILL_6__2648_
timestamp 1701859473
transform 1 0 350 0 1 7550
box -12 -8 32 272
use FILL  FILL_6__2649_
timestamp 1701859473
transform 1 0 330 0 -1 7550
box -12 -8 32 272
use FILL  FILL_6__2650_
timestamp 1701859473
transform -1 0 810 0 -1 7550
box -12 -8 32 272
use FILL  FILL_6__2651_
timestamp 1701859473
transform 1 0 550 0 -1 7550
box -12 -8 32 272
use FILL  FILL_6__2652_
timestamp 1701859473
transform 1 0 550 0 1 7030
box -12 -8 32 272
use FILL  FILL_6__2653_
timestamp 1701859473
transform 1 0 130 0 1 7550
box -12 -8 32 272
use FILL  FILL_6__2654_
timestamp 1701859473
transform -1 0 610 0 1 7550
box -12 -8 32 272
use FILL  FILL_6__2655_
timestamp 1701859473
transform 1 0 1930 0 1 7030
box -12 -8 32 272
use FILL  FILL_6__2656_
timestamp 1701859473
transform 1 0 1570 0 -1 5470
box -12 -8 32 272
use FILL  FILL_6__2657_
timestamp 1701859473
transform -1 0 1770 0 1 5990
box -12 -8 32 272
use FILL  FILL_6__2658_
timestamp 1701859473
transform -1 0 2250 0 1 5470
box -12 -8 32 272
use FILL  FILL_6__2659_
timestamp 1701859473
transform 1 0 2010 0 -1 5990
box -12 -8 32 272
use FILL  FILL_6__2660_
timestamp 1701859473
transform -1 0 2010 0 1 5470
box -12 -8 32 272
use FILL  FILL_6__2661_
timestamp 1701859473
transform -1 0 1690 0 1 5470
box -12 -8 32 272
use FILL  FILL_6__2662_
timestamp 1701859473
transform 1 0 790 0 1 5470
box -12 -8 32 272
use FILL  FILL_6__2663_
timestamp 1701859473
transform -1 0 1070 0 -1 5990
box -12 -8 32 272
use FILL  FILL_6__2664_
timestamp 1701859473
transform 1 0 790 0 -1 7030
box -12 -8 32 272
use FILL  FILL_6__2665_
timestamp 1701859473
transform 1 0 1250 0 -1 7030
box -12 -8 32 272
use FILL  FILL_6__2666_
timestamp 1701859473
transform 1 0 1450 0 1 7030
box -12 -8 32 272
use FILL  FILL_6__2667_
timestamp 1701859473
transform 1 0 990 0 -1 7030
box -12 -8 32 272
use FILL  FILL_6__2668_
timestamp 1701859473
transform -1 0 2790 0 1 7550
box -12 -8 32 272
use FILL  FILL_6__2669_
timestamp 1701859473
transform 1 0 2730 0 -1 8070
box -12 -8 32 272
use FILL  FILL_6__2670_
timestamp 1701859473
transform 1 0 1990 0 -1 8070
box -12 -8 32 272
use FILL  FILL_6__2671_
timestamp 1701859473
transform -1 0 1490 0 1 7550
box -12 -8 32 272
use FILL  FILL_6__2672_
timestamp 1701859473
transform 1 0 1210 0 -1 7550
box -12 -8 32 272
use FILL  FILL_6__2673_
timestamp 1701859473
transform -1 0 1410 0 -1 7550
box -12 -8 32 272
use FILL  FILL_6__2674_
timestamp 1701859473
transform 1 0 1690 0 1 7030
box -12 -8 32 272
use FILL  FILL_6__2675_
timestamp 1701859473
transform 1 0 1630 0 -1 7550
box -12 -8 32 272
use FILL  FILL_6__2676_
timestamp 1701859473
transform -1 0 2070 0 -1 7550
box -12 -8 32 272
use FILL  FILL_6__2677_
timestamp 1701859473
transform 1 0 2470 0 -1 8070
box -12 -8 32 272
use FILL  FILL_6__2678_
timestamp 1701859473
transform -1 0 2250 0 -1 8070
box -12 -8 32 272
use FILL  FILL_6__2679_
timestamp 1701859473
transform -1 0 1690 0 1 8070
box -12 -8 32 272
use FILL  FILL_6__2680_
timestamp 1701859473
transform -1 0 370 0 -1 8590
box -12 -8 32 272
use FILL  FILL_6__2681_
timestamp 1701859473
transform 1 0 990 0 -1 7550
box -12 -8 32 272
use FILL  FILL_6__2682_
timestamp 1701859473
transform -1 0 370 0 -1 8070
box -12 -8 32 272
use FILL  FILL_6__2683_
timestamp 1701859473
transform -1 0 150 0 -1 9630
box -12 -8 32 272
use FILL  FILL_6__2684_
timestamp 1701859473
transform -1 0 150 0 1 10150
box -12 -8 32 272
use FILL  FILL_6__2685_
timestamp 1701859473
transform 1 0 1030 0 1 5990
box -12 -8 32 272
use FILL  FILL_6__2686_
timestamp 1701859473
transform 1 0 1010 0 1 7550
box -12 -8 32 272
use FILL  FILL_6__2687_
timestamp 1701859473
transform -1 0 1010 0 -1 10150
box -12 -8 32 272
use FILL  FILL_6__2688_
timestamp 1701859473
transform 1 0 130 0 -1 10150
box -12 -8 32 272
use FILL  FILL_6__2689_
timestamp 1701859473
transform 1 0 350 0 -1 9630
box -12 -8 32 272
use FILL  FILL_6__2690_
timestamp 1701859473
transform 1 0 350 0 1 9110
box -12 -8 32 272
use FILL  FILL_6__2691_
timestamp 1701859473
transform 1 0 2810 0 1 8590
box -12 -8 32 272
use FILL  FILL_6__2692_
timestamp 1701859473
transform 1 0 2570 0 1 8590
box -12 -8 32 272
use FILL  FILL_6__2693_
timestamp 1701859473
transform -1 0 1230 0 -1 9630
box -12 -8 32 272
use FILL  FILL_6__2694_
timestamp 1701859473
transform 1 0 810 0 -1 9630
box -12 -8 32 272
use FILL  FILL_6__2695_
timestamp 1701859473
transform 1 0 130 0 1 9630
box -12 -8 32 272
use FILL  FILL_6__2696_
timestamp 1701859473
transform -1 0 610 0 -1 10150
box -12 -8 32 272
use FILL  FILL_6__2697_
timestamp 1701859473
transform 1 0 350 0 -1 10150
box -12 -8 32 272
use FILL  FILL_6__2698_
timestamp 1701859473
transform 1 0 370 0 1 9630
box -12 -8 32 272
use FILL  FILL_6__2699_
timestamp 1701859473
transform 1 0 590 0 -1 9630
box -12 -8 32 272
use FILL  FILL_6__2700_
timestamp 1701859473
transform 1 0 610 0 1 9630
box -12 -8 32 272
use FILL  FILL_6__2701_
timestamp 1701859473
transform -1 0 830 0 -1 10670
box -12 -8 32 272
use FILL  FILL_6__2702_
timestamp 1701859473
transform 1 0 3550 0 1 8590
box -12 -8 32 272
use FILL  FILL_6__2703_
timestamp 1701859473
transform -1 0 3090 0 1 8590
box -12 -8 32 272
use FILL  FILL_6__2704_
timestamp 1701859473
transform -1 0 1570 0 1 9630
box -12 -8 32 272
use FILL  FILL_6__2705_
timestamp 1701859473
transform 1 0 1310 0 1 9630
box -12 -8 32 272
use FILL  FILL_6__2706_
timestamp 1701859473
transform 1 0 330 0 1 10150
box -12 -8 32 272
use FILL  FILL_6__2707_
timestamp 1701859473
transform -1 0 570 0 1 10150
box -12 -8 32 272
use FILL  FILL_6__2708_
timestamp 1701859473
transform 1 0 770 0 1 10150
box -12 -8 32 272
use FILL  FILL_6__2709_
timestamp 1701859473
transform -1 0 590 0 -1 10670
box -12 -8 32 272
use FILL  FILL_6__2710_
timestamp 1701859473
transform 1 0 1770 0 1 10150
box -12 -8 32 272
use FILL  FILL_6__2711_
timestamp 1701859473
transform 1 0 2310 0 1 8590
box -12 -8 32 272
use FILL  FILL_6__2712_
timestamp 1701859473
transform -1 0 2090 0 1 8590
box -12 -8 32 272
use FILL  FILL_6__2713_
timestamp 1701859473
transform -1 0 1950 0 -1 9630
box -12 -8 32 272
use FILL  FILL_6__2714_
timestamp 1701859473
transform 1 0 1710 0 -1 10150
box -12 -8 32 272
use FILL  FILL_6__2715_
timestamp 1701859473
transform 1 0 1030 0 1 10150
box -12 -8 32 272
use FILL  FILL_6__2716_
timestamp 1701859473
transform 1 0 1270 0 1 10150
box -12 -8 32 272
use FILL  FILL_6__2717_
timestamp 1701859473
transform 1 0 1530 0 1 10150
box -12 -8 32 272
use FILL  FILL_6__2718_
timestamp 1701859473
transform -1 0 10110 0 1 4950
box -12 -8 32 272
use FILL  FILL_6__2719_
timestamp 1701859473
transform -1 0 9870 0 1 4950
box -12 -8 32 272
use FILL  FILL_6__2720_
timestamp 1701859473
transform -1 0 4650 0 1 4950
box -12 -8 32 272
use FILL  FILL_6__2721_
timestamp 1701859473
transform -1 0 7410 0 -1 2350
box -12 -8 32 272
use FILL  FILL_6__2722_
timestamp 1701859473
transform 1 0 10050 0 -1 790
box -12 -8 32 272
use FILL  FILL_6__2723_
timestamp 1701859473
transform -1 0 7170 0 1 1830
box -12 -8 32 272
use FILL  FILL_6__2724_
timestamp 1701859473
transform -1 0 7170 0 -1 2350
box -12 -8 32 272
use FILL  FILL_6__2725_
timestamp 1701859473
transform 1 0 7030 0 1 3390
box -12 -8 32 272
use FILL  FILL_6__2726_
timestamp 1701859473
transform -1 0 7270 0 1 3390
box -12 -8 32 272
use FILL  FILL_6__2727_
timestamp 1701859473
transform -1 0 5490 0 1 3390
box -12 -8 32 272
use FILL  FILL_6__2728_
timestamp 1701859473
transform -1 0 5710 0 1 3390
box -12 -8 32 272
use FILL  FILL_6__2729_
timestamp 1701859473
transform -1 0 6810 0 -1 3910
box -12 -8 32 272
use FILL  FILL_6__2730_
timestamp 1701859473
transform 1 0 8310 0 -1 3910
box -12 -8 32 272
use FILL  FILL_6__2731_
timestamp 1701859473
transform 1 0 9330 0 1 1830
box -12 -8 32 272
use FILL  FILL_6__2732_
timestamp 1701859473
transform 1 0 7770 0 1 1830
box -12 -8 32 272
use FILL  FILL_6__2733_
timestamp 1701859473
transform 1 0 8650 0 1 2350
box -12 -8 32 272
use FILL  FILL_6__2734_
timestamp 1701859473
transform 1 0 7230 0 -1 5470
box -12 -8 32 272
use FILL  FILL_6__2735_
timestamp 1701859473
transform 1 0 7310 0 -1 2870
box -12 -8 32 272
use FILL  FILL_6__2736_
timestamp 1701859473
transform -1 0 7590 0 1 1310
box -12 -8 32 272
use FILL  FILL_6__2737_
timestamp 1701859473
transform 1 0 8650 0 1 1830
box -12 -8 32 272
use FILL  FILL_6__2738_
timestamp 1701859473
transform -1 0 8030 0 -1 2870
box -12 -8 32 272
use FILL  FILL_6__2739_
timestamp 1701859473
transform -1 0 7850 0 1 2870
box -12 -8 32 272
use FILL  FILL_6__2740_
timestamp 1701859473
transform -1 0 6630 0 -1 1830
box -12 -8 32 272
use FILL  FILL_6__2741_
timestamp 1701859473
transform 1 0 6830 0 -1 1830
box -12 -8 32 272
use FILL  FILL_6__2742_
timestamp 1701859473
transform -1 0 8270 0 -1 2870
box -12 -8 32 272
use FILL  FILL_6__2743_
timestamp 1701859473
transform -1 0 8290 0 1 2870
box -12 -8 32 272
use FILL  FILL_6__2744_
timestamp 1701859473
transform -1 0 7410 0 -1 270
box -12 -8 32 272
use FILL  FILL_6__2745_
timestamp 1701859473
transform -1 0 7370 0 1 1830
box -12 -8 32 272
use FILL  FILL_6__2746_
timestamp 1701859473
transform 1 0 8030 0 1 2870
box -12 -8 32 272
use FILL  FILL_6__2747_
timestamp 1701859473
transform -1 0 7830 0 -1 2350
box -12 -8 32 272
use FILL  FILL_6__2748_
timestamp 1701859473
transform 1 0 8010 0 -1 2350
box -12 -8 32 272
use FILL  FILL_6__2749_
timestamp 1701859473
transform 1 0 5970 0 1 1830
box -12 -8 32 272
use FILL  FILL_6__2750_
timestamp 1701859473
transform -1 0 6730 0 -1 1310
box -12 -8 32 272
use FILL  FILL_6__2751_
timestamp 1701859473
transform -1 0 6450 0 1 1830
box -12 -8 32 272
use FILL  FILL_6__2752_
timestamp 1701859473
transform -1 0 7810 0 1 2350
box -12 -8 32 272
use FILL  FILL_6__2753_
timestamp 1701859473
transform -1 0 7550 0 1 2350
box -12 -8 32 272
use FILL  FILL_6__2754_
timestamp 1701859473
transform 1 0 8890 0 -1 4950
box -12 -8 32 272
use FILL  FILL_6__2755_
timestamp 1701859473
transform 1 0 9790 0 1 790
box -12 -8 32 272
use FILL  FILL_6__2756_
timestamp 1701859473
transform -1 0 10030 0 1 790
box -12 -8 32 272
use FILL  FILL_6__2757_
timestamp 1701859473
transform 1 0 10730 0 -1 2870
box -12 -8 32 272
use FILL  FILL_6__2758_
timestamp 1701859473
transform -1 0 9230 0 -1 2870
box -12 -8 32 272
use FILL  FILL_6__2759_
timestamp 1701859473
transform 1 0 9150 0 1 4430
box -12 -8 32 272
use FILL  FILL_6__2760_
timestamp 1701859473
transform 1 0 10490 0 -1 790
box -12 -8 32 272
use FILL  FILL_6__2761_
timestamp 1701859473
transform 1 0 10250 0 -1 790
box -12 -8 32 272
use FILL  FILL_6__2762_
timestamp 1701859473
transform -1 0 10930 0 -1 1830
box -12 -8 32 272
use FILL  FILL_6__2763_
timestamp 1701859473
transform 1 0 6670 0 1 1830
box -12 -8 32 272
use FILL  FILL_6__2764_
timestamp 1701859473
transform -1 0 6930 0 1 1830
box -12 -8 32 272
use FILL  FILL_6__2765_
timestamp 1701859473
transform -1 0 10230 0 1 1830
box -12 -8 32 272
use FILL  FILL_6__2766_
timestamp 1701859473
transform -1 0 10050 0 -1 1830
box -12 -8 32 272
use FILL  FILL_6__2767_
timestamp 1701859473
transform -1 0 10470 0 -1 1830
box -12 -8 32 272
use FILL  FILL_6__2768_
timestamp 1701859473
transform -1 0 10450 0 1 1830
box -12 -8 32 272
use FILL  FILL_6__2769_
timestamp 1701859473
transform -1 0 10910 0 1 2350
box -12 -8 32 272
use FILL  FILL_6__2770_
timestamp 1701859473
transform -1 0 10690 0 -1 1830
box -12 -8 32 272
use FILL  FILL_6__2771_
timestamp 1701859473
transform 1 0 11110 0 1 2350
box -12 -8 32 272
use FILL  FILL_6__2772_
timestamp 1701859473
transform -1 0 10770 0 1 4950
box -12 -8 32 272
use FILL  FILL_6__2773_
timestamp 1701859473
transform 1 0 10510 0 -1 3910
box -12 -8 32 272
use FILL  FILL_6__2774_
timestamp 1701859473
transform -1 0 10810 0 -1 2350
box -12 -8 32 272
use FILL  FILL_6__2775_
timestamp 1701859473
transform -1 0 9170 0 -1 1310
box -12 -8 32 272
use FILL  FILL_6__2776_
timestamp 1701859473
transform 1 0 10710 0 -1 790
box -12 -8 32 272
use FILL  FILL_6__2777_
timestamp 1701859473
transform -1 0 8470 0 -1 270
box -12 -8 32 272
use FILL  FILL_6__2778_
timestamp 1701859473
transform 1 0 11010 0 1 270
box -12 -8 32 272
use FILL  FILL_6__2779_
timestamp 1701859473
transform 1 0 9090 0 -1 1830
box -12 -8 32 272
use FILL  FILL_6__2780_
timestamp 1701859473
transform -1 0 10110 0 1 1310
box -12 -8 32 272
use FILL  FILL_6__2781_
timestamp 1701859473
transform 1 0 10250 0 -1 1310
box -12 -8 32 272
use FILL  FILL_6__2782_
timestamp 1701859473
transform 1 0 8870 0 1 1830
box -12 -8 32 272
use FILL  FILL_6__2783_
timestamp 1701859473
transform 1 0 8430 0 -1 1310
box -12 -8 32 272
use FILL  FILL_6__2784_
timestamp 1701859473
transform 1 0 8670 0 -1 1310
box -12 -8 32 272
use FILL  FILL_6__2785_
timestamp 1701859473
transform 1 0 8890 0 -1 1830
box -12 -8 32 272
use FILL  FILL_6__2786_
timestamp 1701859473
transform -1 0 9370 0 -1 1310
box -12 -8 32 272
use FILL  FILL_6__2787_
timestamp 1701859473
transform -1 0 9570 0 -1 1830
box -12 -8 32 272
use FILL  FILL_6__2788_
timestamp 1701859473
transform 1 0 10250 0 -1 1830
box -12 -8 32 272
use FILL  FILL_6__2789_
timestamp 1701859473
transform 1 0 10330 0 1 1310
box -12 -8 32 272
use FILL  FILL_6__2790_
timestamp 1701859473
transform -1 0 10130 0 -1 2350
box -12 -8 32 272
use FILL  FILL_6__2791_
timestamp 1701859473
transform 1 0 9890 0 -1 2350
box -12 -8 32 272
use FILL  FILL_6__2792_
timestamp 1701859473
transform -1 0 10350 0 -1 2350
box -12 -8 32 272
use FILL  FILL_6__2793_
timestamp 1701859473
transform -1 0 10590 0 -1 2350
box -12 -8 32 272
use FILL  FILL_6__2794_
timestamp 1701859473
transform -1 0 11010 0 -1 2350
box -12 -8 32 272
use FILL  FILL_6__2795_
timestamp 1701859473
transform -1 0 10970 0 -1 2870
box -12 -8 32 272
use FILL  FILL_6__2796_
timestamp 1701859473
transform -1 0 10310 0 -1 2870
box -12 -8 32 272
use FILL  FILL_6__2797_
timestamp 1701859473
transform -1 0 9810 0 -1 1830
box -12 -8 32 272
use FILL  FILL_6__2798_
timestamp 1701859473
transform -1 0 10690 0 1 2350
box -12 -8 32 272
use FILL  FILL_6__2799_
timestamp 1701859473
transform 1 0 10470 0 -1 2870
box -12 -8 32 272
use FILL  FILL_6__2800_
timestamp 1701859473
transform -1 0 10490 0 -1 4430
box -12 -8 32 272
use FILL  FILL_6__2801_
timestamp 1701859473
transform -1 0 9450 0 -1 2870
box -12 -8 32 272
use FILL  FILL_6__2802_
timestamp 1701859473
transform -1 0 7310 0 -1 1830
box -12 -8 32 272
use FILL  FILL_6__2803_
timestamp 1701859473
transform 1 0 8510 0 -1 2870
box -12 -8 32 272
use FILL  FILL_6__2804_
timestamp 1701859473
transform -1 0 9570 0 -1 3390
box -12 -8 32 272
use FILL  FILL_6__2805_
timestamp 1701859473
transform -1 0 9870 0 -1 2870
box -12 -8 32 272
use FILL  FILL_6__2806_
timestamp 1701859473
transform 1 0 9630 0 -1 2870
box -12 -8 32 272
use FILL  FILL_6__2807_
timestamp 1701859473
transform 1 0 8970 0 -1 2350
box -12 -8 32 272
use FILL  FILL_6__2808_
timestamp 1701859473
transform 1 0 8730 0 -1 2350
box -12 -8 32 272
use FILL  FILL_6__2809_
timestamp 1701859473
transform 1 0 10450 0 1 2350
box -12 -8 32 272
use FILL  FILL_6__2810_
timestamp 1701859473
transform -1 0 10230 0 1 2350
box -12 -8 32 272
use FILL  FILL_6__2811_
timestamp 1701859473
transform 1 0 5010 0 -1 4430
box -12 -8 32 272
use FILL  FILL_6__2812_
timestamp 1701859473
transform -1 0 8970 0 1 4950
box -12 -8 32 272
use FILL  FILL_6__2813_
timestamp 1701859473
transform 1 0 9070 0 1 3390
box -12 -8 32 272
use FILL  FILL_6__2814_
timestamp 1701859473
transform -1 0 8890 0 -1 4430
box -12 -8 32 272
use FILL  FILL_6__2815_
timestamp 1701859473
transform -1 0 8670 0 1 3910
box -12 -8 32 272
use FILL  FILL_6__2816_
timestamp 1701859473
transform -1 0 8290 0 1 4950
box -12 -8 32 272
use FILL  FILL_6__2817_
timestamp 1701859473
transform 1 0 8730 0 1 4950
box -12 -8 32 272
use FILL  FILL_6__2818_
timestamp 1701859473
transform 1 0 8430 0 -1 4430
box -12 -8 32 272
use FILL  FILL_6__2819_
timestamp 1701859473
transform 1 0 8630 0 -1 4430
box -12 -8 32 272
use FILL  FILL_6__2820_
timestamp 1701859473
transform -1 0 9590 0 1 2350
box -12 -8 32 272
use FILL  FILL_6__2821_
timestamp 1701859473
transform 1 0 9110 0 1 2350
box -12 -8 32 272
use FILL  FILL_6__2822_
timestamp 1701859473
transform -1 0 9110 0 1 1830
box -12 -8 32 272
use FILL  FILL_6__2823_
timestamp 1701859473
transform -1 0 8890 0 1 2350
box -12 -8 32 272
use FILL  FILL_6__2824_
timestamp 1701859473
transform 1 0 10010 0 -1 3390
box -12 -8 32 272
use FILL  FILL_6__2825_
timestamp 1701859473
transform -1 0 10730 0 -1 3390
box -12 -8 32 272
use FILL  FILL_6__2826_
timestamp 1701859473
transform 1 0 9590 0 1 790
box -12 -8 32 272
use FILL  FILL_6__2827_
timestamp 1701859473
transform -1 0 9330 0 -1 1830
box -12 -8 32 272
use FILL  FILL_6__2828_
timestamp 1701859473
transform 1 0 7050 0 -1 1830
box -12 -8 32 272
use FILL  FILL_6__2829_
timestamp 1701859473
transform -1 0 10070 0 1 2870
box -12 -8 32 272
use FILL  FILL_6__2830_
timestamp 1701859473
transform 1 0 8370 0 -1 3390
box -12 -8 32 272
use FILL  FILL_6__2831_
timestamp 1701859473
transform 1 0 8410 0 1 3910
box -12 -8 32 272
use FILL  FILL_6__2832_
timestamp 1701859473
transform -1 0 9390 0 1 2350
box -12 -8 32 272
use FILL  FILL_6__2833_
timestamp 1701859473
transform -1 0 9330 0 -1 3390
box -12 -8 32 272
use FILL  FILL_6__2834_
timestamp 1701859473
transform -1 0 9090 0 -1 3390
box -12 -8 32 272
use FILL  FILL_6__2835_
timestamp 1701859473
transform -1 0 9390 0 1 790
box -12 -8 32 272
use FILL  FILL_6__2836_
timestamp 1701859473
transform 1 0 8970 0 1 1310
box -12 -8 32 272
use FILL  FILL_6__2837_
timestamp 1701859473
transform -1 0 9650 0 1 1310
box -12 -8 32 272
use FILL  FILL_6__2838_
timestamp 1701859473
transform -1 0 9770 0 1 3390
box -12 -8 32 272
use FILL  FILL_6__2839_
timestamp 1701859473
transform -1 0 9810 0 -1 3390
box -12 -8 32 272
use FILL  FILL_6__2840_
timestamp 1701859473
transform 1 0 9130 0 -1 270
box -12 -8 32 272
use FILL  FILL_6__2841_
timestamp 1701859473
transform -1 0 8930 0 -1 270
box -12 -8 32 272
use FILL  FILL_6__2842_
timestamp 1701859473
transform 1 0 9350 0 -1 270
box -12 -8 32 272
use FILL  FILL_6__2843_
timestamp 1701859473
transform 1 0 9590 0 -1 270
box -12 -8 32 272
use FILL  FILL_6__2844_
timestamp 1701859473
transform 1 0 9390 0 1 270
box -12 -8 32 272
use FILL  FILL_6__2845_
timestamp 1701859473
transform -1 0 10070 0 1 270
box -12 -8 32 272
use FILL  FILL_6__2846_
timestamp 1701859473
transform 1 0 9810 0 1 270
box -12 -8 32 272
use FILL  FILL_6__2847_
timestamp 1701859473
transform -1 0 11210 0 -1 10670
box -12 -8 32 272
use FILL  FILL_6__2848_
timestamp 1701859473
transform -1 0 10690 0 -1 1310
box -12 -8 32 272
use FILL  FILL_6__2849_
timestamp 1701859473
transform -1 0 11030 0 1 1310
box -12 -8 32 272
use FILL  FILL_6__2850_
timestamp 1701859473
transform -1 0 11170 0 -1 1830
box -12 -8 32 272
use FILL  FILL_6__2851_
timestamp 1701859473
transform 1 0 10770 0 -1 3910
box -12 -8 32 272
use FILL  FILL_6__2852_
timestamp 1701859473
transform -1 0 8970 0 1 270
box -12 -8 32 272
use FILL  FILL_6__2853_
timestamp 1701859473
transform -1 0 9190 0 1 270
box -12 -8 32 272
use FILL  FILL_6__2854_
timestamp 1701859473
transform 1 0 10690 0 1 790
box -12 -8 32 272
use FILL  FILL_6__2855_
timestamp 1701859473
transform -1 0 9890 0 1 1310
box -12 -8 32 272
use FILL  FILL_6__2856_
timestamp 1701859473
transform -1 0 10550 0 1 1310
box -12 -8 32 272
use FILL  FILL_6__2857_
timestamp 1701859473
transform -1 0 10790 0 1 1310
box -12 -8 32 272
use FILL  FILL_6__2858_
timestamp 1701859473
transform -1 0 11150 0 1 1830
box -12 -8 32 272
use FILL  FILL_6__2859_
timestamp 1701859473
transform 1 0 11010 0 -1 3910
box -12 -8 32 272
use FILL  FILL_6__2860_
timestamp 1701859473
transform 1 0 10930 0 -1 3390
box -12 -8 32 272
use FILL  FILL_6__2861_
timestamp 1701859473
transform 1 0 9810 0 -1 270
box -12 -8 32 272
use FILL  FILL_6__2862_
timestamp 1701859473
transform 1 0 8670 0 -1 270
box -12 -8 32 272
use FILL  FILL_6__2863_
timestamp 1701859473
transform -1 0 10310 0 1 270
box -12 -8 32 272
use FILL  FILL_6__2864_
timestamp 1701859473
transform 1 0 10550 0 1 270
box -12 -8 32 272
use FILL  FILL_6__2865_
timestamp 1701859473
transform -1 0 10790 0 1 270
box -12 -8 32 272
use FILL  FILL_6__2866_
timestamp 1701859473
transform -1 0 11170 0 -1 790
box -12 -8 32 272
use FILL  FILL_6__2867_
timestamp 1701859473
transform 1 0 11130 0 -1 3390
box -12 -8 32 272
use FILL  FILL_6__2868_
timestamp 1701859473
transform 1 0 11110 0 1 790
box -12 -8 32 272
use FILL  FILL_6__2869_
timestamp 1701859473
transform 1 0 10230 0 1 790
box -12 -8 32 272
use FILL  FILL_6__2870_
timestamp 1701859473
transform -1 0 10450 0 1 790
box -12 -8 32 272
use FILL  FILL_6__2871_
timestamp 1701859473
transform -1 0 10890 0 1 790
box -12 -8 32 272
use FILL  FILL_6__2872_
timestamp 1701859473
transform -1 0 11230 0 1 1310
box -12 -8 32 272
use FILL  FILL_6__2873_
timestamp 1701859473
transform -1 0 10010 0 1 3390
box -12 -8 32 272
use FILL  FILL_6__2874_
timestamp 1701859473
transform -1 0 10250 0 1 3390
box -12 -8 32 272
use FILL  FILL_6__2875_
timestamp 1701859473
transform -1 0 10830 0 -1 4950
box -12 -8 32 272
use FILL  FILL_6__2876_
timestamp 1701859473
transform -1 0 9790 0 1 1830
box -12 -8 32 272
use FILL  FILL_6__2877_
timestamp 1701859473
transform 1 0 9970 0 1 1830
box -12 -8 32 272
use FILL  FILL_6__2878_
timestamp 1701859473
transform 1 0 9790 0 -1 1310
box -12 -8 32 272
use FILL  FILL_6__2879_
timestamp 1701859473
transform -1 0 10030 0 -1 1310
box -12 -8 32 272
use FILL  FILL_6__2880_
timestamp 1701859473
transform 1 0 9530 0 1 1830
box -12 -8 32 272
use FILL  FILL_6__2881_
timestamp 1701859473
transform 1 0 10910 0 -1 790
box -12 -8 32 272
use FILL  FILL_6__2882_
timestamp 1701859473
transform -1 0 9590 0 -1 1310
box -12 -8 32 272
use FILL  FILL_6__2883_
timestamp 1701859473
transform -1 0 10490 0 -1 1310
box -12 -8 32 272
use FILL  FILL_6__2884_
timestamp 1701859473
transform 1 0 11130 0 -1 1310
box -12 -8 32 272
use FILL  FILL_6__2885_
timestamp 1701859473
transform -1 0 10910 0 -1 1310
box -12 -8 32 272
use FILL  FILL_6__2886_
timestamp 1701859473
transform 1 0 10670 0 1 1830
box -12 -8 32 272
use FILL  FILL_6__2887_
timestamp 1701859473
transform 1 0 10230 0 -1 4430
box -12 -8 32 272
use FILL  FILL_6__2888_
timestamp 1701859473
transform -1 0 4050 0 1 5470
box -12 -8 32 272
use FILL  FILL_6__2889_
timestamp 1701859473
transform 1 0 6170 0 1 2350
box -12 -8 32 272
use FILL  FILL_6__2890_
timestamp 1701859473
transform -1 0 8450 0 1 5990
box -12 -8 32 272
use FILL  FILL_6__2891_
timestamp 1701859473
transform -1 0 8250 0 1 5990
box -12 -8 32 272
use FILL  FILL_6__2892_
timestamp 1701859473
transform 1 0 7470 0 -1 5470
box -12 -8 32 272
use FILL  FILL_6__2893_
timestamp 1701859473
transform 1 0 7290 0 1 5470
box -12 -8 32 272
use FILL  FILL_6__2894_
timestamp 1701859473
transform 1 0 6570 0 -1 6510
box -12 -8 32 272
use FILL  FILL_6__2895_
timestamp 1701859473
transform 1 0 6710 0 1 6510
box -12 -8 32 272
use FILL  FILL_6__2896_
timestamp 1701859473
transform -1 0 7970 0 -1 5470
box -12 -8 32 272
use FILL  FILL_6__2897_
timestamp 1701859473
transform 1 0 7770 0 1 5470
box -12 -8 32 272
use FILL  FILL_6__2898_
timestamp 1701859473
transform 1 0 7290 0 -1 6510
box -12 -8 32 272
use FILL  FILL_6__2899_
timestamp 1701859473
transform 1 0 6810 0 -1 6510
box -12 -8 32 272
use FILL  FILL_6__2900_
timestamp 1701859473
transform -1 0 6350 0 -1 6510
box -12 -8 32 272
use FILL  FILL_6__2901_
timestamp 1701859473
transform 1 0 6090 0 -1 6510
box -12 -8 32 272
use FILL  FILL_6__2902_
timestamp 1701859473
transform -1 0 8010 0 1 5990
box -12 -8 32 272
use FILL  FILL_6__2903_
timestamp 1701859473
transform 1 0 7290 0 1 5990
box -12 -8 32 272
use FILL  FILL_6__2904_
timestamp 1701859473
transform 1 0 8410 0 -1 5470
box -12 -8 32 272
use FILL  FILL_6__2905_
timestamp 1701859473
transform 1 0 8430 0 1 5470
box -12 -8 32 272
use FILL  FILL_6__2906_
timestamp 1701859473
transform 1 0 8170 0 -1 5990
box -12 -8 32 272
use FILL  FILL_6__2907_
timestamp 1701859473
transform -1 0 7950 0 -1 5990
box -12 -8 32 272
use FILL  FILL_6__2908_
timestamp 1701859473
transform -1 0 8270 0 -1 4950
box -12 -8 32 272
use FILL  FILL_6__2909_
timestamp 1701859473
transform 1 0 3410 0 -1 4430
box -12 -8 32 272
use FILL  FILL_6__2910_
timestamp 1701859473
transform -1 0 6570 0 -1 4430
box -12 -8 32 272
use FILL  FILL_6__2911_
timestamp 1701859473
transform -1 0 6910 0 1 4430
box -12 -8 32 272
use FILL  FILL_6__2912_
timestamp 1701859473
transform 1 0 8690 0 -1 4950
box -12 -8 32 272
use FILL  FILL_6__2913_
timestamp 1701859473
transform -1 0 6870 0 -1 4950
box -12 -8 32 272
use FILL  FILL_6__2914_
timestamp 1701859473
transform 1 0 7130 0 -1 8070
box -12 -8 32 272
use FILL  FILL_6__2915_
timestamp 1701859473
transform 1 0 7250 0 -1 5990
box -12 -8 32 272
use FILL  FILL_6__2916_
timestamp 1701859473
transform 1 0 7010 0 -1 5990
box -12 -8 32 272
use FILL  FILL_6__2917_
timestamp 1701859473
transform -1 0 6390 0 -1 5990
box -12 -8 32 272
use FILL  FILL_6__2918_
timestamp 1701859473
transform 1 0 6310 0 1 5470
box -12 -8 32 272
use FILL  FILL_6__2919_
timestamp 1701859473
transform 1 0 6230 0 1 4950
box -12 -8 32 272
use FILL  FILL_6__2920_
timestamp 1701859473
transform 1 0 5990 0 1 4950
box -12 -8 32 272
use FILL  FILL_6__2921_
timestamp 1701859473
transform -1 0 7450 0 -1 3910
box -12 -8 32 272
use FILL  FILL_6__2922_
timestamp 1701859473
transform -1 0 7490 0 1 3910
box -12 -8 32 272
use FILL  FILL_6__2923_
timestamp 1701859473
transform -1 0 6810 0 -1 4430
box -12 -8 32 272
use FILL  FILL_6__2924_
timestamp 1701859473
transform 1 0 6430 0 1 4950
box -12 -8 32 272
use FILL  FILL_6__2925_
timestamp 1701859473
transform 1 0 7330 0 1 7550
box -12 -8 32 272
use FILL  FILL_6__2926_
timestamp 1701859473
transform -1 0 7570 0 1 4430
box -12 -8 32 272
use FILL  FILL_6__2927_
timestamp 1701859473
transform 1 0 7350 0 -1 4950
box -12 -8 32 272
use FILL  FILL_6__2928_
timestamp 1701859473
transform 1 0 7090 0 -1 4950
box -12 -8 32 272
use FILL  FILL_6__2929_
timestamp 1701859473
transform -1 0 6670 0 1 4950
box -12 -8 32 272
use FILL  FILL_6__2930_
timestamp 1701859473
transform 1 0 6210 0 1 1830
box -12 -8 32 272
use FILL  FILL_6__2931_
timestamp 1701859473
transform 1 0 7090 0 -1 2870
box -12 -8 32 272
use FILL  FILL_6__2932_
timestamp 1701859473
transform 1 0 5250 0 -1 4430
box -12 -8 32 272
use FILL  FILL_6__2933_
timestamp 1701859473
transform 1 0 5450 0 -1 4430
box -12 -8 32 272
use FILL  FILL_6__2934_
timestamp 1701859473
transform 1 0 5690 0 -1 4430
box -12 -8 32 272
use FILL  FILL_6__2935_
timestamp 1701859473
transform 1 0 6510 0 1 6510
box -12 -8 32 272
use FILL  FILL_6__2936_
timestamp 1701859473
transform 1 0 6390 0 -1 4950
box -12 -8 32 272
use FILL  FILL_6__2937_
timestamp 1701859473
transform 1 0 6610 0 -1 4950
box -12 -8 32 272
use FILL  FILL_6__2938_
timestamp 1701859473
transform 1 0 5090 0 1 4950
box -12 -8 32 272
use FILL  FILL_6__2939_
timestamp 1701859473
transform 1 0 4870 0 1 4950
box -12 -8 32 272
use FILL  FILL_6__2940_
timestamp 1701859473
transform -1 0 5930 0 -1 5470
box -12 -8 32 272
use FILL  FILL_6__2941_
timestamp 1701859473
transform 1 0 5690 0 -1 5470
box -12 -8 32 272
use FILL  FILL_6__2942_
timestamp 1701859473
transform -1 0 9390 0 1 4430
box -12 -8 32 272
use FILL  FILL_6__2943_
timestamp 1701859473
transform 1 0 6350 0 -1 4430
box -12 -8 32 272
use FILL  FILL_6__2944_
timestamp 1701859473
transform -1 0 6370 0 1 3910
box -12 -8 32 272
use FILL  FILL_6__2945_
timestamp 1701859473
transform -1 0 6450 0 1 4430
box -12 -8 32 272
use FILL  FILL_6__2946_
timestamp 1701859473
transform 1 0 6210 0 1 4430
box -12 -8 32 272
use FILL  FILL_6__2947_
timestamp 1701859473
transform -1 0 6610 0 -1 5990
box -12 -8 32 272
use FILL  FILL_6__2948_
timestamp 1701859473
transform 1 0 6150 0 -1 5990
box -12 -8 32 272
use FILL  FILL_6__2949_
timestamp 1701859473
transform -1 0 5970 0 -1 5990
box -12 -8 32 272
use FILL  FILL_6__2950_
timestamp 1701859473
transform 1 0 5830 0 1 5470
box -12 -8 32 272
use FILL  FILL_6__2951_
timestamp 1701859473
transform -1 0 6090 0 1 5470
box -12 -8 32 272
use FILL  FILL_6__2952_
timestamp 1701859473
transform -1 0 6170 0 -1 4950
box -12 -8 32 272
use FILL  FILL_6__2953_
timestamp 1701859473
transform -1 0 4450 0 1 4950
box -12 -8 32 272
use FILL  FILL_6__2954_
timestamp 1701859473
transform -1 0 6710 0 1 4430
box -12 -8 32 272
use FILL  FILL_6__2955_
timestamp 1701859473
transform -1 0 5990 0 1 4430
box -12 -8 32 272
use FILL  FILL_6__2956_
timestamp 1701859473
transform 1 0 5270 0 1 4430
box -12 -8 32 272
use FILL  FILL_6__2957_
timestamp 1701859473
transform 1 0 5210 0 -1 4950
box -12 -8 32 272
use FILL  FILL_6__2958_
timestamp 1701859473
transform -1 0 5530 0 1 4430
box -12 -8 32 272
use FILL  FILL_6__2959_
timestamp 1701859473
transform 1 0 7030 0 -1 5470
box -12 -8 32 272
use FILL  FILL_6__2960_
timestamp 1701859473
transform -1 0 6570 0 1 5470
box -12 -8 32 272
use FILL  FILL_6__2961_
timestamp 1701859473
transform 1 0 6330 0 -1 5470
box -12 -8 32 272
use FILL  FILL_6__2962_
timestamp 1701859473
transform -1 0 6590 0 -1 5470
box -12 -8 32 272
use FILL  FILL_6__2963_
timestamp 1701859473
transform -1 0 6830 0 -1 5470
box -12 -8 32 272
use FILL  FILL_6__2964_
timestamp 1701859473
transform -1 0 5470 0 -1 4950
box -12 -8 32 272
use FILL  FILL_6__2965_
timestamp 1701859473
transform 1 0 4970 0 -1 4950
box -12 -8 32 272
use FILL  FILL_6__2966_
timestamp 1701859473
transform -1 0 6430 0 1 2350
box -12 -8 32 272
use FILL  FILL_6__2967_
timestamp 1701859473
transform 1 0 7690 0 1 3910
box -12 -8 32 272
use FILL  FILL_6__2968_
timestamp 1701859473
transform -1 0 7010 0 -1 3910
box -12 -8 32 272
use FILL  FILL_6__2969_
timestamp 1701859473
transform -1 0 7230 0 -1 3910
box -12 -8 32 272
use FILL  FILL_6__2970_
timestamp 1701859473
transform -1 0 7270 0 1 3910
box -12 -8 32 272
use FILL  FILL_6__2971_
timestamp 1701859473
transform -1 0 6790 0 1 3910
box -12 -8 32 272
use FILL  FILL_6__2972_
timestamp 1701859473
transform 1 0 7010 0 1 3910
box -12 -8 32 272
use FILL  FILL_6__2973_
timestamp 1701859473
transform -1 0 7130 0 1 4430
box -12 -8 32 272
use FILL  FILL_6__2974_
timestamp 1701859473
transform 1 0 7030 0 -1 4430
box -12 -8 32 272
use FILL  FILL_6__2975_
timestamp 1701859473
transform -1 0 7790 0 -1 4430
box -12 -8 32 272
use FILL  FILL_6__2976_
timestamp 1701859473
transform -1 0 7550 0 -1 4430
box -12 -8 32 272
use FILL  FILL_6__2977_
timestamp 1701859473
transform 1 0 7270 0 -1 4430
box -12 -8 32 272
use FILL  FILL_6__2978_
timestamp 1701859473
transform 1 0 7330 0 1 4430
box -12 -8 32 272
use FILL  FILL_6__2979_
timestamp 1701859473
transform -1 0 3670 0 -1 4950
box -12 -8 32 272
use FILL  FILL_6__2980_
timestamp 1701859473
transform -1 0 3050 0 1 7550
box -12 -8 32 272
use FILL  FILL_6__2981_
timestamp 1701859473
transform 1 0 3570 0 1 4950
box -12 -8 32 272
use FILL  FILL_6__2982_
timestamp 1701859473
transform 1 0 9630 0 1 6510
box -12 -8 32 272
use FILL  FILL_6__2983_
timestamp 1701859473
transform 1 0 1950 0 1 4430
box -12 -8 32 272
use FILL  FILL_6__2984_
timestamp 1701859473
transform -1 0 3570 0 -1 3910
box -12 -8 32 272
use FILL  FILL_6__2985_
timestamp 1701859473
transform 1 0 3730 0 1 4430
box -12 -8 32 272
use FILL  FILL_6__2986_
timestamp 1701859473
transform -1 0 5930 0 -1 4430
box -12 -8 32 272
use FILL  FILL_6__2987_
timestamp 1701859473
transform -1 0 5750 0 1 4430
box -12 -8 32 272
use FILL  FILL_6__2988_
timestamp 1701859473
transform 1 0 9410 0 1 6510
box -12 -8 32 272
use FILL  FILL_6__2989_
timestamp 1701859473
transform 1 0 6030 0 1 6510
box -12 -8 32 272
use FILL  FILL_6__2990_
timestamp 1701859473
transform -1 0 6290 0 1 6510
box -12 -8 32 272
use FILL  FILL_6__2991_
timestamp 1701859473
transform 1 0 7190 0 1 6510
box -12 -8 32 272
use FILL  FILL_6__2992_
timestamp 1701859473
transform 1 0 9710 0 1 7030
box -12 -8 32 272
use FILL  FILL_6__2993_
timestamp 1701859473
transform 1 0 9910 0 1 7030
box -12 -8 32 272
use FILL  FILL_6__2994_
timestamp 1701859473
transform -1 0 10830 0 -1 7550
box -12 -8 32 272
use FILL  FILL_6__2995_
timestamp 1701859473
transform -1 0 7630 0 -1 7550
box -12 -8 32 272
use FILL  FILL_6__2996_
timestamp 1701859473
transform 1 0 7530 0 1 7550
box -12 -8 32 272
use FILL  FILL_6__2997_
timestamp 1701859473
transform -1 0 7410 0 -1 7550
box -12 -8 32 272
use FILL  FILL_6__2998_
timestamp 1701859473
transform -1 0 6470 0 -1 7550
box -12 -8 32 272
use FILL  FILL_6__2999_
timestamp 1701859473
transform 1 0 6190 0 1 7550
box -12 -8 32 272
use FILL  FILL_6__3000_
timestamp 1701859473
transform -1 0 6030 0 -1 7550
box -12 -8 32 272
use FILL  FILL_6__3001_
timestamp 1701859473
transform -1 0 5810 0 -1 7550
box -12 -8 32 272
use FILL  FILL_6__3002_
timestamp 1701859473
transform -1 0 6230 0 -1 7550
box -12 -8 32 272
use FILL  FILL_6__3003_
timestamp 1701859473
transform -1 0 6410 0 1 7550
box -12 -8 32 272
use FILL  FILL_6__3004_
timestamp 1701859473
transform 1 0 8210 0 1 7550
box -12 -8 32 272
use FILL  FILL_6__3005_
timestamp 1701859473
transform 1 0 11030 0 -1 7550
box -12 -8 32 272
use FILL  FILL_6__3006_
timestamp 1701859473
transform -1 0 10510 0 1 7550
box -12 -8 32 272
use FILL  FILL_6__3007_
timestamp 1701859473
transform 1 0 7030 0 1 7030
box -12 -8 32 272
use FILL  FILL_6__3008_
timestamp 1701859473
transform -1 0 6590 0 1 7030
box -12 -8 32 272
use FILL  FILL_6__3009_
timestamp 1701859473
transform -1 0 5990 0 -1 7030
box -12 -8 32 272
use FILL  FILL_6__3010_
timestamp 1701859473
transform 1 0 6210 0 -1 7030
box -12 -8 32 272
use FILL  FILL_6__3011_
timestamp 1701859473
transform 1 0 6790 0 1 7030
box -12 -8 32 272
use FILL  FILL_6__3012_
timestamp 1701859473
transform -1 0 7910 0 -1 7030
box -12 -8 32 272
use FILL  FILL_6__3013_
timestamp 1701859473
transform 1 0 8350 0 -1 7030
box -12 -8 32 272
use FILL  FILL_6__3014_
timestamp 1701859473
transform 1 0 10710 0 1 7550
box -12 -8 32 272
use FILL  FILL_6__3015_
timestamp 1701859473
transform -1 0 6430 0 -1 7030
box -12 -8 32 272
use FILL  FILL_6__3016_
timestamp 1701859473
transform -1 0 7310 0 1 7030
box -12 -8 32 272
use FILL  FILL_6__3017_
timestamp 1701859473
transform 1 0 6650 0 -1 7030
box -12 -8 32 272
use FILL  FILL_6__3018_
timestamp 1701859473
transform -1 0 6950 0 -1 7030
box -12 -8 32 272
use FILL  FILL_6__3019_
timestamp 1701859473
transform -1 0 7190 0 -1 7030
box -12 -8 32 272
use FILL  FILL_6__3020_
timestamp 1701859473
transform 1 0 8350 0 1 7030
box -12 -8 32 272
use FILL  FILL_6__3021_
timestamp 1701859473
transform -1 0 9410 0 -1 8070
box -12 -8 32 272
use FILL  FILL_6__3022_
timestamp 1701859473
transform 1 0 9590 0 -1 8070
box -12 -8 32 272
use FILL  FILL_6__3023_
timestamp 1701859473
transform -1 0 5810 0 1 6510
box -12 -8 32 272
use FILL  FILL_6__3024_
timestamp 1701859473
transform 1 0 5550 0 1 6510
box -12 -8 32 272
use FILL  FILL_6__3025_
timestamp 1701859473
transform -1 0 5570 0 -1 6510
box -12 -8 32 272
use FILL  FILL_6__3026_
timestamp 1701859473
transform 1 0 10990 0 -1 5990
box -12 -8 32 272
use FILL  FILL_6__3027_
timestamp 1701859473
transform -1 0 11230 0 -1 5990
box -12 -8 32 272
use FILL  FILL_6__3028_
timestamp 1701859473
transform -1 0 9850 0 -1 8070
box -12 -8 32 272
use FILL  FILL_6__3029_
timestamp 1701859473
transform -1 0 7170 0 -1 7550
box -12 -8 32 272
use FILL  FILL_6__3030_
timestamp 1701859473
transform -1 0 8150 0 -1 7030
box -12 -8 32 272
use FILL  FILL_6__3031_
timestamp 1701859473
transform 1 0 8130 0 1 7030
box -12 -8 32 272
use FILL  FILL_6__3032_
timestamp 1701859473
transform 1 0 7750 0 1 7550
box -12 -8 32 272
use FILL  FILL_6__3033_
timestamp 1701859473
transform -1 0 6830 0 1 8070
box -12 -8 32 272
use FILL  FILL_6__3034_
timestamp 1701859473
transform -1 0 7810 0 -1 8070
box -12 -8 32 272
use FILL  FILL_6__3035_
timestamp 1701859473
transform 1 0 7550 0 -1 8070
box -12 -8 32 272
use FILL  FILL_6__3036_
timestamp 1701859473
transform -1 0 7030 0 1 8070
box -12 -8 32 272
use FILL  FILL_6__3037_
timestamp 1701859473
transform -1 0 6590 0 1 8070
box -12 -8 32 272
use FILL  FILL_6__3038_
timestamp 1701859473
transform -1 0 7210 0 1 8070
box -12 -8 32 272
use FILL  FILL_6__3039_
timestamp 1701859473
transform 1 0 7430 0 1 8070
box -12 -8 32 272
use FILL  FILL_6__3040_
timestamp 1701859473
transform 1 0 9770 0 1 7550
box -12 -8 32 272
use FILL  FILL_6__3041_
timestamp 1701859473
transform -1 0 9630 0 -1 6510
box -12 -8 32 272
use FILL  FILL_6__3042_
timestamp 1701859473
transform 1 0 7330 0 -1 8070
box -12 -8 32 272
use FILL  FILL_6__3043_
timestamp 1701859473
transform -1 0 6650 0 1 7550
box -12 -8 32 272
use FILL  FILL_6__3044_
timestamp 1701859473
transform -1 0 6690 0 -1 7550
box -12 -8 32 272
use FILL  FILL_6__3045_
timestamp 1701859473
transform 1 0 6910 0 -1 7550
box -12 -8 32 272
use FILL  FILL_6__3046_
timestamp 1701859473
transform -1 0 7870 0 1 6510
box -12 -8 32 272
use FILL  FILL_6__3047_
timestamp 1701859473
transform 1 0 9210 0 1 6510
box -12 -8 32 272
use FILL  FILL_6__3048_
timestamp 1701859473
transform 1 0 9830 0 -1 6510
box -12 -8 32 272
use FILL  FILL_6__3049_
timestamp 1701859473
transform -1 0 6910 0 1 7550
box -12 -8 32 272
use FILL  FILL_6__3050_
timestamp 1701859473
transform -1 0 7130 0 1 7550
box -12 -8 32 272
use FILL  FILL_6__3051_
timestamp 1701859473
transform -1 0 7870 0 1 7030
box -12 -8 32 272
use FILL  FILL_6__3052_
timestamp 1701859473
transform 1 0 7570 0 1 7030
box -12 -8 32 272
use FILL  FILL_6__3053_
timestamp 1701859473
transform 1 0 7410 0 -1 7030
box -12 -8 32 272
use FILL  FILL_6__3054_
timestamp 1701859473
transform -1 0 7670 0 -1 7030
box -12 -8 32 272
use FILL  FILL_6__3055_
timestamp 1701859473
transform 1 0 8090 0 1 6510
box -12 -8 32 272
use FILL  FILL_6__3056_
timestamp 1701859473
transform -1 0 9610 0 1 5470
box -12 -8 32 272
use FILL  FILL_6__3057_
timestamp 1701859473
transform -1 0 9370 0 1 5470
box -12 -8 32 272
use FILL  FILL_6__3058_
timestamp 1701859473
transform 1 0 8790 0 -1 7550
box -12 -8 32 272
use FILL  FILL_6__3059_
timestamp 1701859473
transform -1 0 8670 0 -1 5990
box -12 -8 32 272
use FILL  FILL_6__3060_
timestamp 1701859473
transform 1 0 9850 0 1 6510
box -12 -8 32 272
use FILL  FILL_6__3061_
timestamp 1701859473
transform 1 0 10090 0 1 6510
box -12 -8 32 272
use FILL  FILL_6__3062_
timestamp 1701859473
transform -1 0 9710 0 -1 7550
box -12 -8 32 272
use FILL  FILL_6__3063_
timestamp 1701859473
transform 1 0 9450 0 -1 7550
box -12 -8 32 272
use FILL  FILL_6__3064_
timestamp 1701859473
transform -1 0 10410 0 -1 7030
box -12 -8 32 272
use FILL  FILL_6__3065_
timestamp 1701859473
transform -1 0 10650 0 -1 7030
box -12 -8 32 272
use FILL  FILL_6__3066_
timestamp 1701859473
transform -1 0 8570 0 -1 7550
box -12 -8 32 272
use FILL  FILL_6__3067_
timestamp 1701859473
transform 1 0 8310 0 -1 7550
box -12 -8 32 272
use FILL  FILL_6__3068_
timestamp 1701859473
transform 1 0 10270 0 -1 5990
box -12 -8 32 272
use FILL  FILL_6__3069_
timestamp 1701859473
transform 1 0 10510 0 -1 5990
box -12 -8 32 272
use FILL  FILL_6__3070_
timestamp 1701859473
transform 1 0 8970 0 -1 7550
box -12 -8 32 272
use FILL  FILL_6__3071_
timestamp 1701859473
transform -1 0 9230 0 -1 7550
box -12 -8 32 272
use FILL  FILL_6__3072_
timestamp 1701859473
transform -1 0 9850 0 1 5990
box -12 -8 32 272
use FILL  FILL_6__3073_
timestamp 1701859473
transform -1 0 10070 0 1 5990
box -12 -8 32 272
use FILL  FILL_6__3074_
timestamp 1701859473
transform 1 0 8890 0 1 5990
box -12 -8 32 272
use FILL  FILL_6__3075_
timestamp 1701859473
transform 1 0 8890 0 -1 5990
box -12 -8 32 272
use FILL  FILL_6__3076_
timestamp 1701859473
transform 1 0 10790 0 1 6510
box -12 -8 32 272
use FILL  FILL_6__3077_
timestamp 1701859473
transform 1 0 10990 0 1 6510
box -12 -8 32 272
use FILL  FILL_6__3078_
timestamp 1701859473
transform -1 0 8790 0 -1 7030
box -12 -8 32 272
use FILL  FILL_6__3079_
timestamp 1701859473
transform -1 0 8570 0 -1 7030
box -12 -8 32 272
use FILL  FILL_6__3080_
timestamp 1701859473
transform 1 0 11050 0 -1 8590
box -12 -8 32 272
use FILL  FILL_6__3081_
timestamp 1701859473
transform -1 0 11050 0 -1 270
box -12 -8 32 272
use FILL  FILL_6__3082_
timestamp 1701859473
transform 1 0 10150 0 -1 8590
box -12 -8 32 272
use FILL  FILL_6__3083_
timestamp 1701859473
transform -1 0 9930 0 -1 8590
box -12 -8 32 272
use FILL  FILL_6__3084_
timestamp 1701859473
transform -1 0 9110 0 1 7550
box -12 -8 32 272
use FILL  FILL_6__3085_
timestamp 1701859473
transform 1 0 9010 0 1 7030
box -12 -8 32 272
use FILL  FILL_6__3086_
timestamp 1701859473
transform -1 0 10770 0 1 5990
box -12 -8 32 272
use FILL  FILL_6__3087_
timestamp 1701859473
transform 1 0 10970 0 1 5990
box -12 -8 32 272
use FILL  FILL_6__3088_
timestamp 1701859473
transform 1 0 8330 0 1 8070
box -12 -8 32 272
use FILL  FILL_6__3089_
timestamp 1701859473
transform -1 0 8110 0 1 8070
box -12 -8 32 272
use FILL  FILL_6__3090_
timestamp 1701859473
transform -1 0 11210 0 1 4950
box -12 -8 32 272
use FILL  FILL_6__3091_
timestamp 1701859473
transform 1 0 10950 0 1 4950
box -12 -8 32 272
use FILL  FILL_6__3092_
timestamp 1701859473
transform 1 0 8870 0 -1 5470
box -12 -8 32 272
use FILL  FILL_6__3093_
timestamp 1701859473
transform -1 0 9110 0 -1 5470
box -12 -8 32 272
use FILL  FILL_6__3094_
timestamp 1701859473
transform -1 0 10310 0 -1 5470
box -12 -8 32 272
use FILL  FILL_6__3095_
timestamp 1701859473
transform 1 0 10250 0 1 5470
box -12 -8 32 272
use FILL  FILL_6__3096_
timestamp 1701859473
transform 1 0 8990 0 1 6510
box -12 -8 32 272
use FILL  FILL_6__3097_
timestamp 1701859473
transform -1 0 8770 0 1 6510
box -12 -8 32 272
use FILL  FILL_6__3098_
timestamp 1701859473
transform -1 0 10470 0 1 8070
box -12 -8 32 272
use FILL  FILL_6__3099_
timestamp 1701859473
transform -1 0 11230 0 -1 8070
box -12 -8 32 272
use FILL  FILL_6__3100_
timestamp 1701859473
transform 1 0 10230 0 1 8070
box -12 -8 32 272
use FILL  FILL_6__3101_
timestamp 1701859473
transform 1 0 10370 0 -1 8590
box -12 -8 32 272
use FILL  FILL_6__3102_
timestamp 1701859473
transform 1 0 8450 0 -1 8070
box -12 -8 32 272
use FILL  FILL_6__3103_
timestamp 1701859473
transform -1 0 8430 0 1 7550
box -12 -8 32 272
use FILL  FILL_6__3104_
timestamp 1701859473
transform -1 0 11230 0 1 6510
box -12 -8 32 272
use FILL  FILL_6__3105_
timestamp 1701859473
transform -1 0 11030 0 -1 4950
box -12 -8 32 272
use FILL  FILL_6__3106_
timestamp 1701859473
transform 1 0 9450 0 -1 8590
box -12 -8 32 272
use FILL  FILL_6__3107_
timestamp 1701859473
transform -1 0 9690 0 -1 8590
box -12 -8 32 272
use FILL  FILL_6__3108_
timestamp 1701859473
transform 1 0 10050 0 1 5470
box -12 -8 32 272
use FILL  FILL_6__3109_
timestamp 1701859473
transform -1 0 9830 0 1 5470
box -12 -8 32 272
use FILL  FILL_6__3110_
timestamp 1701859473
transform 1 0 8470 0 -1 6510
box -12 -8 32 272
use FILL  FILL_6__3111_
timestamp 1701859473
transform -1 0 8250 0 -1 6510
box -12 -8 32 272
use FILL  FILL_6__3112_
timestamp 1701859473
transform 1 0 590 0 -1 2870
box -12 -8 32 272
use FILL  FILL_6__3113_
timestamp 1701859473
transform 1 0 130 0 -1 2870
box -12 -8 32 272
use FILL  FILL_6__3114_
timestamp 1701859473
transform -1 0 390 0 -1 2870
box -12 -8 32 272
use FILL  FILL_6__3115_
timestamp 1701859473
transform -1 0 1270 0 1 2350
box -12 -8 32 272
use FILL  FILL_6__3116_
timestamp 1701859473
transform 1 0 1030 0 -1 2350
box -12 -8 32 272
use FILL  FILL_6__3117_
timestamp 1701859473
transform 1 0 2110 0 -1 1310
box -12 -8 32 272
use FILL  FILL_6__3118_
timestamp 1701859473
transform -1 0 1490 0 -1 2350
box -12 -8 32 272
use FILL  FILL_6__3119_
timestamp 1701859473
transform -1 0 1250 0 -1 2350
box -12 -8 32 272
use FILL  FILL_6__3120_
timestamp 1701859473
transform -1 0 550 0 1 2350
box -12 -8 32 272
use FILL  FILL_6__3121_
timestamp 1701859473
transform 1 0 330 0 1 2870
box -12 -8 32 272
use FILL  FILL_6__3122_
timestamp 1701859473
transform 1 0 2590 0 -1 3390
box -12 -8 32 272
use FILL  FILL_6__3123_
timestamp 1701859473
transform 1 0 610 0 1 3390
box -12 -8 32 272
use FILL  FILL_6__3124_
timestamp 1701859473
transform -1 0 390 0 1 3390
box -12 -8 32 272
use FILL  FILL_6__3125_
timestamp 1701859473
transform -1 0 810 0 -1 2350
box -12 -8 32 272
use FILL  FILL_6__3126_
timestamp 1701859473
transform -1 0 1510 0 1 2350
box -12 -8 32 272
use FILL  FILL_6__3127_
timestamp 1701859473
transform -1 0 1030 0 1 2350
box -12 -8 32 272
use FILL  FILL_6__3128_
timestamp 1701859473
transform -1 0 1970 0 1 2350
box -12 -8 32 272
use FILL  FILL_6__3129_
timestamp 1701859473
transform -1 0 1730 0 -1 2350
box -12 -8 32 272
use FILL  FILL_6__3130_
timestamp 1701859473
transform -1 0 1750 0 1 2350
box -12 -8 32 272
use FILL  FILL_6__3131_
timestamp 1701859473
transform -1 0 790 0 1 2350
box -12 -8 32 272
use FILL  FILL_6__3132_
timestamp 1701859473
transform 1 0 550 0 1 2870
box -12 -8 32 272
use FILL  FILL_6__3133_
timestamp 1701859473
transform 1 0 610 0 -1 3910
box -12 -8 32 272
use FILL  FILL_6__3134_
timestamp 1701859473
transform -1 0 1290 0 1 3390
box -12 -8 32 272
use FILL  FILL_6__3135_
timestamp 1701859473
transform 1 0 1050 0 1 3390
box -12 -8 32 272
use FILL  FILL_6__3136_
timestamp 1701859473
transform -1 0 630 0 -1 3390
box -12 -8 32 272
use FILL  FILL_6__3137_
timestamp 1701859473
transform 1 0 350 0 -1 3390
box -12 -8 32 272
use FILL  FILL_6__3138_
timestamp 1701859473
transform -1 0 1750 0 1 4430
box -12 -8 32 272
use FILL  FILL_6__3139_
timestamp 1701859473
transform -1 0 1950 0 -1 3390
box -12 -8 32 272
use FILL  FILL_6__3140_
timestamp 1701859473
transform -1 0 370 0 1 3910
box -12 -8 32 272
use FILL  FILL_6__3141_
timestamp 1701859473
transform 1 0 810 0 1 4430
box -12 -8 32 272
use FILL  FILL_6__3142_
timestamp 1701859473
transform 1 0 1050 0 1 4430
box -12 -8 32 272
use FILL  FILL_6__3143_
timestamp 1701859473
transform 1 0 1070 0 -1 4430
box -12 -8 32 272
use FILL  FILL_6__3144_
timestamp 1701859473
transform -1 0 1310 0 -1 4430
box -12 -8 32 272
use FILL  FILL_6__3145_
timestamp 1701859473
transform -1 0 590 0 1 3910
box -12 -8 32 272
use FILL  FILL_6__3146_
timestamp 1701859473
transform -1 0 810 0 1 3910
box -12 -8 32 272
use FILL  FILL_6__3147_
timestamp 1701859473
transform 1 0 590 0 -1 4430
box -12 -8 32 272
use FILL  FILL_6__3148_
timestamp 1701859473
transform -1 0 850 0 -1 4430
box -12 -8 32 272
use FILL  FILL_6__3149_
timestamp 1701859473
transform -1 0 150 0 -1 3910
box -12 -8 32 272
use FILL  FILL_6__3150_
timestamp 1701859473
transform -1 0 1010 0 1 3910
box -12 -8 32 272
use FILL  FILL_6__3151_
timestamp 1701859473
transform 1 0 130 0 1 3910
box -12 -8 32 272
use FILL  FILL_6__3152_
timestamp 1701859473
transform 1 0 130 0 -1 4430
box -12 -8 32 272
use FILL  FILL_6__3153_
timestamp 1701859473
transform -1 0 370 0 -1 4430
box -12 -8 32 272
use FILL  FILL_6__3154_
timestamp 1701859473
transform -1 0 870 0 -1 3390
box -12 -8 32 272
use FILL  FILL_6__3155_
timestamp 1701859473
transform -1 0 150 0 1 2870
box -12 -8 32 272
use FILL  FILL_6__3156_
timestamp 1701859473
transform 1 0 130 0 -1 3390
box -12 -8 32 272
use FILL  FILL_6__3157_
timestamp 1701859473
transform -1 0 150 0 1 3390
box -12 -8 32 272
use FILL  FILL_6__3158_
timestamp 1701859473
transform 1 0 130 0 1 4430
box -12 -8 32 272
use FILL  FILL_6__3159_
timestamp 1701859473
transform 1 0 350 0 1 4430
box -12 -8 32 272
use FILL  FILL_6__3160_
timestamp 1701859473
transform -1 0 590 0 1 4430
box -12 -8 32 272
use FILL  FILL_6__3161_
timestamp 1701859473
transform 1 0 4230 0 -1 7030
box -12 -8 32 272
use FILL  FILL_6__3162_
timestamp 1701859473
transform -1 0 4470 0 -1 7030
box -12 -8 32 272
use FILL  FILL_6__3163_
timestamp 1701859473
transform 1 0 4690 0 -1 7030
box -12 -8 32 272
use FILL  FILL_6__3164_
timestamp 1701859473
transform 1 0 4930 0 1 7030
box -12 -8 32 272
use FILL  FILL_6__3165_
timestamp 1701859473
transform 1 0 4190 0 1 7550
box -12 -8 32 272
use FILL  FILL_6__3166_
timestamp 1701859473
transform -1 0 4430 0 1 7550
box -12 -8 32 272
use FILL  FILL_6__3167_
timestamp 1701859473
transform 1 0 4910 0 -1 10150
box -12 -8 32 272
use FILL  FILL_6__3168_
timestamp 1701859473
transform 1 0 5110 0 -1 10150
box -12 -8 32 272
use FILL  FILL_6__3169_
timestamp 1701859473
transform -1 0 3750 0 -1 10670
box -12 -8 32 272
use FILL  FILL_6__3170_
timestamp 1701859473
transform -1 0 3970 0 -1 10670
box -12 -8 32 272
use FILL  FILL_6__3171_
timestamp 1701859473
transform 1 0 4390 0 -1 10670
box -12 -8 32 272
use FILL  FILL_6__3172_
timestamp 1701859473
transform -1 0 4630 0 -1 10670
box -12 -8 32 272
use FILL  FILL_6__3173_
timestamp 1701859473
transform 1 0 4230 0 1 10150
box -12 -8 32 272
use FILL  FILL_6__3174_
timestamp 1701859473
transform -1 0 4470 0 1 10150
box -12 -8 32 272
use FILL  FILL_6__3175_
timestamp 1701859473
transform 1 0 5570 0 1 10150
box -12 -8 32 272
use FILL  FILL_6__3176_
timestamp 1701859473
transform 1 0 5330 0 1 10150
box -12 -8 32 272
use FILL  FILL_6__3177_
timestamp 1701859473
transform -1 0 1810 0 -1 5990
box -12 -8 32 272
use FILL  FILL_6__3178_
timestamp 1701859473
transform 1 0 2250 0 -1 5990
box -12 -8 32 272
use FILL  FILL_6__3179_
timestamp 1701859473
transform -1 0 1530 0 1 6510
box -12 -8 32 272
use FILL  FILL_6__3180_
timestamp 1701859473
transform -1 0 1750 0 1 6510
box -12 -8 32 272
use FILL  FILL_6__3181_
timestamp 1701859473
transform -1 0 610 0 -1 6510
box -12 -8 32 272
use FILL  FILL_6__3182_
timestamp 1701859473
transform -1 0 1010 0 -1 6510
box -12 -8 32 272
use FILL  FILL_6__3183_
timestamp 1701859473
transform 1 0 370 0 1 8070
box -12 -8 32 272
use FILL  FILL_6__3184_
timestamp 1701859473
transform -1 0 610 0 1 8070
box -12 -8 32 272
use FILL  FILL_6__3185_
timestamp 1701859473
transform -1 0 150 0 -1 8590
box -12 -8 32 272
use FILL  FILL_6__3186_
timestamp 1701859473
transform -1 0 150 0 1 8070
box -12 -8 32 272
use FILL  FILL_6__3187_
timestamp 1701859473
transform 1 0 770 0 -1 9110
box -12 -8 32 272
use FILL  FILL_6__3188_
timestamp 1701859473
transform 1 0 990 0 -1 9110
box -12 -8 32 272
use FILL  FILL_6__3189_
timestamp 1701859473
transform 1 0 2170 0 -1 9630
box -12 -8 32 272
use FILL  FILL_6__3190_
timestamp 1701859473
transform 1 0 2410 0 1 9110
box -12 -8 32 272
use FILL  FILL_6__3191_
timestamp 1701859473
transform 1 0 1470 0 -1 9110
box -12 -8 32 272
use FILL  FILL_6__3192_
timestamp 1701859473
transform -1 0 1710 0 -1 9110
box -12 -8 32 272
use FILL  FILL_6__3324_
timestamp 1701859473
transform 1 0 5650 0 1 8070
box -12 -8 32 272
use FILL  FILL_6__3325_
timestamp 1701859473
transform -1 0 6370 0 1 8070
box -12 -8 32 272
use FILL  FILL_6__3326_
timestamp 1701859473
transform -1 0 6270 0 -1 8070
box -12 -8 32 272
use FILL  FILL_6__3327_
timestamp 1701859473
transform -1 0 6230 0 -1 8590
box -12 -8 32 272
use FILL  FILL_6__3328_
timestamp 1701859473
transform -1 0 6130 0 1 8070
box -12 -8 32 272
use FILL  FILL_6__3329_
timestamp 1701859473
transform 1 0 5890 0 1 8070
box -12 -8 32 272
use FILL  FILL_6__3330_
timestamp 1701859473
transform -1 0 7070 0 1 8590
box -12 -8 32 272
use FILL  FILL_6__3331_
timestamp 1701859473
transform 1 0 7350 0 -1 8590
box -12 -8 32 272
use FILL  FILL_6__3332_
timestamp 1701859473
transform 1 0 7070 0 -1 8590
box -12 -8 32 272
use FILL  FILL_6__3333_
timestamp 1701859473
transform 1 0 10270 0 1 8590
box -12 -8 32 272
use FILL  FILL_6__3334_
timestamp 1701859473
transform 1 0 9390 0 1 8590
box -12 -8 32 272
use FILL  FILL_6__3335_
timestamp 1701859473
transform 1 0 7930 0 -1 10150
box -12 -8 32 272
use FILL  FILL_6__3336_
timestamp 1701859473
transform -1 0 6770 0 1 9630
box -12 -8 32 272
use FILL  FILL_6__3337_
timestamp 1701859473
transform -1 0 6290 0 1 9630
box -12 -8 32 272
use FILL  FILL_6__3338_
timestamp 1701859473
transform 1 0 7250 0 -1 10150
box -12 -8 32 272
use FILL  FILL_6__3339_
timestamp 1701859473
transform -1 0 8130 0 1 10150
box -12 -8 32 272
use FILL  FILL_6__3340_
timestamp 1701859473
transform 1 0 7890 0 1 10150
box -12 -8 32 272
use FILL  FILL_6__3341_
timestamp 1701859473
transform 1 0 7650 0 1 10150
box -12 -8 32 272
use FILL  FILL_6__3342_
timestamp 1701859473
transform 1 0 6870 0 -1 11190
box -12 -8 32 272
use FILL  FILL_6__3343_
timestamp 1701859473
transform -1 0 7470 0 -1 10150
box -12 -8 32 272
use FILL  FILL_6__3344_
timestamp 1701859473
transform 1 0 7690 0 -1 10150
box -12 -8 32 272
use FILL  FILL_6__3345_
timestamp 1701859473
transform -1 0 9070 0 1 9630
box -12 -8 32 272
use FILL  FILL_6__3346_
timestamp 1701859473
transform 1 0 8590 0 1 10150
box -12 -8 32 272
use FILL  FILL_6__3347_
timestamp 1701859473
transform -1 0 8370 0 1 10150
box -12 -8 32 272
use FILL  FILL_6__3348_
timestamp 1701859473
transform 1 0 9190 0 -1 10670
box -12 -8 32 272
use FILL  FILL_6__3349_
timestamp 1701859473
transform 1 0 7930 0 1 9630
box -12 -8 32 272
use FILL  FILL_6__3350_
timestamp 1701859473
transform 1 0 7630 0 -1 8590
box -12 -8 32 272
use FILL  FILL_6__3351_
timestamp 1701859473
transform -1 0 7810 0 1 8590
box -12 -8 32 272
use FILL  FILL_6__3352_
timestamp 1701859473
transform -1 0 8270 0 -1 9110
box -12 -8 32 272
use FILL  FILL_6__3353_
timestamp 1701859473
transform 1 0 8150 0 -1 10150
box -12 -8 32 272
use FILL  FILL_6__3354_
timestamp 1701859473
transform 1 0 7830 0 -1 10670
box -12 -8 32 272
use FILL  FILL_6__3355_
timestamp 1701859473
transform -1 0 7610 0 -1 10670
box -12 -8 32 272
use FILL  FILL_6__3356_
timestamp 1701859473
transform 1 0 7390 0 -1 10670
box -12 -8 32 272
use FILL  FILL_6__3357_
timestamp 1701859473
transform 1 0 7210 0 1 10670
box -12 -8 32 272
use FILL  FILL_6__3358_
timestamp 1701859473
transform 1 0 7470 0 1 10670
box -12 -8 32 272
use FILL  FILL_6__3359_
timestamp 1701859473
transform 1 0 7710 0 1 10670
box -12 -8 32 272
use FILL  FILL_6__3360_
timestamp 1701859473
transform -1 0 7970 0 1 10670
box -12 -8 32 272
use FILL  FILL_6__3361_
timestamp 1701859473
transform 1 0 8990 0 -1 10670
box -12 -8 32 272
use FILL  FILL_6__3362_
timestamp 1701859473
transform 1 0 8050 0 -1 10670
box -12 -8 32 272
use FILL  FILL_6__3363_
timestamp 1701859473
transform 1 0 8170 0 1 10670
box -12 -8 32 272
use FILL  FILL_6__3364_
timestamp 1701859473
transform 1 0 8010 0 -1 11190
box -12 -8 32 272
use FILL  FILL_6__3365_
timestamp 1701859473
transform -1 0 7550 0 -1 11190
box -12 -8 32 272
use FILL  FILL_6__3366_
timestamp 1701859473
transform 1 0 7070 0 -1 11190
box -12 -8 32 272
use FILL  FILL_6__3367_
timestamp 1701859473
transform 1 0 6950 0 1 10670
box -12 -8 32 272
use FILL  FILL_6__3368_
timestamp 1701859473
transform 1 0 7290 0 -1 11190
box -12 -8 32 272
use FILL  FILL_6__3369_
timestamp 1701859473
transform 1 0 7770 0 -1 11190
box -12 -8 32 272
use FILL  FILL_6__3370_
timestamp 1701859473
transform 1 0 8290 0 -1 10670
box -12 -8 32 272
use FILL  FILL_6__3371_
timestamp 1701859473
transform 1 0 8390 0 1 10670
box -12 -8 32 272
use FILL  FILL_6__3372_
timestamp 1701859473
transform 1 0 9570 0 1 10670
box -12 -8 32 272
use FILL  FILL_6__3373_
timestamp 1701859473
transform -1 0 6670 0 -1 11190
box -12 -8 32 272
use FILL  FILL_6__3374_
timestamp 1701859473
transform 1 0 5770 0 1 10670
box -12 -8 32 272
use FILL  FILL_6__3375_
timestamp 1701859473
transform -1 0 6030 0 1 10670
box -12 -8 32 272
use FILL  FILL_6__3376_
timestamp 1701859473
transform -1 0 6250 0 1 10670
box -12 -8 32 272
use FILL  FILL_6__3377_
timestamp 1701859473
transform 1 0 6490 0 1 10670
box -12 -8 32 272
use FILL  FILL_6__3378_
timestamp 1701859473
transform 1 0 6430 0 -1 11190
box -12 -8 32 272
use FILL  FILL_6__3379_
timestamp 1701859473
transform 1 0 8750 0 -1 10670
box -12 -8 32 272
use FILL  FILL_6__3380_
timestamp 1701859473
transform 1 0 8870 0 1 10670
box -12 -8 32 272
use FILL  FILL_6__3381_
timestamp 1701859473
transform -1 0 6750 0 1 10670
box -12 -8 32 272
use FILL  FILL_6__3382_
timestamp 1701859473
transform 1 0 6210 0 -1 10670
box -12 -8 32 272
use FILL  FILL_6__3383_
timestamp 1701859473
transform -1 0 6470 0 -1 10670
box -12 -8 32 272
use FILL  FILL_6__3384_
timestamp 1701859473
transform -1 0 6910 0 -1 10670
box -12 -8 32 272
use FILL  FILL_6__3385_
timestamp 1701859473
transform 1 0 6670 0 -1 10670
box -12 -8 32 272
use FILL  FILL_6__3386_
timestamp 1701859473
transform 1 0 7150 0 -1 10670
box -12 -8 32 272
use FILL  FILL_6__3387_
timestamp 1701859473
transform 1 0 8510 0 -1 10670
box -12 -8 32 272
use FILL  FILL_6__3388_
timestamp 1701859473
transform 1 0 8630 0 1 10670
box -12 -8 32 272
use FILL  FILL_6__3389_
timestamp 1701859473
transform 1 0 10290 0 -1 10670
box -12 -8 32 272
use FILL  FILL_6__3390_
timestamp 1701859473
transform 1 0 9850 0 -1 10670
box -12 -8 32 272
use FILL  FILL_6__3391_
timestamp 1701859473
transform 1 0 10050 0 -1 10670
box -12 -8 32 272
use FILL  FILL_6__3392_
timestamp 1701859473
transform 1 0 10510 0 -1 10670
box -12 -8 32 272
use FILL  FILL_6__3393_
timestamp 1701859473
transform -1 0 11250 0 -1 10150
box -12 -8 32 272
use FILL  FILL_6__3394_
timestamp 1701859473
transform 1 0 7430 0 1 10150
box -12 -8 32 272
use FILL  FILL_6__3395_
timestamp 1701859473
transform 1 0 6490 0 1 10150
box -12 -8 32 272
use FILL  FILL_6__3396_
timestamp 1701859473
transform -1 0 6750 0 1 10150
box -12 -8 32 272
use FILL  FILL_6__3397_
timestamp 1701859473
transform -1 0 7070 0 -1 10150
box -12 -8 32 272
use FILL  FILL_6__3398_
timestamp 1701859473
transform 1 0 6350 0 -1 10150
box -12 -8 32 272
use FILL  FILL_6__3399_
timestamp 1701859473
transform -1 0 6830 0 -1 10150
box -12 -8 32 272
use FILL  FILL_6__3400_
timestamp 1701859473
transform -1 0 7010 0 1 10150
box -12 -8 32 272
use FILL  FILL_6__3401_
timestamp 1701859473
transform 1 0 7190 0 1 10150
box -12 -8 32 272
use FILL  FILL_6__3402_
timestamp 1701859473
transform -1 0 9130 0 1 10150
box -12 -8 32 272
use FILL  FILL_6__3403_
timestamp 1701859473
transform 1 0 9570 0 1 10150
box -12 -8 32 272
use FILL  FILL_6__3404_
timestamp 1701859473
transform -1 0 5830 0 1 9630
box -12 -8 32 272
use FILL  FILL_6__3405_
timestamp 1701859473
transform -1 0 6110 0 -1 10150
box -12 -8 32 272
use FILL  FILL_6__3406_
timestamp 1701859473
transform 1 0 6470 0 -1 9630
box -12 -8 32 272
use FILL  FILL_6__3407_
timestamp 1701859473
transform -1 0 6690 0 -1 9630
box -12 -8 32 272
use FILL  FILL_6__3408_
timestamp 1701859473
transform 1 0 6950 0 1 9630
box -12 -8 32 272
use FILL  FILL_6__3409_
timestamp 1701859473
transform -1 0 6570 0 -1 10150
box -12 -8 32 272
use FILL  FILL_6__3410_
timestamp 1701859473
transform 1 0 9310 0 -1 10150
box -12 -8 32 272
use FILL  FILL_6__3411_
timestamp 1701859473
transform 1 0 9330 0 1 10150
box -12 -8 32 272
use FILL  FILL_6__3412_
timestamp 1701859473
transform 1 0 10050 0 1 10150
box -12 -8 32 272
use FILL  FILL_6__3413_
timestamp 1701859473
transform -1 0 6070 0 1 9630
box -12 -8 32 272
use FILL  FILL_6__3414_
timestamp 1701859473
transform 1 0 8210 0 1 9110
box -12 -8 32 272
use FILL  FILL_6__3415_
timestamp 1701859473
transform 1 0 6490 0 1 9630
box -12 -8 32 272
use FILL  FILL_6__3416_
timestamp 1701859473
transform 1 0 7330 0 1 8590
box -12 -8 32 272
use FILL  FILL_6__3417_
timestamp 1701859473
transform 1 0 7410 0 -1 9110
box -12 -8 32 272
use FILL  FILL_6__3418_
timestamp 1701859473
transform -1 0 7550 0 -1 9630
box -12 -8 32 272
use FILL  FILL_6__3419_
timestamp 1701859473
transform 1 0 7310 0 -1 9630
box -12 -8 32 272
use FILL  FILL_6__3420_
timestamp 1701859473
transform -1 0 6890 0 -1 9630
box -12 -8 32 272
use FILL  FILL_6__3421_
timestamp 1701859473
transform -1 0 7110 0 -1 9630
box -12 -8 32 272
use FILL  FILL_6__3422_
timestamp 1701859473
transform -1 0 7210 0 1 9630
box -12 -8 32 272
use FILL  FILL_6__3423_
timestamp 1701859473
transform -1 0 8270 0 -1 9630
box -12 -8 32 272
use FILL  FILL_6__3424_
timestamp 1701859473
transform -1 0 7790 0 -1 9630
box -12 -8 32 272
use FILL  FILL_6__3425_
timestamp 1701859473
transform -1 0 7450 0 1 9630
box -12 -8 32 272
use FILL  FILL_6__3426_
timestamp 1701859473
transform -1 0 9090 0 -1 10150
box -12 -8 32 272
use FILL  FILL_6__3427_
timestamp 1701859473
transform 1 0 8850 0 -1 10150
box -12 -8 32 272
use FILL  FILL_6__3428_
timestamp 1701859473
transform 1 0 7530 0 1 8590
box -12 -8 32 272
use FILL  FILL_6__3429_
timestamp 1701859473
transform 1 0 7610 0 -1 9110
box -12 -8 32 272
use FILL  FILL_6__3430_
timestamp 1701859473
transform -1 0 7830 0 -1 9110
box -12 -8 32 272
use FILL  FILL_6__3431_
timestamp 1701859473
transform 1 0 7750 0 1 9110
box -12 -8 32 272
use FILL  FILL_6__3432_
timestamp 1701859473
transform 1 0 7990 0 1 9110
box -12 -8 32 272
use FILL  FILL_6__3433_
timestamp 1701859473
transform -1 0 8030 0 -1 9630
box -12 -8 32 272
use FILL  FILL_6__3434_
timestamp 1701859473
transform 1 0 7670 0 1 9630
box -12 -8 32 272
use FILL  FILL_6__3435_
timestamp 1701859473
transform 1 0 10290 0 1 10150
box -12 -8 32 272
use FILL  FILL_6__3436_
timestamp 1701859473
transform -1 0 10290 0 -1 10150
box -12 -8 32 272
use FILL  FILL_6__3437_
timestamp 1701859473
transform 1 0 10730 0 1 10150
box -12 -8 32 272
use FILL  FILL_6__3438_
timestamp 1701859473
transform 1 0 10510 0 1 10150
box -12 -8 32 272
use FILL  FILL_6__3439_
timestamp 1701859473
transform 1 0 10950 0 1 10150
box -12 -8 32 272
use FILL  FILL_6__3440_
timestamp 1701859473
transform -1 0 10770 0 -1 10150
box -12 -8 32 272
use FILL  FILL_6__3441_
timestamp 1701859473
transform -1 0 10630 0 1 9630
box -12 -8 32 272
use FILL  FILL_6__3442_
timestamp 1701859473
transform -1 0 10510 0 -1 10150
box -12 -8 32 272
use FILL  FILL_6__3443_
timestamp 1701859473
transform -1 0 11070 0 1 9630
box -12 -8 32 272
use FILL  FILL_6__3444_
timestamp 1701859473
transform -1 0 8470 0 -1 9630
box -12 -8 32 272
use FILL  FILL_6__3445_
timestamp 1701859473
transform -1 0 8170 0 1 9630
box -12 -8 32 272
use FILL  FILL_6__3446_
timestamp 1701859473
transform 1 0 8610 0 1 9630
box -12 -8 32 272
use FILL  FILL_6__3447_
timestamp 1701859473
transform 1 0 8390 0 1 9630
box -12 -8 32 272
use FILL  FILL_6__3448_
timestamp 1701859473
transform -1 0 8830 0 1 9630
box -12 -8 32 272
use FILL  FILL_6__3449_
timestamp 1701859473
transform -1 0 9870 0 1 10150
box -12 -8 32 272
use FILL  FILL_6__3450_
timestamp 1701859473
transform -1 0 9830 0 -1 10150
box -12 -8 32 272
use FILL  FILL_6__3451_
timestamp 1701859473
transform 1 0 9550 0 -1 10150
box -12 -8 32 272
use FILL  FILL_6__3452_
timestamp 1701859473
transform -1 0 9290 0 1 9630
box -12 -8 32 272
use FILL  FILL_6__3453_
timestamp 1701859473
transform -1 0 10050 0 -1 10150
box -12 -8 32 272
use FILL  FILL_6__3454_
timestamp 1701859473
transform 1 0 9490 0 1 9630
box -12 -8 32 272
use FILL  FILL_6__3455_
timestamp 1701859473
transform 1 0 9710 0 1 9630
box -12 -8 32 272
use FILL  FILL_6__3456_
timestamp 1701859473
transform -1 0 10410 0 1 9630
box -12 -8 32 272
use FILL  FILL_6__3457_
timestamp 1701859473
transform -1 0 9950 0 1 9630
box -12 -8 32 272
use FILL  FILL_6__3458_
timestamp 1701859473
transform -1 0 10190 0 1 9630
box -12 -8 32 272
use FILL  FILL_6__3459_
timestamp 1701859473
transform -1 0 10330 0 -1 9630
box -12 -8 32 272
use FILL  FILL_6__3460_
timestamp 1701859473
transform 1 0 10990 0 -1 10150
box -12 -8 32 272
use FILL  FILL_6__3461_
timestamp 1701859473
transform -1 0 11230 0 -1 9630
box -12 -8 32 272
use FILL  FILL_6__3462_
timestamp 1701859473
transform -1 0 10770 0 -1 9630
box -12 -8 32 272
use FILL  FILL_6__3463_
timestamp 1701859473
transform 1 0 10450 0 -1 11190
box -12 -8 32 272
use FILL  FILL_6__3464_
timestamp 1701859473
transform 1 0 9790 0 -1 11190
box -12 -8 32 272
use FILL  FILL_6__3465_
timestamp 1701859473
transform 1 0 10030 0 -1 11190
box -12 -8 32 272
use FILL  FILL_6__3466_
timestamp 1701859473
transform 1 0 10210 0 -1 11190
box -12 -8 32 272
use FILL  FILL_6__3467_
timestamp 1701859473
transform -1 0 11190 0 1 10670
box -12 -8 32 272
use FILL  FILL_6__3468_
timestamp 1701859473
transform 1 0 10690 0 1 10670
box -12 -8 32 272
use FILL  FILL_6__3469_
timestamp 1701859473
transform 1 0 9410 0 -1 10670
box -12 -8 32 272
use FILL  FILL_6__3470_
timestamp 1701859473
transform 1 0 9650 0 -1 10670
box -12 -8 32 272
use FILL  FILL_6__3471_
timestamp 1701859473
transform 1 0 9790 0 1 10670
box -12 -8 32 272
use FILL  FILL_6__3472_
timestamp 1701859473
transform -1 0 10050 0 1 10670
box -12 -8 32 272
use FILL  FILL_6__3473_
timestamp 1701859473
transform 1 0 8670 0 -1 11190
box -12 -8 32 272
use FILL  FILL_6__3474_
timestamp 1701859473
transform 1 0 8230 0 -1 11190
box -12 -8 32 272
use FILL  FILL_6__3475_
timestamp 1701859473
transform 1 0 8470 0 -1 11190
box -12 -8 32 272
use FILL  FILL_6__3476_
timestamp 1701859473
transform -1 0 8910 0 -1 11190
box -12 -8 32 272
use FILL  FILL_6__3477_
timestamp 1701859473
transform 1 0 9130 0 -1 11190
box -12 -8 32 272
use FILL  FILL_6__3478_
timestamp 1701859473
transform 1 0 9110 0 1 10670
box -12 -8 32 272
use FILL  FILL_6__3479_
timestamp 1701859473
transform 1 0 8390 0 -1 10150
box -12 -8 32 272
use FILL  FILL_6__3480_
timestamp 1701859473
transform -1 0 8650 0 -1 10150
box -12 -8 32 272
use FILL  FILL_6__3481_
timestamp 1701859473
transform -1 0 8430 0 1 9110
box -12 -8 32 272
use FILL  FILL_6__3482_
timestamp 1701859473
transform -1 0 8650 0 1 9110
box -12 -8 32 272
use FILL  FILL_6__3483_
timestamp 1701859473
transform 1 0 8830 0 1 10150
box -12 -8 32 272
use FILL  FILL_6__3484_
timestamp 1701859473
transform -1 0 10130 0 -1 9630
box -12 -8 32 272
use FILL  FILL_6__3485_
timestamp 1701859473
transform 1 0 11150 0 1 10150
box -12 -8 32 272
use FILL  FILL_6__3486_
timestamp 1701859473
transform 1 0 10490 0 1 9110
box -12 -8 32 272
use FILL  FILL_6__3487_
timestamp 1701859473
transform 1 0 10530 0 -1 9630
box -12 -8 32 272
use FILL  FILL_6__3488_
timestamp 1701859473
transform -1 0 10830 0 1 9630
box -12 -8 32 272
use FILL  FILL_6__3489_
timestamp 1701859473
transform 1 0 10670 0 -1 11190
box -12 -8 32 272
use FILL  FILL_6__3490_
timestamp 1701859473
transform 1 0 11130 0 -1 11190
box -12 -8 32 272
use FILL  FILL_6__3491_
timestamp 1701859473
transform -1 0 10930 0 -1 11190
box -12 -8 32 272
use FILL  FILL_6__3492_
timestamp 1701859473
transform -1 0 10490 0 1 10670
box -12 -8 32 272
use FILL  FILL_6__3493_
timestamp 1701859473
transform -1 0 10270 0 1 10670
box -12 -8 32 272
use FILL  FILL_6__3494_
timestamp 1701859473
transform 1 0 9370 0 1 10670
box -12 -8 32 272
use FILL  FILL_6__3495_
timestamp 1701859473
transform -1 0 9570 0 -1 11190
box -12 -8 32 272
use FILL  FILL_6__3496_
timestamp 1701859473
transform 1 0 9330 0 -1 11190
box -12 -8 32 272
use FILL  FILL_6__3497_
timestamp 1701859473
transform -1 0 9430 0 -1 9630
box -12 -8 32 272
use FILL  FILL_6__3498_
timestamp 1701859473
transform -1 0 8930 0 1 9110
box -12 -8 32 272
use FILL  FILL_6__3499_
timestamp 1701859473
transform 1 0 8450 0 -1 9110
box -12 -8 32 272
use FILL  FILL_6__3500_
timestamp 1701859473
transform 1 0 9830 0 1 9110
box -12 -8 32 272
use FILL  FILL_6__3501_
timestamp 1701859473
transform -1 0 10070 0 1 9110
box -12 -8 32 272
use FILL  FILL_6__3502_
timestamp 1701859473
transform -1 0 8330 0 -1 8590
box -12 -8 32 272
use FILL  FILL_6__3503_
timestamp 1701859473
transform -1 0 8710 0 -1 9630
box -12 -8 32 272
use FILL  FILL_6__3504_
timestamp 1701859473
transform 1 0 8930 0 -1 9630
box -12 -8 32 272
use FILL  FILL_6__3505_
timestamp 1701859473
transform -1 0 9190 0 -1 9630
box -12 -8 32 272
use FILL  FILL_6__3506_
timestamp 1701859473
transform -1 0 8710 0 1 8590
box -12 -8 32 272
use FILL  FILL_6__3507_
timestamp 1701859473
transform 1 0 10790 0 -1 9110
box -12 -8 32 272
use FILL  FILL_6__3508_
timestamp 1701859473
transform 1 0 10550 0 -1 9110
box -12 -8 32 272
use FILL  FILL_6__3509_
timestamp 1701859473
transform 1 0 8490 0 1 8590
box -12 -8 32 272
use FILL  FILL_6__3510_
timestamp 1701859473
transform -1 0 8950 0 1 8590
box -12 -8 32 272
use FILL  FILL_6__3511_
timestamp 1701859473
transform 1 0 10010 0 -1 270
box -12 -8 32 272
use FILL  FILL_6__3512_
timestamp 1701859473
transform 1 0 11010 0 -1 9110
box -12 -8 32 272
use FILL  FILL_6__3513_
timestamp 1701859473
transform 1 0 10990 0 -1 9630
box -12 -8 32 272
use FILL  FILL_6__3514_
timestamp 1701859473
transform 1 0 10950 0 1 10670
box -12 -8 32 272
use FILL  FILL_6__3515_
timestamp 1701859473
transform -1 0 10750 0 -1 10670
box -12 -8 32 272
use FILL  FILL_6__3516_
timestamp 1701859473
transform 1 0 10970 0 -1 10670
box -12 -8 32 272
use FILL  FILL_6__3517_
timestamp 1701859473
transform 1 0 9650 0 -1 9630
box -12 -8 32 272
use FILL  FILL_6__3518_
timestamp 1701859473
transform 1 0 9870 0 -1 9630
box -12 -8 32 272
use FILL  FILL_6__3519_
timestamp 1701859473
transform 1 0 9150 0 1 9110
box -12 -8 32 272
use FILL  FILL_6__3520_
timestamp 1701859473
transform -1 0 9390 0 1 9110
box -12 -8 32 272
use FILL  FILL_6__3521_
timestamp 1701859473
transform 1 0 6630 0 1 8590
box -12 -8 32 272
use FILL  FILL_6__3522_
timestamp 1701859473
transform 1 0 8030 0 -1 9110
box -12 -8 32 272
use FILL  FILL_6__3523_
timestamp 1701859473
transform 1 0 6830 0 1 8590
box -12 -8 32 272
use FILL  FILL_6__3524_
timestamp 1701859473
transform 1 0 7550 0 1 9110
box -12 -8 32 272
use FILL  FILL_6__3525_
timestamp 1701859473
transform 1 0 7090 0 1 9110
box -12 -8 32 272
use FILL  FILL_6__3526_
timestamp 1701859473
transform -1 0 7330 0 1 9110
box -12 -8 32 272
use FILL  FILL_6__3539_
timestamp 1701859473
transform 1 0 11190 0 -1 7030
box -12 -8 32 272
use FILL  FILL_6__3540_
timestamp 1701859473
transform 1 0 4690 0 1 10670
box -12 -8 32 272
use FILL  FILL_6__3541_
timestamp 1701859473
transform -1 0 150 0 1 5990
box -12 -8 32 272
use FILL  FILL_6__3542_
timestamp 1701859473
transform -1 0 150 0 -1 8070
box -12 -8 32 272
use FILL  FILL_6__3543_
timestamp 1701859473
transform -1 0 150 0 1 8590
box -12 -8 32 272
use FILL  FILL_6__3544_
timestamp 1701859473
transform -1 0 150 0 1 9110
box -12 -8 32 272
use FILL  FILL_6__3545_
timestamp 1701859473
transform -1 0 1990 0 -1 11190
box -12 -8 32 272
use FILL  FILL_6__3546_
timestamp 1701859473
transform -1 0 610 0 1 9110
box -12 -8 32 272
use FILL  FILL_6__3547_
timestamp 1701859473
transform 1 0 4730 0 -1 11190
box -12 -8 32 272
use FILL  FILL_6__3548_
timestamp 1701859473
transform 1 0 5330 0 1 10670
box -12 -8 32 272
use FILL  FILL_6__3549_
timestamp 1701859473
transform -1 0 4330 0 -1 11190
box -12 -8 32 272
use FILL  FILL_6__3550_
timestamp 1701859473
transform -1 0 5170 0 -1 11190
box -12 -8 32 272
use FILL  FILL_6__3551_
timestamp 1701859473
transform 1 0 5570 0 -1 11190
box -12 -8 32 272
use FILL  FILL_6__3552_
timestamp 1701859473
transform 1 0 5350 0 -1 11190
box -12 -8 32 272
use FILL  FILL_6__3553_
timestamp 1701859473
transform -1 0 150 0 -1 5990
box -12 -8 32 272
use FILL  FILL_6__3554_
timestamp 1701859473
transform -1 0 350 0 1 7030
box -12 -8 32 272
use FILL  FILL_6__3555_
timestamp 1701859473
transform -1 0 5130 0 1 10670
box -12 -8 32 272
use FILL  FILL_6__3556_
timestamp 1701859473
transform 1 0 6270 0 1 10150
box -12 -8 32 272
use FILL  FILL_6__3557_
timestamp 1701859473
transform -1 0 5810 0 -1 11190
box -12 -8 32 272
use FILL  FILL_6__3558_
timestamp 1701859473
transform 1 0 6210 0 -1 11190
box -12 -8 32 272
use FILL  FILL_6__3559_
timestamp 1701859473
transform -1 0 4870 0 -1 10670
box -12 -8 32 272
use FILL  FILL_6__3560_
timestamp 1701859473
transform 1 0 5550 0 1 10670
box -12 -8 32 272
use FILL  FILL_6__3561_
timestamp 1701859473
transform 1 0 5990 0 -1 11190
box -12 -8 32 272
use FILL  FILL_6__3562_
timestamp 1701859473
transform 1 0 5790 0 1 10150
box -12 -8 32 272
use FILL  FILL_6__3563_
timestamp 1701859473
transform 1 0 5250 0 1 3390
box -12 -8 32 272
use FILL  FILL_6_BUFX2_insert0
timestamp 1701859473
transform 1 0 5870 0 -1 10150
box -12 -8 32 272
use FILL  FILL_6_BUFX2_insert1
timestamp 1701859473
transform 1 0 6630 0 1 2350
box -12 -8 32 272
use FILL  FILL_6_BUFX2_insert2
timestamp 1701859473
transform 1 0 5470 0 -1 1830
box -12 -8 32 272
use FILL  FILL_6_BUFX2_insert3
timestamp 1701859473
transform -1 0 610 0 -1 5470
box -12 -8 32 272
use FILL  FILL_6_BUFX2_insert4
timestamp 1701859473
transform 1 0 3350 0 1 4950
box -12 -8 32 272
use FILL  FILL_6_BUFX2_insert5
timestamp 1701859473
transform 1 0 1410 0 -1 1830
box -12 -8 32 272
use FILL  FILL_6_BUFX2_insert6
timestamp 1701859473
transform -1 0 150 0 -1 11190
box -12 -8 32 272
use FILL  FILL_6_BUFX2_insert7
timestamp 1701859473
transform 1 0 1710 0 1 10670
box -12 -8 32 272
use FILL  FILL_6_BUFX2_insert8
timestamp 1701859473
transform 1 0 1670 0 1 1830
box -12 -8 32 272
use FILL  FILL_6_BUFX2_insert9
timestamp 1701859473
transform 1 0 1970 0 -1 3910
box -12 -8 32 272
use FILL  FILL_6_BUFX2_insert10
timestamp 1701859473
transform 1 0 1790 0 -1 4430
box -12 -8 32 272
use FILL  FILL_6_BUFX2_insert11
timestamp 1701859473
transform -1 0 1770 0 -1 3910
box -12 -8 32 272
use FILL  FILL_6_BUFX2_insert12
timestamp 1701859473
transform -1 0 1550 0 -1 3910
box -12 -8 32 272
use FILL  FILL_6_BUFX2_insert13
timestamp 1701859473
transform -1 0 1450 0 -1 1310
box -12 -8 32 272
use FILL  FILL_6_BUFX2_insert14
timestamp 1701859473
transform -1 0 3690 0 1 3390
box -12 -8 32 272
use FILL  FILL_6_BUFX2_insert15
timestamp 1701859473
transform 1 0 4570 0 -1 5470
box -12 -8 32 272
use FILL  FILL_6_BUFX2_insert16
timestamp 1701859473
transform 1 0 1370 0 -1 4950
box -12 -8 32 272
use FILL  FILL_6_BUFX2_insert17
timestamp 1701859473
transform 1 0 3650 0 1 1310
box -12 -8 32 272
use FILL  FILL_6_BUFX2_insert18
timestamp 1701859473
transform -1 0 9790 0 1 2350
box -12 -8 32 272
use FILL  FILL_6_BUFX2_insert19
timestamp 1701859473
transform -1 0 8530 0 -1 790
box -12 -8 32 272
use FILL  FILL_6_BUFX2_insert20
timestamp 1701859473
transform 1 0 9990 0 1 2350
box -12 -8 32 272
use FILL  FILL_6_BUFX2_insert21
timestamp 1701859473
transform -1 0 7830 0 -1 1310
box -12 -8 32 272
use FILL  FILL_6_BUFX2_insert22
timestamp 1701859473
transform -1 0 3230 0 -1 2870
box -12 -8 32 272
use FILL  FILL_6_BUFX2_insert23
timestamp 1701859473
transform -1 0 2770 0 -1 4950
box -12 -8 32 272
use FILL  FILL_6_BUFX2_insert24
timestamp 1701859473
transform -1 0 3670 0 -1 4430
box -12 -8 32 272
use FILL  FILL_6_BUFX2_insert25
timestamp 1701859473
transform 1 0 4410 0 1 4430
box -12 -8 32 272
use FILL  FILL_6_BUFX2_insert26
timestamp 1701859473
transform 1 0 4230 0 1 2870
box -12 -8 32 272
use FILL  FILL_6_BUFX2_insert27
timestamp 1701859473
transform 1 0 9630 0 1 4950
box -12 -8 32 272
use FILL  FILL_6_BUFX2_insert28
timestamp 1701859473
transform -1 0 7510 0 -1 5990
box -12 -8 32 272
use FILL  FILL_6_BUFX2_insert29
timestamp 1701859473
transform -1 0 1310 0 1 6510
box -12 -8 32 272
use FILL  FILL_6_BUFX2_insert30
timestamp 1701859473
transform -1 0 8810 0 -1 3910
box -12 -8 32 272
use FILL  FILL_6_BUFX2_insert31
timestamp 1701859473
transform -1 0 9590 0 1 3910
box -12 -8 32 272
use FILL  FILL_6_BUFX2_insert32
timestamp 1701859473
transform 1 0 5890 0 -1 3910
box -12 -8 32 272
use FILL  FILL_6_BUFX2_insert33
timestamp 1701859473
transform -1 0 9570 0 -1 4950
box -12 -8 32 272
use FILL  FILL_6_BUFX2_insert34
timestamp 1701859473
transform 1 0 5230 0 1 8590
box -12 -8 32 272
use FILL  FILL_6_BUFX2_insert35
timestamp 1701859473
transform -1 0 5990 0 1 7550
box -12 -8 32 272
use FILL  FILL_6_BUFX2_insert36
timestamp 1701859473
transform -1 0 1230 0 1 8590
box -12 -8 32 272
use FILL  FILL_6_BUFX2_insert37
timestamp 1701859473
transform -1 0 9610 0 1 8590
box -12 -8 32 272
use FILL  FILL_6_BUFX2_insert49
timestamp 1701859473
transform -1 0 3070 0 1 6510
box -12 -8 32 272
use FILL  FILL_6_BUFX2_insert50
timestamp 1701859473
transform 1 0 2370 0 -1 8590
box -12 -8 32 272
use FILL  FILL_6_BUFX2_insert51
timestamp 1701859473
transform 1 0 3230 0 -1 8590
box -12 -8 32 272
use FILL  FILL_6_BUFX2_insert52
timestamp 1701859473
transform 1 0 3410 0 1 5470
box -12 -8 32 272
use FILL  FILL_6_BUFX2_insert53
timestamp 1701859473
transform -1 0 11250 0 1 9110
box -12 -8 32 272
use FILL  FILL_6_BUFX2_insert54
timestamp 1701859473
transform -1 0 9190 0 1 8590
box -12 -8 32 272
use FILL  FILL_6_BUFX2_insert55
timestamp 1701859473
transform -1 0 9630 0 1 9110
box -12 -8 32 272
use FILL  FILL_6_BUFX2_insert56
timestamp 1701859473
transform -1 0 10290 0 1 9110
box -12 -8 32 272
use FILL  FILL_6_BUFX2_insert57
timestamp 1701859473
transform -1 0 11250 0 -1 2350
box -12 -8 32 272
use FILL  FILL_6_BUFX2_insert58
timestamp 1701859473
transform -1 0 8990 0 1 2870
box -12 -8 32 272
use FILL  FILL_6_BUFX2_insert59
timestamp 1701859473
transform -1 0 7570 0 1 1830
box -12 -8 32 272
use FILL  FILL_6_BUFX2_insert60
timestamp 1701859473
transform 1 0 10910 0 1 1830
box -12 -8 32 272
use FILL  FILL_6_BUFX2_insert61
timestamp 1701859473
transform -1 0 11190 0 1 2870
box -12 -8 32 272
use FILL  FILL_6_BUFX2_insert62
timestamp 1701859473
transform 1 0 2230 0 1 3910
box -12 -8 32 272
use FILL  FILL_6_BUFX2_insert63
timestamp 1701859473
transform 1 0 2150 0 1 3390
box -12 -8 32 272
use FILL  FILL_6_BUFX2_insert64
timestamp 1701859473
transform -1 0 1810 0 1 3910
box -12 -8 32 272
use FILL  FILL_6_BUFX2_insert65
timestamp 1701859473
transform -1 0 1750 0 1 3390
box -12 -8 32 272
use FILL  FILL_6_BUFX2_insert66
timestamp 1701859473
transform -1 0 4330 0 1 1310
box -12 -8 32 272
use FILL  FILL_6_BUFX2_insert67
timestamp 1701859473
transform -1 0 3630 0 -1 10150
box -12 -8 32 272
use FILL  FILL_6_BUFX2_insert68
timestamp 1701859473
transform -1 0 7190 0 1 2870
box -12 -8 32 272
use FILL  FILL_6_BUFX2_insert69
timestamp 1701859473
transform -1 0 5670 0 -1 3390
box -12 -8 32 272
use FILL  FILL_6_BUFX2_insert70
timestamp 1701859473
transform -1 0 3690 0 -1 1830
box -12 -8 32 272
use FILL  FILL_6_BUFX2_insert71
timestamp 1701859473
transform -1 0 7330 0 1 2350
box -12 -8 32 272
use FILL  FILL_6_BUFX2_insert72
timestamp 1701859473
transform -1 0 6510 0 1 1310
box -12 -8 32 272
use FILL  FILL_6_BUFX2_insert73
timestamp 1701859473
transform 1 0 3630 0 1 5470
box -12 -8 32 272
use FILL  FILL_6_BUFX2_insert74
timestamp 1701859473
transform 1 0 7590 0 -1 2350
box -12 -8 32 272
use FILL  FILL_6_BUFX2_insert75
timestamp 1701859473
transform 1 0 7610 0 1 2870
box -12 -8 32 272
use FILL  FILL_6_BUFX2_insert76
timestamp 1701859473
transform 1 0 7390 0 1 2870
box -12 -8 32 272
use FILL  FILL_6_BUFX2_insert77
timestamp 1701859473
transform -1 0 3450 0 -1 2870
box -12 -8 32 272
use FILL  FILL_6_BUFX2_insert78
timestamp 1701859473
transform 1 0 1950 0 -1 2870
box -12 -8 32 272
use FILL  FILL_6_BUFX2_insert79
timestamp 1701859473
transform -1 0 2190 0 -1 2870
box -12 -8 32 272
use FILL  FILL_6_BUFX2_insert80
timestamp 1701859473
transform 1 0 2430 0 1 4430
box -12 -8 32 272
use FILL  FILL_6_BUFX2_insert81
timestamp 1701859473
transform -1 0 2030 0 1 3910
box -12 -8 32 272
use FILL  FILL_6_BUFX2_insert82
timestamp 1701859473
transform -1 0 350 0 1 8590
box -12 -8 32 272
use FILL  FILL_6_BUFX2_insert83
timestamp 1701859473
transform 1 0 4230 0 -1 10150
box -12 -8 32 272
use FILL  FILL_6_BUFX2_insert84
timestamp 1701859473
transform 1 0 4190 0 -1 7550
box -12 -8 32 272
use FILL  FILL_6_BUFX2_insert85
timestamp 1701859473
transform -1 0 150 0 -1 6510
box -12 -8 32 272
use FILL  FILL_6_BUFX2_insert86
timestamp 1701859473
transform 1 0 1950 0 -1 10150
box -12 -8 32 272
use FILL  FILL_6_CLKBUF1_insert38
timestamp 1701859473
transform 1 0 2950 0 -1 7550
box -12 -8 32 272
use FILL  FILL_6_CLKBUF1_insert39
timestamp 1701859473
transform -1 0 4750 0 -1 6510
box -12 -8 32 272
use FILL  FILL_6_CLKBUF1_insert40
timestamp 1701859473
transform -1 0 1050 0 -1 4950
box -12 -8 32 272
use FILL  FILL_6_CLKBUF1_insert41
timestamp 1701859473
transform -1 0 10710 0 -1 270
box -12 -8 32 272
use FILL  FILL_6_CLKBUF1_insert42
timestamp 1701859473
transform 1 0 9770 0 -1 4950
box -12 -8 32 272
use FILL  FILL_6_CLKBUF1_insert43
timestamp 1701859473
transform -1 0 11090 0 1 7030
box -12 -8 32 272
use FILL  FILL_6_CLKBUF1_insert44
timestamp 1701859473
transform -1 0 10830 0 1 4430
box -12 -8 32 272
use FILL  FILL_6_CLKBUF1_insert45
timestamp 1701859473
transform 1 0 5750 0 -1 6510
box -12 -8 32 272
use FILL  FILL_6_CLKBUF1_insert46
timestamp 1701859473
transform 1 0 4070 0 1 5990
box -12 -8 32 272
use FILL  FILL_6_CLKBUF1_insert47
timestamp 1701859473
transform -1 0 2190 0 1 7550
box -12 -8 32 272
use FILL  FILL_6_CLKBUF1_insert48
timestamp 1701859473
transform -1 0 10870 0 -1 7030
box -12 -8 32 272
use FILL  FILL_7__1669_
timestamp 1701859473
transform -1 0 6870 0 -1 790
box -12 -8 32 272
use FILL  FILL_7__1670_
timestamp 1701859473
transform 1 0 6650 0 -1 2870
box -12 -8 32 272
use FILL  FILL_7__1671_
timestamp 1701859473
transform -1 0 6450 0 -1 8590
box -12 -8 32 272
use FILL  FILL_7__1672_
timestamp 1701859473
transform 1 0 6010 0 -1 10670
box -12 -8 32 272
use FILL  FILL_7__1673_
timestamp 1701859473
transform 1 0 6410 0 1 8590
box -12 -8 32 272
use FILL  FILL_7__1674_
timestamp 1701859473
transform -1 0 6490 0 -1 9110
box -12 -8 32 272
use FILL  FILL_7__1676_
timestamp 1701859473
transform -1 0 390 0 -1 5470
box -12 -8 32 272
use FILL  FILL_7__1677_
timestamp 1701859473
transform -1 0 630 0 1 5470
box -12 -8 32 272
use FILL  FILL_7__1678_
timestamp 1701859473
transform 1 0 150 0 -1 10670
box -12 -8 32 272
use FILL  FILL_7__1679_
timestamp 1701859473
transform -1 0 370 0 -1 11190
box -12 -8 32 272
use FILL  FILL_7__1680_
timestamp 1701859473
transform 1 0 350 0 -1 10670
box -12 -8 32 272
use FILL  FILL_7__1681_
timestamp 1701859473
transform -1 0 170 0 -1 7030
box -12 -8 32 272
use FILL  FILL_7__1683_
timestamp 1701859473
transform 1 0 150 0 1 6510
box -12 -8 32 272
use FILL  FILL_7__1684_
timestamp 1701859473
transform 1 0 1030 0 -1 11190
box -12 -8 32 272
use FILL  FILL_7__1685_
timestamp 1701859473
transform -1 0 1290 0 -1 11190
box -12 -8 32 272
use FILL  FILL_7__1686_
timestamp 1701859473
transform -1 0 1090 0 1 10670
box -12 -8 32 272
use FILL  FILL_7__1687_
timestamp 1701859473
transform 1 0 1510 0 -1 11190
box -12 -8 32 272
use FILL  FILL_7__1688_
timestamp 1701859473
transform -1 0 1770 0 -1 11190
box -12 -8 32 272
use FILL  FILL_7__1689_
timestamp 1701859473
transform -1 0 2030 0 1 10150
box -12 -8 32 272
use FILL  FILL_7__1691_
timestamp 1701859473
transform -1 0 2210 0 -1 9110
box -12 -8 32 272
use FILL  FILL_7__1692_
timestamp 1701859473
transform 1 0 150 0 1 790
box -12 -8 32 272
use FILL  FILL_7__1693_
timestamp 1701859473
transform 1 0 150 0 -1 1310
box -12 -8 32 272
use FILL  FILL_7__1694_
timestamp 1701859473
transform 1 0 570 0 -1 270
box -12 -8 32 272
use FILL  FILL_7__1695_
timestamp 1701859473
transform -1 0 790 0 -1 270
box -12 -8 32 272
use FILL  FILL_7__1696_
timestamp 1701859473
transform 1 0 1210 0 1 2870
box -12 -8 32 272
use FILL  FILL_7__1698_
timestamp 1701859473
transform -1 0 1970 0 1 3390
box -12 -8 32 272
use FILL  FILL_7__1699_
timestamp 1701859473
transform 1 0 3890 0 1 3390
box -12 -8 32 272
use FILL  FILL_7__1700_
timestamp 1701859473
transform -1 0 2690 0 -1 3910
box -12 -8 32 272
use FILL  FILL_7__1701_
timestamp 1701859473
transform -1 0 1230 0 1 270
box -12 -8 32 272
use FILL  FILL_7__1702_
timestamp 1701859473
transform 1 0 990 0 1 270
box -12 -8 32 272
use FILL  FILL_7__1703_
timestamp 1701859473
transform -1 0 1470 0 1 1830
box -12 -8 32 272
use FILL  FILL_7__1705_
timestamp 1701859473
transform 1 0 9850 0 -1 790
box -12 -8 32 272
use FILL  FILL_7__1706_
timestamp 1701859473
transform -1 0 8070 0 -1 4950
box -12 -8 32 272
use FILL  FILL_7__1707_
timestamp 1701859473
transform 1 0 8510 0 -1 4950
box -12 -8 32 272
use FILL  FILL_7__1708_
timestamp 1701859473
transform 1 0 5130 0 -1 5990
box -12 -8 32 272
use FILL  FILL_7__1709_
timestamp 1701859473
transform -1 0 11230 0 1 5990
box -12 -8 32 272
use FILL  FILL_7__1710_
timestamp 1701859473
transform 1 0 5510 0 -1 5470
box -12 -8 32 272
use FILL  FILL_7__1712_
timestamp 1701859473
transform -1 0 5170 0 1 5470
box -12 -8 32 272
use FILL  FILL_7__1713_
timestamp 1701859473
transform 1 0 8030 0 1 4430
box -12 -8 32 272
use FILL  FILL_7__1714_
timestamp 1701859473
transform 1 0 7830 0 1 4950
box -12 -8 32 272
use FILL  FILL_7__1715_
timestamp 1701859473
transform -1 0 8070 0 1 4950
box -12 -8 32 272
use FILL  FILL_7__1716_
timestamp 1701859473
transform -1 0 8290 0 1 4430
box -12 -8 32 272
use FILL  FILL_7__1717_
timestamp 1701859473
transform -1 0 8070 0 1 1310
box -12 -8 32 272
use FILL  FILL_7__1718_
timestamp 1701859473
transform -1 0 6010 0 1 5990
box -12 -8 32 272
use FILL  FILL_7__1720_
timestamp 1701859473
transform -1 0 6850 0 1 5470
box -12 -8 32 272
use FILL  FILL_7__1721_
timestamp 1701859473
transform -1 0 7090 0 1 5470
box -12 -8 32 272
use FILL  FILL_7__1722_
timestamp 1701859473
transform -1 0 7790 0 1 4430
box -12 -8 32 272
use FILL  FILL_7__1723_
timestamp 1701859473
transform 1 0 8010 0 1 1830
box -12 -8 32 272
use FILL  FILL_7__1724_
timestamp 1701859473
transform -1 0 8050 0 -1 1310
box -12 -8 32 272
use FILL  FILL_7__1725_
timestamp 1701859473
transform 1 0 6650 0 1 5990
box -12 -8 32 272
use FILL  FILL_7__1727_
timestamp 1701859473
transform -1 0 7090 0 1 5990
box -12 -8 32 272
use FILL  FILL_7__1728_
timestamp 1701859473
transform 1 0 7790 0 1 5990
box -12 -8 32 272
use FILL  FILL_7__1729_
timestamp 1701859473
transform -1 0 7730 0 -1 5990
box -12 -8 32 272
use FILL  FILL_7__1730_
timestamp 1701859473
transform -1 0 8210 0 1 3390
box -12 -8 32 272
use FILL  FILL_7__1731_
timestamp 1701859473
transform -1 0 8070 0 -1 270
box -12 -8 32 272
use FILL  FILL_7__1732_
timestamp 1701859473
transform -1 0 8030 0 1 5470
box -12 -8 32 272
use FILL  FILL_7__1734_
timestamp 1701859473
transform 1 0 8210 0 -1 5470
box -12 -8 32 272
use FILL  FILL_7__1735_
timestamp 1701859473
transform 1 0 8670 0 -1 5470
box -12 -8 32 272
use FILL  FILL_7__1736_
timestamp 1701859473
transform 1 0 8510 0 1 4950
box -12 -8 32 272
use FILL  FILL_7__1737_
timestamp 1701859473
transform -1 0 8590 0 -1 3910
box -12 -8 32 272
use FILL  FILL_7__1738_
timestamp 1701859473
transform 1 0 8990 0 1 790
box -12 -8 32 272
use FILL  FILL_7__1739_
timestamp 1701859473
transform -1 0 9210 0 -1 790
box -12 -8 32 272
use FILL  FILL_7__1740_
timestamp 1701859473
transform 1 0 6570 0 1 270
box -12 -8 32 272
use FILL  FILL_7__1742_
timestamp 1701859473
transform -1 0 6410 0 -1 790
box -12 -8 32 272
use FILL  FILL_7__1743_
timestamp 1701859473
transform -1 0 2410 0 -1 3390
box -12 -8 32 272
use FILL  FILL_7__1744_
timestamp 1701859473
transform 1 0 390 0 -1 4950
box -12 -8 32 272
use FILL  FILL_7__1745_
timestamp 1701859473
transform 1 0 2210 0 -1 3910
box -12 -8 32 272
use FILL  FILL_7__1746_
timestamp 1701859473
transform -1 0 5230 0 -1 3390
box -12 -8 32 272
use FILL  FILL_7__1747_
timestamp 1701859473
transform -1 0 390 0 -1 270
box -12 -8 32 272
use FILL  FILL_7__1749_
timestamp 1701859473
transform -1 0 1030 0 1 1310
box -12 -8 32 272
use FILL  FILL_7__1750_
timestamp 1701859473
transform -1 0 1250 0 1 1310
box -12 -8 32 272
use FILL  FILL_7__1751_
timestamp 1701859473
transform -1 0 4610 0 -1 2870
box -12 -8 32 272
use FILL  FILL_7__1752_
timestamp 1701859473
transform 1 0 4810 0 -1 2870
box -12 -8 32 272
use FILL  FILL_7__1753_
timestamp 1701859473
transform -1 0 4430 0 1 790
box -12 -8 32 272
use FILL  FILL_7__1754_
timestamp 1701859473
transform 1 0 370 0 -1 790
box -12 -8 32 272
use FILL  FILL_7__1756_
timestamp 1701859473
transform -1 0 170 0 -1 270
box -12 -8 32 272
use FILL  FILL_7__1757_
timestamp 1701859473
transform 1 0 770 0 -1 790
box -12 -8 32 272
use FILL  FILL_7__1758_
timestamp 1701859473
transform 1 0 150 0 1 2350
box -12 -8 32 272
use FILL  FILL_7__1759_
timestamp 1701859473
transform -1 0 2650 0 -1 2870
box -12 -8 32 272
use FILL  FILL_7__1760_
timestamp 1701859473
transform 1 0 3030 0 -1 2870
box -12 -8 32 272
use FILL  FILL_7__1761_
timestamp 1701859473
transform -1 0 3350 0 -1 3390
box -12 -8 32 272
use FILL  FILL_7__1763_
timestamp 1701859473
transform 1 0 150 0 -1 790
box -12 -8 32 272
use FILL  FILL_7__1764_
timestamp 1701859473
transform 1 0 590 0 1 1310
box -12 -8 32 272
use FILL  FILL_7__1765_
timestamp 1701859473
transform 1 0 1450 0 1 1310
box -12 -8 32 272
use FILL  FILL_7__1766_
timestamp 1701859473
transform -1 0 3250 0 -1 1830
box -12 -8 32 272
use FILL  FILL_7__1767_
timestamp 1701859473
transform 1 0 1550 0 -1 4430
box -12 -8 32 272
use FILL  FILL_7__1768_
timestamp 1701859473
transform 1 0 370 0 -1 1310
box -12 -8 32 272
use FILL  FILL_7__1769_
timestamp 1701859473
transform -1 0 590 0 1 1830
box -12 -8 32 272
use FILL  FILL_7__1771_
timestamp 1701859473
transform -1 0 2450 0 -1 3910
box -12 -8 32 272
use FILL  FILL_7__1772_
timestamp 1701859473
transform -1 0 3110 0 -1 3910
box -12 -8 32 272
use FILL  FILL_7__1773_
timestamp 1701859473
transform 1 0 4010 0 1 2870
box -12 -8 32 272
use FILL  FILL_7__1774_
timestamp 1701859473
transform -1 0 5390 0 -1 2350
box -12 -8 32 272
use FILL  FILL_7__1775_
timestamp 1701859473
transform 1 0 350 0 1 790
box -12 -8 32 272
use FILL  FILL_7__1776_
timestamp 1701859473
transform -1 0 390 0 1 1310
box -12 -8 32 272
use FILL  FILL_7__1778_
timestamp 1701859473
transform -1 0 4530 0 1 5470
box -12 -8 32 272
use FILL  FILL_7__1779_
timestamp 1701859473
transform -1 0 6170 0 -1 5470
box -12 -8 32 272
use FILL  FILL_7__1780_
timestamp 1701859473
transform 1 0 4890 0 1 2870
box -12 -8 32 272
use FILL  FILL_7__1781_
timestamp 1701859473
transform 1 0 4470 0 1 2870
box -12 -8 32 272
use FILL  FILL_7__1782_
timestamp 1701859473
transform -1 0 170 0 1 1310
box -12 -8 32 272
use FILL  FILL_7__1783_
timestamp 1701859473
transform -1 0 1450 0 1 2870
box -12 -8 32 272
use FILL  FILL_7__1785_
timestamp 1701859473
transform 1 0 5070 0 -1 2870
box -12 -8 32 272
use FILL  FILL_7__1786_
timestamp 1701859473
transform -1 0 5150 0 -1 2350
box -12 -8 32 272
use FILL  FILL_7__1787_
timestamp 1701859473
transform 1 0 5130 0 1 2350
box -12 -8 32 272
use FILL  FILL_7__1788_
timestamp 1701859473
transform -1 0 4930 0 -1 2350
box -12 -8 32 272
use FILL  FILL_7__1789_
timestamp 1701859473
transform 1 0 150 0 1 1830
box -12 -8 32 272
use FILL  FILL_7__1790_
timestamp 1701859473
transform -1 0 390 0 -1 2350
box -12 -8 32 272
use FILL  FILL_7__1791_
timestamp 1701859473
transform -1 0 2190 0 -1 2350
box -12 -8 32 272
use FILL  FILL_7__1793_
timestamp 1701859473
transform -1 0 4670 0 1 1830
box -12 -8 32 272
use FILL  FILL_7__1794_
timestamp 1701859473
transform 1 0 990 0 1 1830
box -12 -8 32 272
use FILL  FILL_7__1795_
timestamp 1701859473
transform -1 0 2250 0 1 2350
box -12 -8 32 272
use FILL  FILL_7__1796_
timestamp 1701859473
transform -1 0 1870 0 -1 1830
box -12 -8 32 272
use FILL  FILL_7__1797_
timestamp 1701859473
transform 1 0 2090 0 -1 1830
box -12 -8 32 272
use FILL  FILL_7__1798_
timestamp 1701859473
transform 1 0 1010 0 -1 1310
box -12 -8 32 272
use FILL  FILL_7__1800_
timestamp 1701859473
transform 1 0 3510 0 1 1830
box -12 -8 32 272
use FILL  FILL_7__1801_
timestamp 1701859473
transform -1 0 1250 0 1 1830
box -12 -8 32 272
use FILL  FILL_7__1802_
timestamp 1701859473
transform -1 0 3790 0 1 2350
box -12 -8 32 272
use FILL  FILL_7__1803_
timestamp 1701859473
transform -1 0 4010 0 1 2350
box -12 -8 32 272
use FILL  FILL_7__1804_
timestamp 1701859473
transform -1 0 4250 0 1 2350
box -12 -8 32 272
use FILL  FILL_7__1805_
timestamp 1701859473
transform 1 0 5550 0 1 2350
box -12 -8 32 272
use FILL  FILL_7__1807_
timestamp 1701859473
transform -1 0 5350 0 1 2350
box -12 -8 32 272
use FILL  FILL_7__1808_
timestamp 1701859473
transform 1 0 4870 0 1 1830
box -12 -8 32 272
use FILL  FILL_7__1809_
timestamp 1701859473
transform -1 0 7230 0 -1 270
box -12 -8 32 272
use FILL  FILL_7__1810_
timestamp 1701859473
transform -1 0 7210 0 1 1310
box -12 -8 32 272
use FILL  FILL_7__1811_
timestamp 1701859473
transform 1 0 7550 0 -1 1830
box -12 -8 32 272
use FILL  FILL_7__1812_
timestamp 1701859473
transform -1 0 7630 0 -1 1310
box -12 -8 32 272
use FILL  FILL_7__1814_
timestamp 1701859473
transform -1 0 8250 0 -1 1830
box -12 -8 32 272
use FILL  FILL_7__1815_
timestamp 1701859473
transform 1 0 8450 0 1 2350
box -12 -8 32 272
use FILL  FILL_7__1816_
timestamp 1701859473
transform -1 0 9730 0 -1 2350
box -12 -8 32 272
use FILL  FILL_7__1817_
timestamp 1701859473
transform -1 0 9450 0 1 1310
box -12 -8 32 272
use FILL  FILL_7__1818_
timestamp 1701859473
transform -1 0 9650 0 1 270
box -12 -8 32 272
use FILL  FILL_7__1819_
timestamp 1701859473
transform -1 0 8470 0 -1 1830
box -12 -8 32 272
use FILL  FILL_7__1820_
timestamp 1701859473
transform -1 0 8550 0 1 1310
box -12 -8 32 272
use FILL  FILL_7__1822_
timestamp 1701859473
transform -1 0 4790 0 -1 790
box -12 -8 32 272
use FILL  FILL_7__1823_
timestamp 1701859473
transform -1 0 4330 0 -1 790
box -12 -8 32 272
use FILL  FILL_7__1824_
timestamp 1701859473
transform 1 0 4710 0 1 2350
box -12 -8 32 272
use FILL  FILL_7__1825_
timestamp 1701859473
transform 1 0 5770 0 1 1830
box -12 -8 32 272
use FILL  FILL_7__1826_
timestamp 1701859473
transform 1 0 8270 0 -1 270
box -12 -8 32 272
use FILL  FILL_7__1827_
timestamp 1701859473
transform 1 0 9410 0 -1 790
box -12 -8 32 272
use FILL  FILL_7__1829_
timestamp 1701859473
transform 1 0 5870 0 1 270
box -12 -8 32 272
use FILL  FILL_7__1830_
timestamp 1701859473
transform 1 0 3310 0 1 4430
box -12 -8 32 272
use FILL  FILL_7__1831_
timestamp 1701859473
transform -1 0 8090 0 -1 790
box -12 -8 32 272
use FILL  FILL_7__1832_
timestamp 1701859473
transform 1 0 6590 0 -1 790
box -12 -8 32 272
use FILL  FILL_7__1833_
timestamp 1701859473
transform -1 0 790 0 1 270
box -12 -8 32 272
use FILL  FILL_7__1834_
timestamp 1701859473
transform 1 0 1230 0 -1 1310
box -12 -8 32 272
use FILL  FILL_7__1836_
timestamp 1701859473
transform 1 0 1170 0 1 790
box -12 -8 32 272
use FILL  FILL_7__1837_
timestamp 1701859473
transform -1 0 2570 0 1 790
box -12 -8 32 272
use FILL  FILL_7__1838_
timestamp 1701859473
transform 1 0 2310 0 1 790
box -12 -8 32 272
use FILL  FILL_7__1839_
timestamp 1701859473
transform -1 0 370 0 1 270
box -12 -8 32 272
use FILL  FILL_7__1840_
timestamp 1701859473
transform -1 0 1010 0 1 2870
box -12 -8 32 272
use FILL  FILL_7__1841_
timestamp 1701859473
transform 1 0 3790 0 1 2870
box -12 -8 32 272
use FILL  FILL_7__1843_
timestamp 1701859473
transform -1 0 4010 0 -1 2350
box -12 -8 32 272
use FILL  FILL_7__1844_
timestamp 1701859473
transform 1 0 3910 0 -1 2870
box -12 -8 32 272
use FILL  FILL_7__1845_
timestamp 1701859473
transform -1 0 1850 0 -1 4950
box -12 -8 32 272
use FILL  FILL_7__1846_
timestamp 1701859473
transform 1 0 4210 0 1 4430
box -12 -8 32 272
use FILL  FILL_7__1847_
timestamp 1701859473
transform 1 0 3530 0 1 4430
box -12 -8 32 272
use FILL  FILL_7__1848_
timestamp 1701859473
transform 1 0 3970 0 1 4430
box -12 -8 32 272
use FILL  FILL_7__1849_
timestamp 1701859473
transform -1 0 4170 0 -1 2870
box -12 -8 32 272
use FILL  FILL_7__1851_
timestamp 1701859473
transform 1 0 1650 0 -1 1830
box -12 -8 32 272
use FILL  FILL_7__1852_
timestamp 1701859473
transform -1 0 2470 0 1 2350
box -12 -8 32 272
use FILL  FILL_7__1853_
timestamp 1701859473
transform 1 0 150 0 -1 2350
box -12 -8 32 272
use FILL  FILL_7__1854_
timestamp 1701859473
transform 1 0 2390 0 -1 2350
box -12 -8 32 272
use FILL  FILL_7__1855_
timestamp 1701859473
transform -1 0 2650 0 -1 2350
box -12 -8 32 272
use FILL  FILL_7__1856_
timestamp 1701859473
transform 1 0 1550 0 -1 790
box -12 -8 32 272
use FILL  FILL_7__1858_
timestamp 1701859473
transform 1 0 2490 0 -1 790
box -12 -8 32 272
use FILL  FILL_7__1859_
timestamp 1701859473
transform 1 0 2270 0 -1 790
box -12 -8 32 272
use FILL  FILL_7__1860_
timestamp 1701859473
transform -1 0 1810 0 -1 790
box -12 -8 32 272
use FILL  FILL_7__1861_
timestamp 1701859473
transform -1 0 2050 0 -1 790
box -12 -8 32 272
use FILL  FILL_7__1862_
timestamp 1701859473
transform -1 0 2130 0 1 270
box -12 -8 32 272
use FILL  FILL_7__1863_
timestamp 1701859473
transform 1 0 2350 0 1 270
box -12 -8 32 272
use FILL  FILL_7__1865_
timestamp 1701859473
transform 1 0 7390 0 -1 1310
box -12 -8 32 272
use FILL  FILL_7__1866_
timestamp 1701859473
transform 1 0 3750 0 -1 1310
box -12 -8 32 272
use FILL  FILL_7__1867_
timestamp 1701859473
transform 1 0 1210 0 -1 1830
box -12 -8 32 272
use FILL  FILL_7__1868_
timestamp 1701859473
transform 1 0 1650 0 1 1310
box -12 -8 32 272
use FILL  FILL_7__1869_
timestamp 1701859473
transform 1 0 2070 0 1 1310
box -12 -8 32 272
use FILL  FILL_7__1870_
timestamp 1701859473
transform -1 0 1690 0 -1 1310
box -12 -8 32 272
use FILL  FILL_7__1871_
timestamp 1701859473
transform -1 0 2810 0 -1 1310
box -12 -8 32 272
use FILL  FILL_7__1873_
timestamp 1701859473
transform 1 0 770 0 1 790
box -12 -8 32 272
use FILL  FILL_7__1874_
timestamp 1701859473
transform -1 0 1410 0 1 790
box -12 -8 32 272
use FILL  FILL_7__1875_
timestamp 1701859473
transform 1 0 990 0 -1 790
box -12 -8 32 272
use FILL  FILL_7__1876_
timestamp 1701859473
transform 1 0 1310 0 -1 790
box -12 -8 32 272
use FILL  FILL_7__1877_
timestamp 1701859473
transform 1 0 2250 0 1 4950
box -12 -8 32 272
use FILL  FILL_7__1878_
timestamp 1701859473
transform 1 0 590 0 -1 1310
box -12 -8 32 272
use FILL  FILL_7__1880_
timestamp 1701859473
transform -1 0 2070 0 -1 4950
box -12 -8 32 272
use FILL  FILL_7__1881_
timestamp 1701859473
transform -1 0 2310 0 -1 4950
box -12 -8 32 272
use FILL  FILL_7__1882_
timestamp 1701859473
transform 1 0 1630 0 -1 3390
box -12 -8 32 272
use FILL  FILL_7__1883_
timestamp 1701859473
transform 1 0 1110 0 -1 3390
box -12 -8 32 272
use FILL  FILL_7__1884_
timestamp 1701859473
transform -1 0 4130 0 1 3390
box -12 -8 32 272
use FILL  FILL_7__1885_
timestamp 1701859473
transform -1 0 3850 0 -1 3390
box -12 -8 32 272
use FILL  FILL_7__1887_
timestamp 1701859473
transform -1 0 3570 0 1 2870
box -12 -8 32 272
use FILL  FILL_7__1888_
timestamp 1701859473
transform -1 0 2610 0 1 270
box -12 -8 32 272
use FILL  FILL_7__1889_
timestamp 1701859473
transform 1 0 1750 0 -1 2870
box -12 -8 32 272
use FILL  FILL_7__1890_
timestamp 1701859473
transform -1 0 390 0 -1 1830
box -12 -8 32 272
use FILL  FILL_7__1891_
timestamp 1701859473
transform 1 0 150 0 -1 1830
box -12 -8 32 272
use FILL  FILL_7__1892_
timestamp 1701859473
transform 1 0 4990 0 -1 3390
box -12 -8 32 272
use FILL  FILL_7__1894_
timestamp 1701859473
transform 1 0 4190 0 1 1830
box -12 -8 32 272
use FILL  FILL_7__1895_
timestamp 1701859473
transform -1 0 1930 0 1 1830
box -12 -8 32 272
use FILL  FILL_7__1896_
timestamp 1701859473
transform 1 0 1950 0 -1 2350
box -12 -8 32 272
use FILL  FILL_7__1897_
timestamp 1701859473
transform 1 0 3570 0 1 2350
box -12 -8 32 272
use FILL  FILL_7__1898_
timestamp 1701859473
transform 1 0 3350 0 1 2350
box -12 -8 32 272
use FILL  FILL_7__1899_
timestamp 1701859473
transform -1 0 3330 0 -1 2350
box -12 -8 32 272
use FILL  FILL_7__1900_
timestamp 1701859473
transform -1 0 4170 0 -1 1830
box -12 -8 32 272
use FILL  FILL_7__1902_
timestamp 1701859473
transform 1 0 5110 0 1 1830
box -12 -8 32 272
use FILL  FILL_7__1903_
timestamp 1701859473
transform 1 0 3430 0 1 1310
box -12 -8 32 272
use FILL  FILL_7__1904_
timestamp 1701859473
transform -1 0 3530 0 -1 1310
box -12 -8 32 272
use FILL  FILL_7__1905_
timestamp 1701859473
transform 1 0 3070 0 1 270
box -12 -8 32 272
use FILL  FILL_7__1906_
timestamp 1701859473
transform 1 0 350 0 1 2350
box -12 -8 32 272
use FILL  FILL_7__1907_
timestamp 1701859473
transform -1 0 3110 0 -1 2350
box -12 -8 32 272
use FILL  FILL_7__1909_
timestamp 1701859473
transform -1 0 6130 0 -1 2350
box -12 -8 32 272
use FILL  FILL_7__1910_
timestamp 1701859473
transform -1 0 5630 0 -1 2350
box -12 -8 32 272
use FILL  FILL_7__1911_
timestamp 1701859473
transform -1 0 790 0 1 2870
box -12 -8 32 272
use FILL  FILL_7__1912_
timestamp 1701859473
transform -1 0 3390 0 1 3910
box -12 -8 32 272
use FILL  FILL_7__1913_
timestamp 1701859473
transform -1 0 1110 0 -1 2870
box -12 -8 32 272
use FILL  FILL_7__1914_
timestamp 1701859473
transform -1 0 1550 0 1 3390
box -12 -8 32 272
use FILL  FILL_7__1916_
timestamp 1701859473
transform -1 0 3490 0 1 3390
box -12 -8 32 272
use FILL  FILL_7__1917_
timestamp 1701859473
transform -1 0 4770 0 -1 3390
box -12 -8 32 272
use FILL  FILL_7__1918_
timestamp 1701859473
transform 1 0 1810 0 1 4950
box -12 -8 32 272
use FILL  FILL_7__1919_
timestamp 1701859473
transform -1 0 1330 0 -1 2870
box -12 -8 32 272
use FILL  FILL_7__1920_
timestamp 1701859473
transform -1 0 5110 0 1 4430
box -12 -8 32 272
use FILL  FILL_7__1921_
timestamp 1701859473
transform 1 0 4870 0 1 4430
box -12 -8 32 272
use FILL  FILL_7__1923_
timestamp 1701859473
transform 1 0 4530 0 -1 3390
box -12 -8 32 272
use FILL  FILL_7__1924_
timestamp 1701859473
transform 1 0 2030 0 1 4950
box -12 -8 32 272
use FILL  FILL_7__1925_
timestamp 1701859473
transform 1 0 6170 0 -1 4430
box -12 -8 32 272
use FILL  FILL_7__1926_
timestamp 1701859473
transform 1 0 790 0 -1 1310
box -12 -8 32 272
use FILL  FILL_7__1927_
timestamp 1701859473
transform 1 0 3030 0 -1 1310
box -12 -8 32 272
use FILL  FILL_7__1928_
timestamp 1701859473
transform -1 0 3290 0 -1 1310
box -12 -8 32 272
use FILL  FILL_7__1929_
timestamp 1701859473
transform 1 0 3470 0 1 790
box -12 -8 32 272
use FILL  FILL_7__1931_
timestamp 1701859473
transform 1 0 3890 0 1 270
box -12 -8 32 272
use FILL  FILL_7__1932_
timestamp 1701859473
transform -1 0 4130 0 1 270
box -12 -8 32 272
use FILL  FILL_7__1933_
timestamp 1701859473
transform -1 0 1930 0 1 270
box -12 -8 32 272
use FILL  FILL_7__1934_
timestamp 1701859473
transform -1 0 5550 0 1 790
box -12 -8 32 272
use FILL  FILL_7__1935_
timestamp 1701859473
transform 1 0 5670 0 -1 270
box -12 -8 32 272
use FILL  FILL_7__1936_
timestamp 1701859473
transform -1 0 8430 0 1 3390
box -12 -8 32 272
use FILL  FILL_7__1938_
timestamp 1701859473
transform -1 0 7850 0 -1 270
box -12 -8 32 272
use FILL  FILL_7__1939_
timestamp 1701859473
transform -1 0 6770 0 -1 270
box -12 -8 32 272
use FILL  FILL_7__1940_
timestamp 1701859473
transform -1 0 5890 0 -1 270
box -12 -8 32 272
use FILL  FILL_7__1941_
timestamp 1701859473
transform 1 0 5910 0 -1 790
box -12 -8 32 272
use FILL  FILL_7__1942_
timestamp 1701859473
transform 1 0 4890 0 -1 1310
box -12 -8 32 272
use FILL  FILL_7__1943_
timestamp 1701859473
transform 1 0 8150 0 1 270
box -12 -8 32 272
use FILL  FILL_7__1945_
timestamp 1701859473
transform 1 0 7930 0 1 270
box -12 -8 32 272
use FILL  FILL_7__1946_
timestamp 1701859473
transform -1 0 6130 0 1 270
box -12 -8 32 272
use FILL  FILL_7__1947_
timestamp 1701859473
transform -1 0 6150 0 -1 790
box -12 -8 32 272
use FILL  FILL_7__1948_
timestamp 1701859473
transform 1 0 5430 0 -1 790
box -12 -8 32 272
use FILL  FILL_7__1949_
timestamp 1701859473
transform 1 0 4670 0 -1 1310
box -12 -8 32 272
use FILL  FILL_7__1950_
timestamp 1701859473
transform -1 0 8310 0 -1 790
box -12 -8 32 272
use FILL  FILL_7__1951_
timestamp 1701859473
transform 1 0 590 0 -1 2350
box -12 -8 32 272
use FILL  FILL_7__1953_
timestamp 1701859473
transform 1 0 5870 0 -1 2350
box -12 -8 32 272
use FILL  FILL_7__1954_
timestamp 1701859473
transform 1 0 8250 0 -1 1310
box -12 -8 32 272
use FILL  FILL_7__1955_
timestamp 1701859473
transform -1 0 8790 0 1 1310
box -12 -8 32 272
use FILL  FILL_7__1956_
timestamp 1701859473
transform -1 0 6330 0 -1 1310
box -12 -8 32 272
use FILL  FILL_7__1957_
timestamp 1701859473
transform -1 0 6090 0 -1 1310
box -12 -8 32 272
use FILL  FILL_7__1958_
timestamp 1701859473
transform 1 0 5350 0 -1 1310
box -12 -8 32 272
use FILL  FILL_7__1960_
timestamp 1701859473
transform -1 0 6230 0 -1 2870
box -12 -8 32 272
use FILL  FILL_7__1961_
timestamp 1701859473
transform -1 0 4490 0 1 2350
box -12 -8 32 272
use FILL  FILL_7__1962_
timestamp 1701859473
transform 1 0 5950 0 1 2350
box -12 -8 32 272
use FILL  FILL_7__1963_
timestamp 1701859473
transform 1 0 5410 0 1 1310
box -12 -8 32 272
use FILL  FILL_7__1964_
timestamp 1701859473
transform 1 0 9230 0 1 1310
box -12 -8 32 272
use FILL  FILL_7__1965_
timestamp 1701859473
transform 1 0 7630 0 1 790
box -12 -8 32 272
use FILL  FILL_7__1967_
timestamp 1701859473
transform -1 0 6810 0 1 270
box -12 -8 32 272
use FILL  FILL_7__1968_
timestamp 1701859473
transform 1 0 5590 0 -1 1310
box -12 -8 32 272
use FILL  FILL_7__1969_
timestamp 1701859473
transform 1 0 5790 0 1 2870
box -12 -8 32 272
use FILL  FILL_7__1970_
timestamp 1701859473
transform 1 0 5430 0 -1 3390
box -12 -8 32 272
use FILL  FILL_7__1971_
timestamp 1701859473
transform 1 0 5870 0 1 3910
box -12 -8 32 272
use FILL  FILL_7__1972_
timestamp 1701859473
transform 1 0 5810 0 1 4950
box -12 -8 32 272
use FILL  FILL_7__1974_
timestamp 1701859473
transform 1 0 6330 0 -1 3910
box -12 -8 32 272
use FILL  FILL_7__1975_
timestamp 1701859473
transform -1 0 6130 0 1 3910
box -12 -8 32 272
use FILL  FILL_7__1976_
timestamp 1701859473
transform -1 0 6590 0 -1 3910
box -12 -8 32 272
use FILL  FILL_7__1977_
timestamp 1701859473
transform 1 0 6910 0 1 2870
box -12 -8 32 272
use FILL  FILL_7__1978_
timestamp 1701859473
transform -1 0 6450 0 -1 2870
box -12 -8 32 272
use FILL  FILL_7__1979_
timestamp 1701859473
transform 1 0 6490 0 1 2870
box -12 -8 32 272
use FILL  FILL_7__1980_
timestamp 1701859473
transform 1 0 6690 0 1 2870
box -12 -8 32 272
use FILL  FILL_7__1982_
timestamp 1701859473
transform -1 0 5730 0 -1 1830
box -12 -8 32 272
use FILL  FILL_7__1983_
timestamp 1701859473
transform -1 0 4830 0 -1 270
box -12 -8 32 272
use FILL  FILL_7__1984_
timestamp 1701859473
transform -1 0 6530 0 -1 1310
box -12 -8 32 272
use FILL  FILL_7__1985_
timestamp 1701859473
transform 1 0 5090 0 -1 1310
box -12 -8 32 272
use FILL  FILL_7__1986_
timestamp 1701859473
transform 1 0 8290 0 1 790
box -12 -8 32 272
use FILL  FILL_7__1987_
timestamp 1701859473
transform 1 0 6970 0 1 1310
box -12 -8 32 272
use FILL  FILL_7__1989_
timestamp 1701859473
transform 1 0 2790 0 -1 5470
box -12 -8 32 272
use FILL  FILL_7__1990_
timestamp 1701859473
transform 1 0 2110 0 1 1830
box -12 -8 32 272
use FILL  FILL_7__1991_
timestamp 1701859473
transform -1 0 2830 0 1 1830
box -12 -8 32 272
use FILL  FILL_7__1992_
timestamp 1701859473
transform -1 0 4230 0 -1 2350
box -12 -8 32 272
use FILL  FILL_7__1993_
timestamp 1701859473
transform -1 0 4470 0 -1 2350
box -12 -8 32 272
use FILL  FILL_7__1994_
timestamp 1701859473
transform 1 0 2570 0 1 1830
box -12 -8 32 272
use FILL  FILL_7__1996_
timestamp 1701859473
transform -1 0 6730 0 1 790
box -12 -8 32 272
use FILL  FILL_7__1997_
timestamp 1701859473
transform -1 0 5070 0 1 790
box -12 -8 32 272
use FILL  FILL_7__1998_
timestamp 1701859473
transform 1 0 4330 0 1 270
box -12 -8 32 272
use FILL  FILL_7__1999_
timestamp 1701859473
transform -1 0 3930 0 -1 270
box -12 -8 32 272
use FILL  FILL_7__2000_
timestamp 1701859473
transform -1 0 4610 0 -1 270
box -12 -8 32 272
use FILL  FILL_7__2001_
timestamp 1701859473
transform -1 0 5990 0 -1 2870
box -12 -8 32 272
use FILL  FILL_7__2002_
timestamp 1701859473
transform -1 0 1930 0 1 2870
box -12 -8 32 272
use FILL  FILL_7__2004_
timestamp 1701859473
transform 1 0 2850 0 -1 3390
box -12 -8 32 272
use FILL  FILL_7__2005_
timestamp 1701859473
transform -1 0 3130 0 1 2870
box -12 -8 32 272
use FILL  FILL_7__2006_
timestamp 1701859473
transform 1 0 2870 0 1 2870
box -12 -8 32 272
use FILL  FILL_7__2007_
timestamp 1701859473
transform 1 0 6890 0 -1 2870
box -12 -8 32 272
use FILL  FILL_7__2008_
timestamp 1701859473
transform 1 0 570 0 -1 1830
box -12 -8 32 272
use FILL  FILL_7__2009_
timestamp 1701859473
transform -1 0 4090 0 -1 3390
box -12 -8 32 272
use FILL  FILL_7__2011_
timestamp 1701859473
transform -1 0 2130 0 1 790
box -12 -8 32 272
use FILL  FILL_7__2012_
timestamp 1701859473
transform 1 0 1630 0 1 790
box -12 -8 32 272
use FILL  FILL_7__2013_
timestamp 1701859473
transform -1 0 1890 0 1 790
box -12 -8 32 272
use FILL  FILL_7__2014_
timestamp 1701859473
transform 1 0 4550 0 1 1310
box -12 -8 32 272
use FILL  FILL_7__2015_
timestamp 1701859473
transform 1 0 3270 0 1 1830
box -12 -8 32 272
use FILL  FILL_7__2016_
timestamp 1701859473
transform -1 0 3770 0 1 1830
box -12 -8 32 272
use FILL  FILL_7__2018_
timestamp 1701859473
transform 1 0 5050 0 -1 1830
box -12 -8 32 272
use FILL  FILL_7__2019_
timestamp 1701859473
transform -1 0 5570 0 -1 2870
box -12 -8 32 272
use FILL  FILL_7__2020_
timestamp 1701859473
transform -1 0 5330 0 -1 2870
box -12 -8 32 272
use FILL  FILL_7__2021_
timestamp 1701859473
transform -1 0 6970 0 -1 1310
box -12 -8 32 272
use FILL  FILL_7__2022_
timestamp 1701859473
transform -1 0 7210 0 1 790
box -12 -8 32 272
use FILL  FILL_7__2023_
timestamp 1701859473
transform 1 0 8250 0 1 1830
box -12 -8 32 272
use FILL  FILL_7__2025_
timestamp 1701859473
transform 1 0 9630 0 -1 790
box -12 -8 32 272
use FILL  FILL_7__2026_
timestamp 1701859473
transform -1 0 8770 0 1 790
box -12 -8 32 272
use FILL  FILL_7__2027_
timestamp 1701859473
transform -1 0 6970 0 1 790
box -12 -8 32 272
use FILL  FILL_7__2028_
timestamp 1701859473
transform 1 0 7070 0 -1 790
box -12 -8 32 272
use FILL  FILL_7__2029_
timestamp 1701859473
transform 1 0 7510 0 1 270
box -12 -8 32 272
use FILL  FILL_7__2030_
timestamp 1701859473
transform -1 0 7190 0 -1 1310
box -12 -8 32 272
use FILL  FILL_7__2031_
timestamp 1701859473
transform 1 0 7510 0 -1 790
box -12 -8 32 272
use FILL  FILL_7__2033_
timestamp 1701859473
transform 1 0 8290 0 1 1310
box -12 -8 32 272
use FILL  FILL_7__2034_
timestamp 1701859473
transform -1 0 8970 0 -1 1310
box -12 -8 32 272
use FILL  FILL_7__2035_
timestamp 1701859473
transform -1 0 8550 0 1 790
box -12 -8 32 272
use FILL  FILL_7__2036_
timestamp 1701859473
transform -1 0 8710 0 -1 1830
box -12 -8 32 272
use FILL  FILL_7__2037_
timestamp 1701859473
transform -1 0 8770 0 -1 790
box -12 -8 32 272
use FILL  FILL_7__2038_
timestamp 1701859473
transform 1 0 8070 0 1 790
box -12 -8 32 272
use FILL  FILL_7__2040_
timestamp 1701859473
transform -1 0 7770 0 -1 790
box -12 -8 32 272
use FILL  FILL_7__2041_
timestamp 1701859473
transform -1 0 6990 0 -1 270
box -12 -8 32 272
use FILL  FILL_7__2042_
timestamp 1701859473
transform 1 0 8970 0 -1 790
box -12 -8 32 272
use FILL  FILL_7__2043_
timestamp 1701859473
transform 1 0 7290 0 1 270
box -12 -8 32 272
use FILL  FILL_7__2044_
timestamp 1701859473
transform 1 0 7030 0 1 270
box -12 -8 32 272
use FILL  FILL_7__2045_
timestamp 1701859473
transform -1 0 6350 0 1 270
box -12 -8 32 272
use FILL  FILL_7__2047_
timestamp 1701859473
transform -1 0 6310 0 -1 270
box -12 -8 32 272
use FILL  FILL_7__2048_
timestamp 1701859473
transform -1 0 6110 0 -1 270
box -12 -8 32 272
use FILL  FILL_7__2049_
timestamp 1701859473
transform -1 0 7290 0 -1 790
box -12 -8 32 272
use FILL  FILL_7__2050_
timestamp 1701859473
transform 1 0 1530 0 -1 2870
box -12 -8 32 272
use FILL  FILL_7__2051_
timestamp 1701859473
transform 1 0 6330 0 -1 2350
box -12 -8 32 272
use FILL  FILL_7__2052_
timestamp 1701859473
transform -1 0 6230 0 1 790
box -12 -8 32 272
use FILL  FILL_7__2054_
timestamp 1701859473
transform 1 0 2950 0 1 1310
box -12 -8 32 272
use FILL  FILL_7__2055_
timestamp 1701859473
transform -1 0 3210 0 1 1310
box -12 -8 32 272
use FILL  FILL_7__2056_
timestamp 1701859473
transform -1 0 1930 0 -1 1310
box -12 -8 32 272
use FILL  FILL_7__2057_
timestamp 1701859473
transform 1 0 2790 0 1 790
box -12 -8 32 272
use FILL  FILL_7__2058_
timestamp 1701859473
transform 1 0 3710 0 1 790
box -12 -8 32 272
use FILL  FILL_7__2059_
timestamp 1701859473
transform 1 0 3950 0 1 790
box -12 -8 32 272
use FILL  FILL_7__2060_
timestamp 1701859473
transform -1 0 4190 0 1 790
box -12 -8 32 272
use FILL  FILL_7__2062_
timestamp 1701859473
transform 1 0 2830 0 1 270
box -12 -8 32 272
use FILL  FILL_7__2063_
timestamp 1701859473
transform 1 0 3210 0 -1 270
box -12 -8 32 272
use FILL  FILL_7__2064_
timestamp 1701859473
transform 1 0 3450 0 -1 270
box -12 -8 32 272
use FILL  FILL_7__2065_
timestamp 1701859473
transform -1 0 3690 0 -1 270
box -12 -8 32 272
use FILL  FILL_7__2066_
timestamp 1701859473
transform -1 0 5470 0 -1 270
box -12 -8 32 272
use FILL  FILL_7__2067_
timestamp 1701859473
transform 1 0 7410 0 1 790
box -12 -8 32 272
use FILL  FILL_7__2069_
timestamp 1701859473
transform 1 0 3450 0 -1 1830
box -12 -8 32 272
use FILL  FILL_7__2070_
timestamp 1701859473
transform -1 0 3930 0 -1 1830
box -12 -8 32 272
use FILL  FILL_7__2071_
timestamp 1701859473
transform -1 0 5770 0 1 790
box -12 -8 32 272
use FILL  FILL_7__2072_
timestamp 1701859473
transform -1 0 7830 0 1 1310
box -12 -8 32 272
use FILL  FILL_7__2073_
timestamp 1701859473
transform 1 0 6710 0 1 1310
box -12 -8 32 272
use FILL  FILL_7__2074_
timestamp 1701859473
transform 1 0 1850 0 1 1310
box -12 -8 32 272
use FILL  FILL_7__2076_
timestamp 1701859473
transform -1 0 2370 0 -1 1310
box -12 -8 32 272
use FILL  FILL_7__2077_
timestamp 1701859473
transform 1 0 4230 0 -1 1310
box -12 -8 32 272
use FILL  FILL_7__2078_
timestamp 1701859473
transform -1 0 2370 0 1 1830
box -12 -8 32 272
use FILL  FILL_7__2079_
timestamp 1701859473
transform -1 0 1010 0 -1 1830
box -12 -8 32 272
use FILL  FILL_7__2080_
timestamp 1701859473
transform 1 0 2330 0 -1 1830
box -12 -8 32 272
use FILL  FILL_7__2081_
timestamp 1701859473
transform 1 0 2570 0 -1 1830
box -12 -8 32 272
use FILL  FILL_7__2082_
timestamp 1701859473
transform -1 0 2790 0 -1 1830
box -12 -8 32 272
use FILL  FILL_7__2084_
timestamp 1701859473
transform -1 0 5310 0 1 790
box -12 -8 32 272
use FILL  FILL_7__2085_
timestamp 1701859473
transform -1 0 5150 0 -1 270
box -12 -8 32 272
use FILL  FILL_7__2086_
timestamp 1701859473
transform -1 0 4370 0 -1 270
box -12 -8 32 272
use FILL  FILL_7__2087_
timestamp 1701859473
transform -1 0 4850 0 1 790
box -12 -8 32 272
use FILL  FILL_7__2088_
timestamp 1701859473
transform -1 0 5690 0 1 270
box -12 -8 32 272
use FILL  FILL_7__2089_
timestamp 1701859473
transform 1 0 5450 0 1 270
box -12 -8 32 272
use FILL  FILL_7__2091_
timestamp 1701859473
transform 1 0 3250 0 1 790
box -12 -8 32 272
use FILL  FILL_7__2092_
timestamp 1701859473
transform 1 0 2810 0 -1 270
box -12 -8 32 272
use FILL  FILL_7__2093_
timestamp 1701859473
transform -1 0 2970 0 -1 790
box -12 -8 32 272
use FILL  FILL_7__2094_
timestamp 1701859473
transform 1 0 2370 0 -1 270
box -12 -8 32 272
use FILL  FILL_7__2095_
timestamp 1701859473
transform 1 0 2570 0 -1 270
box -12 -8 32 272
use FILL  FILL_7__2096_
timestamp 1701859473
transform -1 0 5030 0 1 270
box -12 -8 32 272
use FILL  FILL_7__2098_
timestamp 1701859473
transform 1 0 4790 0 1 270
box -12 -8 32 272
use FILL  FILL_7__2099_
timestamp 1701859473
transform 1 0 4110 0 -1 270
box -12 -8 32 272
use FILL  FILL_7__2100_
timestamp 1701859473
transform -1 0 5970 0 -1 1830
box -12 -8 32 272
use FILL  FILL_7__2101_
timestamp 1701859473
transform -1 0 5890 0 1 1310
box -12 -8 32 272
use FILL  FILL_7__2102_
timestamp 1701859473
transform -1 0 6290 0 1 1310
box -12 -8 32 272
use FILL  FILL_7__2103_
timestamp 1701859473
transform 1 0 5850 0 -1 1310
box -12 -8 32 272
use FILL  FILL_7__2105_
timestamp 1701859473
transform -1 0 4390 0 -1 1830
box -12 -8 32 272
use FILL  FILL_7__2106_
timestamp 1701859473
transform 1 0 4070 0 -1 790
box -12 -8 32 272
use FILL  FILL_7__2107_
timestamp 1701859473
transform -1 0 3650 0 -1 790
box -12 -8 32 272
use FILL  FILL_7__2108_
timestamp 1701859473
transform 1 0 3010 0 1 790
box -12 -8 32 272
use FILL  FILL_7__2109_
timestamp 1701859473
transform -1 0 3430 0 -1 790
box -12 -8 32 272
use FILL  FILL_7__2110_
timestamp 1701859473
transform 1 0 3190 0 -1 790
box -12 -8 32 272
use FILL  FILL_7__2111_
timestamp 1701859473
transform -1 0 3870 0 -1 790
box -12 -8 32 272
use FILL  FILL_7__2113_
timestamp 1701859473
transform -1 0 5210 0 1 1310
box -12 -8 32 272
use FILL  FILL_7__2114_
timestamp 1701859473
transform -1 0 5650 0 1 1310
box -12 -8 32 272
use FILL  FILL_7__2115_
timestamp 1701859473
transform -1 0 5690 0 -1 790
box -12 -8 32 272
use FILL  FILL_7__2116_
timestamp 1701859473
transform 1 0 2510 0 1 1310
box -12 -8 32 272
use FILL  FILL_7__2117_
timestamp 1701859473
transform 1 0 2710 0 1 1310
box -12 -8 32 272
use FILL  FILL_7__2118_
timestamp 1701859473
transform 1 0 3890 0 1 1310
box -12 -8 32 272
use FILL  FILL_7__2120_
timestamp 1701859473
transform 1 0 4010 0 -1 1310
box -12 -8 32 272
use FILL  FILL_7__2121_
timestamp 1701859473
transform -1 0 4590 0 1 270
box -12 -8 32 272
use FILL  FILL_7__2122_
timestamp 1701859473
transform -1 0 2930 0 1 2350
box -12 -8 32 272
use FILL  FILL_7__2123_
timestamp 1701859473
transform 1 0 2870 0 -1 2350
box -12 -8 32 272
use FILL  FILL_7__2124_
timestamp 1701859473
transform -1 0 3770 0 -1 2350
box -12 -8 32 272
use FILL  FILL_7__2125_
timestamp 1701859473
transform 1 0 5890 0 -1 3390
box -12 -8 32 272
use FILL  FILL_7__2127_
timestamp 1701859473
transform -1 0 6050 0 1 2870
box -12 -8 32 272
use FILL  FILL_7__2128_
timestamp 1701859473
transform 1 0 4670 0 1 2870
box -12 -8 32 272
use FILL  FILL_7__2129_
timestamp 1701859473
transform 1 0 5350 0 1 2870
box -12 -8 32 272
use FILL  FILL_7__2130_
timestamp 1701859473
transform -1 0 4710 0 -1 2350
box -12 -8 32 272
use FILL  FILL_7__2131_
timestamp 1701859473
transform 1 0 4750 0 1 1310
box -12 -8 32 272
use FILL  FILL_7__2132_
timestamp 1701859473
transform -1 0 4630 0 1 790
box -12 -8 32 272
use FILL  FILL_7__2134_
timestamp 1701859473
transform 1 0 3670 0 -1 2870
box -12 -8 32 272
use FILL  FILL_7__2135_
timestamp 1701859473
transform 1 0 4290 0 -1 3390
box -12 -8 32 272
use FILL  FILL_7__2136_
timestamp 1701859473
transform -1 0 2830 0 1 3390
box -12 -8 32 272
use FILL  FILL_7__2137_
timestamp 1701859473
transform 1 0 2390 0 1 3390
box -12 -8 32 272
use FILL  FILL_7__2138_
timestamp 1701859473
transform 1 0 3190 0 -1 4430
box -12 -8 32 272
use FILL  FILL_7__2139_
timestamp 1701859473
transform -1 0 2970 0 -1 4430
box -12 -8 32 272
use FILL  FILL_7__2140_
timestamp 1701859473
transform 1 0 2890 0 1 4430
box -12 -8 32 272
use FILL  FILL_7__2142_
timestamp 1701859473
transform 1 0 3010 0 1 3390
box -12 -8 32 272
use FILL  FILL_7__2143_
timestamp 1701859473
transform -1 0 7510 0 -1 3390
box -12 -8 32 272
use FILL  FILL_7__2144_
timestamp 1701859473
transform 1 0 2150 0 1 2870
box -12 -8 32 272
use FILL  FILL_7__2145_
timestamp 1701859473
transform -1 0 10130 0 -1 2870
box -12 -8 32 272
use FILL  FILL_7__2146_
timestamp 1701859473
transform -1 0 7710 0 -1 3390
box -12 -8 32 272
use FILL  FILL_7__2147_
timestamp 1701859473
transform 1 0 7670 0 -1 3910
box -12 -8 32 272
use FILL  FILL_7__2149_
timestamp 1701859473
transform 1 0 7710 0 1 3390
box -12 -8 32 272
use FILL  FILL_7__2150_
timestamp 1701859473
transform -1 0 7970 0 1 3390
box -12 -8 32 272
use FILL  FILL_7__2151_
timestamp 1701859473
transform 1 0 7250 0 -1 3390
box -12 -8 32 272
use FILL  FILL_7__2152_
timestamp 1701859473
transform 1 0 7010 0 -1 3390
box -12 -8 32 272
use FILL  FILL_7__2153_
timestamp 1701859473
transform -1 0 6150 0 -1 3390
box -12 -8 32 272
use FILL  FILL_7__2154_
timestamp 1701859473
transform 1 0 2910 0 -1 7030
box -12 -8 32 272
use FILL  FILL_7__2156_
timestamp 1701859473
transform -1 0 4690 0 1 3910
box -12 -8 32 272
use FILL  FILL_7__2157_
timestamp 1701859473
transform -1 0 4830 0 -1 4430
box -12 -8 32 272
use FILL  FILL_7__2158_
timestamp 1701859473
transform -1 0 2690 0 1 2350
box -12 -8 32 272
use FILL  FILL_7__2159_
timestamp 1701859473
transform 1 0 3590 0 1 3910
box -12 -8 32 272
use FILL  FILL_7__2160_
timestamp 1701859473
transform -1 0 3910 0 -1 4430
box -12 -8 32 272
use FILL  FILL_7__2161_
timestamp 1701859473
transform -1 0 4050 0 1 3910
box -12 -8 32 272
use FILL  FILL_7__2162_
timestamp 1701859473
transform -1 0 4490 0 1 3910
box -12 -8 32 272
use FILL  FILL_7__2164_
timestamp 1701859473
transform -1 0 630 0 -1 4950
box -12 -8 32 272
use FILL  FILL_7__2165_
timestamp 1701859473
transform -1 0 3330 0 -1 3910
box -12 -8 32 272
use FILL  FILL_7__2166_
timestamp 1701859473
transform 1 0 4030 0 -1 3910
box -12 -8 32 272
use FILL  FILL_7__2167_
timestamp 1701859473
transform 1 0 4230 0 1 3910
box -12 -8 32 272
use FILL  FILL_7__2168_
timestamp 1701859473
transform 1 0 3150 0 1 3910
box -12 -8 32 272
use FILL  FILL_7__2169_
timestamp 1701859473
transform 1 0 2510 0 -1 4430
box -12 -8 32 272
use FILL  FILL_7__2171_
timestamp 1701859473
transform 1 0 4110 0 -1 4430
box -12 -8 32 272
use FILL  FILL_7__2172_
timestamp 1701859473
transform 1 0 4350 0 -1 4430
box -12 -8 32 272
use FILL  FILL_7__2173_
timestamp 1701859473
transform -1 0 4590 0 -1 4430
box -12 -8 32 272
use FILL  FILL_7__2174_
timestamp 1701859473
transform 1 0 6090 0 1 7030
box -12 -8 32 272
use FILL  FILL_7__2175_
timestamp 1701859473
transform -1 0 2590 0 1 8070
box -12 -8 32 272
use FILL  FILL_7__2176_
timestamp 1701859473
transform -1 0 6510 0 -1 8070
box -12 -8 32 272
use FILL  FILL_7__2178_
timestamp 1701859473
transform -1 0 4210 0 -1 8590
box -12 -8 32 272
use FILL  FILL_7__2179_
timestamp 1701859473
transform -1 0 6030 0 -1 8070
box -12 -8 32 272
use FILL  FILL_7__2180_
timestamp 1701859473
transform -1 0 3050 0 -1 9630
box -12 -8 32 272
use FILL  FILL_7__2181_
timestamp 1701859473
transform 1 0 5110 0 1 7550
box -12 -8 32 272
use FILL  FILL_7__2182_
timestamp 1701859473
transform 1 0 5630 0 -1 10150
box -12 -8 32 272
use FILL  FILL_7__2183_
timestamp 1701859473
transform -1 0 3610 0 1 10150
box -12 -8 32 272
use FILL  FILL_7__2185_
timestamp 1701859473
transform 1 0 6030 0 1 10150
box -12 -8 32 272
use FILL  FILL_7__2186_
timestamp 1701859473
transform 1 0 3590 0 1 10670
box -12 -8 32 272
use FILL  FILL_7__2187_
timestamp 1701859473
transform -1 0 5510 0 -1 10670
box -12 -8 32 272
use FILL  FILL_7__2188_
timestamp 1701859473
transform 1 0 2190 0 -1 10670
box -12 -8 32 272
use FILL  FILL_7__2189_
timestamp 1701859473
transform 1 0 5750 0 -1 10670
box -12 -8 32 272
use FILL  FILL_7__2190_
timestamp 1701859473
transform -1 0 2910 0 1 10150
box -12 -8 32 272
use FILL  FILL_7__2191_
timestamp 1701859473
transform -1 0 5390 0 -1 10150
box -12 -8 32 272
use FILL  FILL_7__2193_
timestamp 1701859473
transform 1 0 1310 0 -1 3910
box -12 -8 32 272
use FILL  FILL_7__2194_
timestamp 1701859473
transform 1 0 1110 0 -1 3910
box -12 -8 32 272
use FILL  FILL_7__2195_
timestamp 1701859473
transform 1 0 2690 0 1 3910
box -12 -8 32 272
use FILL  FILL_7__2196_
timestamp 1701859473
transform 1 0 2930 0 1 3910
box -12 -8 32 272
use FILL  FILL_7__2197_
timestamp 1701859473
transform 1 0 5410 0 1 3910
box -12 -8 32 272
use FILL  FILL_7__2198_
timestamp 1701859473
transform 1 0 350 0 1 1830
box -12 -8 32 272
use FILL  FILL_7__2200_
timestamp 1701859473
transform 1 0 5430 0 -1 3910
box -12 -8 32 272
use FILL  FILL_7__2201_
timestamp 1701859473
transform -1 0 5670 0 1 3910
box -12 -8 32 272
use FILL  FILL_7__2202_
timestamp 1701859473
transform -1 0 8250 0 -1 4430
box -12 -8 32 272
use FILL  FILL_7__2203_
timestamp 1701859473
transform -1 0 4970 0 -1 3910
box -12 -8 32 272
use FILL  FILL_7__2204_
timestamp 1701859473
transform 1 0 5190 0 -1 3910
box -12 -8 32 272
use FILL  FILL_7__2205_
timestamp 1701859473
transform -1 0 9050 0 -1 3910
box -12 -8 32 272
use FILL  FILL_7__2207_
timestamp 1701859473
transform 1 0 9590 0 -1 3910
box -12 -8 32 272
use FILL  FILL_7__2208_
timestamp 1701859473
transform -1 0 9850 0 -1 3910
box -12 -8 32 272
use FILL  FILL_7__2209_
timestamp 1701859473
transform -1 0 9650 0 1 4430
box -12 -8 32 272
use FILL  FILL_7__2210_
timestamp 1701859473
transform -1 0 10650 0 -1 4950
box -12 -8 32 272
use FILL  FILL_7__2211_
timestamp 1701859473
transform 1 0 9350 0 -1 3910
box -12 -8 32 272
use FILL  FILL_7__2212_
timestamp 1701859473
transform -1 0 8930 0 1 3910
box -12 -8 32 272
use FILL  FILL_7__2213_
timestamp 1701859473
transform -1 0 9370 0 1 3910
box -12 -8 32 272
use FILL  FILL_7__2215_
timestamp 1701859473
transform 1 0 9770 0 -1 4430
box -12 -8 32 272
use FILL  FILL_7__2216_
timestamp 1701859473
transform -1 0 9530 0 -1 7030
box -12 -8 32 272
use FILL  FILL_7__2217_
timestamp 1701859473
transform 1 0 9310 0 -1 4430
box -12 -8 32 272
use FILL  FILL_7__2218_
timestamp 1701859473
transform -1 0 9830 0 1 3910
box -12 -8 32 272
use FILL  FILL_7__2219_
timestamp 1701859473
transform 1 0 10010 0 1 3910
box -12 -8 32 272
use FILL  FILL_7__2220_
timestamp 1701859473
transform 1 0 10390 0 -1 4950
box -12 -8 32 272
use FILL  FILL_7__2222_
timestamp 1701859473
transform 1 0 10130 0 1 4430
box -12 -8 32 272
use FILL  FILL_7__2223_
timestamp 1701859473
transform -1 0 10030 0 -1 4430
box -12 -8 32 272
use FILL  FILL_7__2224_
timestamp 1701859473
transform -1 0 9890 0 1 4430
box -12 -8 32 272
use FILL  FILL_7__2225_
timestamp 1701859473
transform 1 0 10130 0 -1 4950
box -12 -8 32 272
use FILL  FILL_7__2226_
timestamp 1701859473
transform 1 0 9010 0 -1 7030
box -12 -8 32 272
use FILL  FILL_7__2227_
timestamp 1701859473
transform -1 0 9290 0 -1 7030
box -12 -8 32 272
use FILL  FILL_7__2229_
timestamp 1701859473
transform 1 0 4390 0 1 3390
box -12 -8 32 272
use FILL  FILL_7__2230_
timestamp 1701859473
transform -1 0 4490 0 -1 3910
box -12 -8 32 272
use FILL  FILL_7__2231_
timestamp 1701859473
transform -1 0 4270 0 -1 3910
box -12 -8 32 272
use FILL  FILL_7__2232_
timestamp 1701859473
transform 1 0 1670 0 1 2870
box -12 -8 32 272
use FILL  FILL_7__2233_
timestamp 1701859473
transform 1 0 2390 0 1 2870
box -12 -8 32 272
use FILL  FILL_7__2234_
timestamp 1701859473
transform -1 0 2650 0 1 2870
box -12 -8 32 272
use FILL  FILL_7__2236_
timestamp 1701859473
transform -1 0 5690 0 -1 3910
box -12 -8 32 272
use FILL  FILL_7__2237_
timestamp 1701859473
transform -1 0 4730 0 -1 3910
box -12 -8 32 272
use FILL  FILL_7__2238_
timestamp 1701859473
transform 1 0 4790 0 -1 4950
box -12 -8 32 272
use FILL  FILL_7__2239_
timestamp 1701859473
transform 1 0 2910 0 1 4950
box -12 -8 32 272
use FILL  FILL_7__2240_
timestamp 1701859473
transform 1 0 2470 0 1 3910
box -12 -8 32 272
use FILL  FILL_7__2241_
timestamp 1701859473
transform -1 0 2490 0 1 4950
box -12 -8 32 272
use FILL  FILL_7__2242_
timestamp 1701859473
transform 1 0 2530 0 -1 4950
box -12 -8 32 272
use FILL  FILL_7__2244_
timestamp 1701859473
transform 1 0 3130 0 1 4950
box -12 -8 32 272
use FILL  FILL_7__2245_
timestamp 1701859473
transform 1 0 2970 0 1 5990
box -12 -8 32 272
use FILL  FILL_7__2246_
timestamp 1701859473
transform 1 0 2990 0 -1 4950
box -12 -8 32 272
use FILL  FILL_7__2247_
timestamp 1701859473
transform -1 0 3110 0 -1 6510
box -12 -8 32 272
use FILL  FILL_7__2248_
timestamp 1701859473
transform 1 0 3570 0 -1 7030
box -12 -8 32 272
use FILL  FILL_7__2249_
timestamp 1701859473
transform 1 0 6350 0 1 7030
box -12 -8 32 272
use FILL  FILL_7__2251_
timestamp 1701859473
transform -1 0 10710 0 1 8070
box -12 -8 32 272
use FILL  FILL_7__2252_
timestamp 1701859473
transform -1 0 11010 0 -1 8070
box -12 -8 32 272
use FILL  FILL_7__2253_
timestamp 1701859473
transform -1 0 10770 0 -1 8070
box -12 -8 32 272
use FILL  FILL_7__2254_
timestamp 1701859473
transform 1 0 5470 0 1 8070
box -12 -8 32 272
use FILL  FILL_7__2255_
timestamp 1701859473
transform 1 0 3090 0 1 7030
box -12 -8 32 272
use FILL  FILL_7__2256_
timestamp 1701859473
transform -1 0 5210 0 1 7030
box -12 -8 32 272
use FILL  FILL_7__2258_
timestamp 1701859473
transform 1 0 5790 0 -1 8590
box -12 -8 32 272
use FILL  FILL_7__2259_
timestamp 1701859473
transform 1 0 10410 0 -1 7550
box -12 -8 32 272
use FILL  FILL_7__2260_
timestamp 1701859473
transform 1 0 9990 0 1 8070
box -12 -8 32 272
use FILL  FILL_7__2261_
timestamp 1701859473
transform -1 0 10290 0 1 7550
box -12 -8 32 272
use FILL  FILL_7__2262_
timestamp 1701859473
transform -1 0 10050 0 1 7550
box -12 -8 32 272
use FILL  FILL_7__2263_
timestamp 1701859473
transform 1 0 5550 0 1 7550
box -12 -8 32 272
use FILL  FILL_7__2265_
timestamp 1701859473
transform 1 0 1890 0 -1 6510
box -12 -8 32 272
use FILL  FILL_7__2266_
timestamp 1701859473
transform 1 0 3990 0 1 6510
box -12 -8 32 272
use FILL  FILL_7__2267_
timestamp 1701859473
transform -1 0 3750 0 -1 7550
box -12 -8 32 272
use FILL  FILL_7__2268_
timestamp 1701859473
transform 1 0 4430 0 -1 7550
box -12 -8 32 272
use FILL  FILL_7__2269_
timestamp 1701859473
transform 1 0 5750 0 1 7550
box -12 -8 32 272
use FILL  FILL_7__2270_
timestamp 1701859473
transform 1 0 8670 0 1 7550
box -12 -8 32 272
use FILL  FILL_7__2271_
timestamp 1701859473
transform -1 0 8950 0 -1 8070
box -12 -8 32 272
use FILL  FILL_7__2273_
timestamp 1701859473
transform -1 0 8710 0 -1 8070
box -12 -8 32 272
use FILL  FILL_7__2274_
timestamp 1701859473
transform -1 0 6070 0 -1 9630
box -12 -8 32 272
use FILL  FILL_7__2275_
timestamp 1701859473
transform -1 0 2370 0 1 8070
box -12 -8 32 272
use FILL  FILL_7__2276_
timestamp 1701859473
transform -1 0 3250 0 1 8070
box -12 -8 32 272
use FILL  FILL_7__2277_
timestamp 1701859473
transform -1 0 3730 0 -1 8590
box -12 -8 32 272
use FILL  FILL_7__2278_
timestamp 1701859473
transform 1 0 6630 0 1 9110
box -12 -8 32 272
use FILL  FILL_7__2280_
timestamp 1701859473
transform 1 0 10510 0 1 5990
box -12 -8 32 272
use FILL  FILL_7__2281_
timestamp 1701859473
transform -1 0 10790 0 -1 5990
box -12 -8 32 272
use FILL  FILL_7__2282_
timestamp 1701859473
transform -1 0 10570 0 -1 6510
box -12 -8 32 272
use FILL  FILL_7__2283_
timestamp 1701859473
transform 1 0 6030 0 -1 8590
box -12 -8 32 272
use FILL  FILL_7__2284_
timestamp 1701859473
transform -1 0 2150 0 1 8070
box -12 -8 32 272
use FILL  FILL_7__2285_
timestamp 1701859473
transform -1 0 4210 0 1 8070
box -12 -8 32 272
use FILL  FILL_7__2287_
timestamp 1701859473
transform -1 0 6190 0 1 8590
box -12 -8 32 272
use FILL  FILL_7__2288_
timestamp 1701859473
transform -1 0 8910 0 1 7550
box -12 -8 32 272
use FILL  FILL_7__2289_
timestamp 1701859473
transform 1 0 8570 0 1 8070
box -12 -8 32 272
use FILL  FILL_7__2290_
timestamp 1701859473
transform -1 0 10070 0 -1 8070
box -12 -8 32 272
use FILL  FILL_7__2291_
timestamp 1701859473
transform -1 0 8850 0 1 8070
box -12 -8 32 272
use FILL  FILL_7__2292_
timestamp 1701859473
transform -1 0 6290 0 -1 9110
box -12 -8 32 272
use FILL  FILL_7__2293_
timestamp 1701859473
transform -1 0 2610 0 -1 8590
box -12 -8 32 272
use FILL  FILL_7__2295_
timestamp 1701859473
transform 1 0 5010 0 1 8590
box -12 -8 32 272
use FILL  FILL_7__2296_
timestamp 1701859473
transform 1 0 6730 0 -1 9110
box -12 -8 32 272
use FILL  FILL_7__2297_
timestamp 1701859473
transform -1 0 9630 0 -1 5990
box -12 -8 32 272
use FILL  FILL_7__2298_
timestamp 1701859473
transform -1 0 10070 0 -1 5470
box -12 -8 32 272
use FILL  FILL_7__2299_
timestamp 1701859473
transform -1 0 9410 0 -1 6510
box -12 -8 32 272
use FILL  FILL_7__2300_
timestamp 1701859473
transform 1 0 9610 0 1 5990
box -12 -8 32 272
use FILL  FILL_7__2302_
timestamp 1701859473
transform -1 0 3550 0 -1 9110
box -12 -8 32 272
use FILL  FILL_7__2303_
timestamp 1701859473
transform 1 0 2670 0 1 9110
box -12 -8 32 272
use FILL  FILL_7__2304_
timestamp 1701859473
transform 1 0 2870 0 -1 9110
box -12 -8 32 272
use FILL  FILL_7__2305_
timestamp 1701859473
transform -1 0 3850 0 1 8590
box -12 -8 32 272
use FILL  FILL_7__2306_
timestamp 1701859473
transform 1 0 4530 0 1 8590
box -12 -8 32 272
use FILL  FILL_7__2307_
timestamp 1701859473
transform 1 0 6390 0 1 9110
box -12 -8 32 272
use FILL  FILL_7__2309_
timestamp 1701859473
transform -1 0 8670 0 1 5990
box -12 -8 32 272
use FILL  FILL_7__2310_
timestamp 1701859473
transform -1 0 9170 0 -1 6510
box -12 -8 32 272
use FILL  FILL_7__2311_
timestamp 1701859473
transform -1 0 8730 0 -1 6510
box -12 -8 32 272
use FILL  FILL_7__2312_
timestamp 1701859473
transform -1 0 5630 0 -1 9630
box -12 -8 32 272
use FILL  FILL_7__2313_
timestamp 1701859473
transform -1 0 1910 0 1 8590
box -12 -8 32 272
use FILL  FILL_7__2314_
timestamp 1701859473
transform 1 0 1510 0 -1 8590
box -12 -8 32 272
use FILL  FILL_7__2316_
timestamp 1701859473
transform -1 0 4310 0 1 8590
box -12 -8 32 272
use FILL  FILL_7__2317_
timestamp 1701859473
transform 1 0 4770 0 1 8590
box -12 -8 32 272
use FILL  FILL_7__2318_
timestamp 1701859473
transform 1 0 6870 0 1 9110
box -12 -8 32 272
use FILL  FILL_7__2319_
timestamp 1701859473
transform -1 0 11190 0 1 4430
box -12 -8 32 272
use FILL  FILL_7__2320_
timestamp 1701859473
transform 1 0 5170 0 1 3910
box -12 -8 32 272
use FILL  FILL_7__2321_
timestamp 1701859473
transform 1 0 6590 0 1 3910
box -12 -8 32 272
use FILL  FILL_7__2322_
timestamp 1701859473
transform -1 0 7970 0 1 3910
box -12 -8 32 272
use FILL  FILL_7__2324_
timestamp 1701859473
transform -1 0 11230 0 -1 2870
box -12 -8 32 272
use FILL  FILL_7__2325_
timestamp 1701859473
transform -1 0 8210 0 1 3910
box -12 -8 32 272
use FILL  FILL_7__2326_
timestamp 1701859473
transform -1 0 3250 0 -1 4950
box -12 -8 32 272
use FILL  FILL_7__2327_
timestamp 1701859473
transform -1 0 3450 0 -1 4950
box -12 -8 32 272
use FILL  FILL_7__2328_
timestamp 1701859473
transform 1 0 3930 0 -1 5470
box -12 -8 32 272
use FILL  FILL_7__2329_
timestamp 1701859473
transform 1 0 3690 0 -1 5470
box -12 -8 32 272
use FILL  FILL_7__2331_
timestamp 1701859473
transform 1 0 4910 0 1 3910
box -12 -8 32 272
use FILL  FILL_7__2332_
timestamp 1701859473
transform -1 0 4250 0 1 4950
box -12 -8 32 272
use FILL  FILL_7__2333_
timestamp 1701859473
transform -1 0 11210 0 -1 4430
box -12 -8 32 272
use FILL  FILL_7__2334_
timestamp 1701859473
transform 1 0 9090 0 -1 4430
box -12 -8 32 272
use FILL  FILL_7__2335_
timestamp 1701859473
transform 1 0 5270 0 -1 5470
box -12 -8 32 272
use FILL  FILL_7__2336_
timestamp 1701859473
transform -1 0 5130 0 1 5990
box -12 -8 32 272
use FILL  FILL_7__2338_
timestamp 1701859473
transform 1 0 3230 0 1 3390
box -12 -8 32 272
use FILL  FILL_7__2339_
timestamp 1701859473
transform 1 0 4810 0 1 3390
box -12 -8 32 272
use FILL  FILL_7__2340_
timestamp 1701859473
transform 1 0 5050 0 1 3390
box -12 -8 32 272
use FILL  FILL_7__2341_
timestamp 1701859473
transform -1 0 630 0 1 5990
box -12 -8 32 272
use FILL  FILL_7__2342_
timestamp 1701859473
transform 1 0 2730 0 1 5470
box -12 -8 32 272
use FILL  FILL_7__2343_
timestamp 1701859473
transform -1 0 4670 0 1 6510
box -12 -8 32 272
use FILL  FILL_7__2345_
timestamp 1701859473
transform -1 0 4750 0 1 5470
box -12 -8 32 272
use FILL  FILL_7__2346_
timestamp 1701859473
transform -1 0 4910 0 -1 5990
box -12 -8 32 272
use FILL  FILL_7__2347_
timestamp 1701859473
transform -1 0 5770 0 -1 5990
box -12 -8 32 272
use FILL  FILL_7__2348_
timestamp 1701859473
transform 1 0 5330 0 -1 6510
box -12 -8 32 272
use FILL  FILL_7__2349_
timestamp 1701859473
transform -1 0 5110 0 -1 6510
box -12 -8 32 272
use FILL  FILL_7__2350_
timestamp 1701859473
transform -1 0 4530 0 -1 6510
box -12 -8 32 272
use FILL  FILL_7__2351_
timestamp 1701859473
transform 1 0 5670 0 1 7030
box -12 -8 32 272
use FILL  FILL_7__2353_
timestamp 1701859473
transform -1 0 830 0 1 7030
box -12 -8 32 272
use FILL  FILL_7__2354_
timestamp 1701859473
transform 1 0 5530 0 -1 5990
box -12 -8 32 272
use FILL  FILL_7__2355_
timestamp 1701859473
transform 1 0 5430 0 1 7030
box -12 -8 32 272
use FILL  FILL_7__2356_
timestamp 1701859473
transform -1 0 4930 0 -1 7550
box -12 -8 32 272
use FILL  FILL_7__2357_
timestamp 1701859473
transform 1 0 4790 0 1 8070
box -12 -8 32 272
use FILL  FILL_7__2358_
timestamp 1701859473
transform 1 0 5270 0 1 8070
box -12 -8 32 272
use FILL  FILL_7__2360_
timestamp 1701859473
transform -1 0 830 0 -1 6510
box -12 -8 32 272
use FILL  FILL_7__2361_
timestamp 1701859473
transform -1 0 5330 0 1 5990
box -12 -8 32 272
use FILL  FILL_7__2362_
timestamp 1701859473
transform 1 0 5330 0 1 6510
box -12 -8 32 272
use FILL  FILL_7__2363_
timestamp 1701859473
transform 1 0 5350 0 -1 7030
box -12 -8 32 272
use FILL  FILL_7__2364_
timestamp 1701859473
transform 1 0 5350 0 -1 8070
box -12 -8 32 272
use FILL  FILL_7__2365_
timestamp 1701859473
transform 1 0 5590 0 -1 8070
box -12 -8 32 272
use FILL  FILL_7__2367_
timestamp 1701859473
transform 1 0 2770 0 -1 7550
box -12 -8 32 272
use FILL  FILL_7__2368_
timestamp 1701859473
transform -1 0 5610 0 -1 7030
box -12 -8 32 272
use FILL  FILL_7__2369_
timestamp 1701859473
transform 1 0 5310 0 1 7550
box -12 -8 32 272
use FILL  FILL_7__2370_
timestamp 1701859473
transform -1 0 5350 0 -1 8590
box -12 -8 32 272
use FILL  FILL_7__2371_
timestamp 1701859473
transform 1 0 6030 0 -1 9110
box -12 -8 32 272
use FILL  FILL_7__2372_
timestamp 1701859473
transform 1 0 6190 0 1 9110
box -12 -8 32 272
use FILL  FILL_7__2373_
timestamp 1701859473
transform -1 0 6270 0 -1 9630
box -12 -8 32 272
use FILL  FILL_7__2375_
timestamp 1701859473
transform -1 0 4290 0 1 5470
box -12 -8 32 272
use FILL  FILL_7__2376_
timestamp 1701859473
transform 1 0 4630 0 -1 5990
box -12 -8 32 272
use FILL  FILL_7__2377_
timestamp 1701859473
transform -1 0 4050 0 -1 6510
box -12 -8 32 272
use FILL  FILL_7__2378_
timestamp 1701859473
transform 1 0 3790 0 -1 6510
box -12 -8 32 272
use FILL  FILL_7__2379_
timestamp 1701859473
transform -1 0 5110 0 1 6510
box -12 -8 32 272
use FILL  FILL_7__2380_
timestamp 1701859473
transform -1 0 4890 0 -1 8590
box -12 -8 32 272
use FILL  FILL_7__2382_
timestamp 1701859473
transform -1 0 4650 0 -1 8590
box -12 -8 32 272
use FILL  FILL_7__2383_
timestamp 1701859473
transform -1 0 5730 0 1 8590
box -12 -8 32 272
use FILL  FILL_7__2384_
timestamp 1701859473
transform -1 0 5950 0 1 8590
box -12 -8 32 272
use FILL  FILL_7__2385_
timestamp 1701859473
transform 1 0 1330 0 -1 10150
box -12 -8 32 272
use FILL  FILL_7__2386_
timestamp 1701859473
transform 1 0 5590 0 -1 7550
box -12 -8 32 272
use FILL  FILL_7__2387_
timestamp 1701859473
transform 1 0 5570 0 -1 9110
box -12 -8 32 272
use FILL  FILL_7__2389_
timestamp 1701859473
transform -1 0 5150 0 -1 9630
box -12 -8 32 272
use FILL  FILL_7__2390_
timestamp 1701859473
transform 1 0 5210 0 1 9630
box -12 -8 32 272
use FILL  FILL_7__2391_
timestamp 1701859473
transform -1 0 5430 0 1 9630
box -12 -8 32 272
use FILL  FILL_7__2392_
timestamp 1701859473
transform 1 0 1530 0 -1 10150
box -12 -8 32 272
use FILL  FILL_7__2393_
timestamp 1701859473
transform -1 0 5390 0 -1 7550
box -12 -8 32 272
use FILL  FILL_7__2394_
timestamp 1701859473
transform 1 0 5470 0 1 8590
box -12 -8 32 272
use FILL  FILL_7__2396_
timestamp 1701859473
transform 1 0 5750 0 1 9110
box -12 -8 32 272
use FILL  FILL_7__2397_
timestamp 1701859473
transform 1 0 5990 0 1 9110
box -12 -8 32 272
use FILL  FILL_7__2398_
timestamp 1701859473
transform 1 0 5810 0 -1 9630
box -12 -8 32 272
use FILL  FILL_7__2399_
timestamp 1701859473
transform -1 0 3250 0 -1 5470
box -12 -8 32 272
use FILL  FILL_7__2400_
timestamp 1701859473
transform -1 0 3430 0 1 5990
box -12 -8 32 272
use FILL  FILL_7__2401_
timestamp 1701859473
transform 1 0 3350 0 -1 6510
box -12 -8 32 272
use FILL  FILL_7__2402_
timestamp 1701859473
transform -1 0 2290 0 -1 4430
box -12 -8 32 272
use FILL  FILL_7__2404_
timestamp 1701859473
transform -1 0 3010 0 -1 5470
box -12 -8 32 272
use FILL  FILL_7__2405_
timestamp 1701859473
transform 1 0 2390 0 -1 2870
box -12 -8 32 272
use FILL  FILL_7__2406_
timestamp 1701859473
transform 1 0 3090 0 -1 3390
box -12 -8 32 272
use FILL  FILL_7__2407_
timestamp 1701859473
transform -1 0 3230 0 1 5470
box -12 -8 32 272
use FILL  FILL_7__2408_
timestamp 1701859473
transform 1 0 850 0 -1 2870
box -12 -8 32 272
use FILL  FILL_7__2409_
timestamp 1701859473
transform 1 0 870 0 -1 3910
box -12 -8 32 272
use FILL  FILL_7__2411_
timestamp 1701859473
transform -1 0 830 0 -1 4950
box -12 -8 32 272
use FILL  FILL_7__2412_
timestamp 1701859473
transform 1 0 2510 0 -1 5990
box -12 -8 32 272
use FILL  FILL_7__2413_
timestamp 1701859473
transform 1 0 2970 0 1 5470
box -12 -8 32 272
use FILL  FILL_7__2414_
timestamp 1701859473
transform 1 0 4130 0 -1 5470
box -12 -8 32 272
use FILL  FILL_7__2415_
timestamp 1701859473
transform -1 0 4070 0 1 7030
box -12 -8 32 272
use FILL  FILL_7__2416_
timestamp 1701859473
transform 1 0 4030 0 1 4950
box -12 -8 32 272
use FILL  FILL_7__2418_
timestamp 1701859473
transform -1 0 1630 0 -1 4950
box -12 -8 32 272
use FILL  FILL_7__2419_
timestamp 1701859473
transform 1 0 2210 0 1 4430
box -12 -8 32 272
use FILL  FILL_7__2420_
timestamp 1701859473
transform 1 0 3870 0 1 5990
box -12 -8 32 272
use FILL  FILL_7__2421_
timestamp 1701859473
transform -1 0 3650 0 1 5990
box -12 -8 32 272
use FILL  FILL_7__2422_
timestamp 1701859473
transform -1 0 3530 0 -1 5990
box -12 -8 32 272
use FILL  FILL_7__2423_
timestamp 1701859473
transform -1 0 3750 0 -1 5990
box -12 -8 32 272
use FILL  FILL_7__2424_
timestamp 1701859473
transform 1 0 3290 0 -1 5990
box -12 -8 32 272
use FILL  FILL_7__2426_
timestamp 1701859473
transform 1 0 4030 0 -1 7030
box -12 -8 32 272
use FILL  FILL_7__2427_
timestamp 1701859473
transform 1 0 4850 0 1 5990
box -12 -8 32 272
use FILL  FILL_7__2428_
timestamp 1701859473
transform 1 0 4610 0 1 5990
box -12 -8 32 272
use FILL  FILL_7__2429_
timestamp 1701859473
transform -1 0 4290 0 -1 6510
box -12 -8 32 272
use FILL  FILL_7__2430_
timestamp 1701859473
transform 1 0 4850 0 1 6510
box -12 -8 32 272
use FILL  FILL_7__2431_
timestamp 1701859473
transform -1 0 4950 0 -1 7030
box -12 -8 32 272
use FILL  FILL_7__2433_
timestamp 1701859473
transform -1 0 4430 0 -1 8070
box -12 -8 32 272
use FILL  FILL_7__2434_
timestamp 1701859473
transform 1 0 4910 0 1 7550
box -12 -8 32 272
use FILL  FILL_7__2435_
timestamp 1701859473
transform 1 0 4250 0 1 7030
box -12 -8 32 272
use FILL  FILL_7__2436_
timestamp 1701859473
transform -1 0 4690 0 -1 7550
box -12 -8 32 272
use FILL  FILL_7__2437_
timestamp 1701859473
transform -1 0 4670 0 -1 8070
box -12 -8 32 272
use FILL  FILL_7__2438_
timestamp 1701859473
transform -1 0 4910 0 -1 8070
box -12 -8 32 272
use FILL  FILL_7__2440_
timestamp 1701859473
transform 1 0 4690 0 1 10150
box -12 -8 32 272
use FILL  FILL_7__2441_
timestamp 1701859473
transform 1 0 3970 0 -1 7550
box -12 -8 32 272
use FILL  FILL_7__2442_
timestamp 1701859473
transform -1 0 4190 0 -1 8070
box -12 -8 32 272
use FILL  FILL_7__2443_
timestamp 1701859473
transform -1 0 3970 0 1 8070
box -12 -8 32 272
use FILL  FILL_7__2444_
timestamp 1701859473
transform 1 0 3710 0 1 8070
box -12 -8 32 272
use FILL  FILL_7__2445_
timestamp 1701859473
transform -1 0 4690 0 1 7550
box -12 -8 32 272
use FILL  FILL_7__2447_
timestamp 1701859473
transform 1 0 4350 0 1 9110
box -12 -8 32 272
use FILL  FILL_7__2448_
timestamp 1701859473
transform 1 0 5010 0 1 9110
box -12 -8 32 272
use FILL  FILL_7__2449_
timestamp 1701859473
transform 1 0 5270 0 1 9110
box -12 -8 32 272
use FILL  FILL_7__2450_
timestamp 1701859473
transform 1 0 5510 0 1 9110
box -12 -8 32 272
use FILL  FILL_7__2451_
timestamp 1701859473
transform -1 0 5390 0 -1 9630
box -12 -8 32 272
use FILL  FILL_7__2452_
timestamp 1701859473
transform -1 0 5310 0 -1 10670
box -12 -8 32 272
use FILL  FILL_7__2453_
timestamp 1701859473
transform 1 0 3850 0 -1 10150
box -12 -8 32 272
use FILL  FILL_7__2455_
timestamp 1701859473
transform 1 0 3930 0 -1 8070
box -12 -8 32 272
use FILL  FILL_7__2456_
timestamp 1701859473
transform -1 0 3710 0 -1 8070
box -12 -8 32 272
use FILL  FILL_7__2457_
timestamp 1701859473
transform 1 0 3470 0 1 8070
box -12 -8 32 272
use FILL  FILL_7__2458_
timestamp 1701859473
transform -1 0 4410 0 -1 8590
box -12 -8 32 272
use FILL  FILL_7__2459_
timestamp 1701859473
transform -1 0 4570 0 -1 11190
box -12 -8 32 272
use FILL  FILL_7__2460_
timestamp 1701859473
transform 1 0 4210 0 -1 10670
box -12 -8 32 272
use FILL  FILL_7__2462_
timestamp 1701859473
transform -1 0 4650 0 -1 9110
box -12 -8 32 272
use FILL  FILL_7__2463_
timestamp 1701859473
transform -1 0 4890 0 -1 9110
box -12 -8 32 272
use FILL  FILL_7__2464_
timestamp 1701859473
transform -1 0 5130 0 -1 9110
box -12 -8 32 272
use FILL  FILL_7__2465_
timestamp 1701859473
transform -1 0 4990 0 -1 11190
box -12 -8 32 272
use FILL  FILL_7__2466_
timestamp 1701859473
transform -1 0 4070 0 -1 10150
box -12 -8 32 272
use FILL  FILL_7__2467_
timestamp 1701859473
transform -1 0 4170 0 -1 9630
box -12 -8 32 272
use FILL  FILL_7__2469_
timestamp 1701859473
transform -1 0 4290 0 1 9630
box -12 -8 32 272
use FILL  FILL_7__2470_
timestamp 1701859473
transform -1 0 4530 0 1 9630
box -12 -8 32 272
use FILL  FILL_7__2471_
timestamp 1701859473
transform -1 0 5110 0 -1 10670
box -12 -8 32 272
use FILL  FILL_7__2472_
timestamp 1701859473
transform 1 0 4070 0 1 9630
box -12 -8 32 272
use FILL  FILL_7__2473_
timestamp 1701859473
transform 1 0 4630 0 -1 9630
box -12 -8 32 272
use FILL  FILL_7__2474_
timestamp 1701859473
transform -1 0 4910 0 -1 9630
box -12 -8 32 272
use FILL  FILL_7__2476_
timestamp 1701859473
transform -1 0 4990 0 1 9630
box -12 -8 32 272
use FILL  FILL_7__2477_
timestamp 1701859473
transform 1 0 4930 0 1 10670
box -12 -8 32 272
use FILL  FILL_7__2478_
timestamp 1701859473
transform 1 0 3170 0 1 5990
box -12 -8 32 272
use FILL  FILL_7__2479_
timestamp 1701859473
transform -1 0 2730 0 1 5990
box -12 -8 32 272
use FILL  FILL_7__2480_
timestamp 1701859473
transform -1 0 2750 0 -1 5990
box -12 -8 32 272
use FILL  FILL_7__2481_
timestamp 1701859473
transform -1 0 2990 0 -1 5990
box -12 -8 32 272
use FILL  FILL_7__2482_
timestamp 1701859473
transform 1 0 1570 0 -1 5990
box -12 -8 32 272
use FILL  FILL_7__2484_
timestamp 1701859473
transform -1 0 2010 0 1 6510
box -12 -8 32 272
use FILL  FILL_7__2485_
timestamp 1701859473
transform -1 0 2210 0 1 6510
box -12 -8 32 272
use FILL  FILL_7__2486_
timestamp 1701859473
transform 1 0 2410 0 -1 7030
box -12 -8 32 272
use FILL  FILL_7__2487_
timestamp 1701859473
transform 1 0 2170 0 -1 7030
box -12 -8 32 272
use FILL  FILL_7__2488_
timestamp 1701859473
transform -1 0 1970 0 -1 7030
box -12 -8 32 272
use FILL  FILL_7__2489_
timestamp 1701859473
transform 1 0 1470 0 -1 7030
box -12 -8 32 272
use FILL  FILL_7__2491_
timestamp 1701859473
transform 1 0 1270 0 1 5470
box -12 -8 32 272
use FILL  FILL_7__2492_
timestamp 1701859473
transform -1 0 2130 0 -1 6510
box -12 -8 32 272
use FILL  FILL_7__2493_
timestamp 1701859473
transform 1 0 2010 0 1 5990
box -12 -8 32 272
use FILL  FILL_7__2494_
timestamp 1701859473
transform -1 0 1570 0 1 5990
box -12 -8 32 272
use FILL  FILL_7__2495_
timestamp 1701859473
transform 1 0 1310 0 1 5990
box -12 -8 32 272
use FILL  FILL_7__2496_
timestamp 1701859473
transform 1 0 1710 0 -1 7030
box -12 -8 32 272
use FILL  FILL_7__2498_
timestamp 1701859473
transform 1 0 850 0 1 8070
box -12 -8 32 272
use FILL  FILL_7__2499_
timestamp 1701859473
transform 1 0 2530 0 1 7550
box -12 -8 32 272
use FILL  FILL_7__2500_
timestamp 1701859473
transform 1 0 1950 0 1 7550
box -12 -8 32 272
use FILL  FILL_7__2501_
timestamp 1701859473
transform 1 0 1730 0 1 7550
box -12 -8 32 272
use FILL  FILL_7__2502_
timestamp 1701859473
transform -1 0 1270 0 1 7550
box -12 -8 32 272
use FILL  FILL_7__2503_
timestamp 1701859473
transform -1 0 1510 0 1 8070
box -12 -8 32 272
use FILL  FILL_7__2504_
timestamp 1701859473
transform -1 0 1930 0 1 8070
box -12 -8 32 272
use FILL  FILL_7__2506_
timestamp 1701859473
transform -1 0 1790 0 -1 8070
box -12 -8 32 272
use FILL  FILL_7__2507_
timestamp 1701859473
transform 1 0 1530 0 -1 8070
box -12 -8 32 272
use FILL  FILL_7__2508_
timestamp 1701859473
transform 1 0 1050 0 1 8070
box -12 -8 32 272
use FILL  FILL_7__2509_
timestamp 1701859473
transform 1 0 610 0 -1 8590
box -12 -8 32 272
use FILL  FILL_7__2510_
timestamp 1701859473
transform -1 0 1550 0 1 9110
box -12 -8 32 272
use FILL  FILL_7__2511_
timestamp 1701859473
transform -1 0 1490 0 -1 9630
box -12 -8 32 272
use FILL  FILL_7__2513_
timestamp 1701859473
transform -1 0 1050 0 1 8590
box -12 -8 32 272
use FILL  FILL_7__2514_
timestamp 1701859473
transform 1 0 2130 0 -1 8590
box -12 -8 32 272
use FILL  FILL_7__2515_
timestamp 1701859473
transform 1 0 1250 0 -1 9110
box -12 -8 32 272
use FILL  FILL_7__2516_
timestamp 1701859473
transform -1 0 1090 0 1 9110
box -12 -8 32 272
use FILL  FILL_7__2517_
timestamp 1701859473
transform -1 0 850 0 1 9110
box -12 -8 32 272
use FILL  FILL_7__2518_
timestamp 1701859473
transform 1 0 1710 0 -1 9630
box -12 -8 32 272
use FILL  FILL_7__2520_
timestamp 1701859473
transform -1 0 2650 0 -1 9110
box -12 -8 32 272
use FILL  FILL_7__2521_
timestamp 1701859473
transform 1 0 2390 0 -1 9110
box -12 -8 32 272
use FILL  FILL_7__2522_
timestamp 1701859473
transform -1 0 2010 0 1 9630
box -12 -8 32 272
use FILL  FILL_7__2523_
timestamp 1701859473
transform -1 0 2230 0 1 9630
box -12 -8 32 272
use FILL  FILL_7__2524_
timestamp 1701859473
transform -1 0 1970 0 -1 9110
box -12 -8 32 272
use FILL  FILL_7__2525_
timestamp 1701859473
transform 1 0 850 0 -1 8590
box -12 -8 32 272
use FILL  FILL_7__2527_
timestamp 1701859473
transform -1 0 1290 0 -1 8590
box -12 -8 32 272
use FILL  FILL_7__2528_
timestamp 1701859473
transform -1 0 1070 0 -1 8590
box -12 -8 32 272
use FILL  FILL_7__2529_
timestamp 1701859473
transform -1 0 1310 0 1 9110
box -12 -8 32 272
use FILL  FILL_7__2530_
timestamp 1701859473
transform -1 0 7570 0 -1 6510
box -12 -8 32 272
use FILL  FILL_7__2531_
timestamp 1701859473
transform 1 0 7990 0 1 7550
box -12 -8 32 272
use FILL  FILL_7__2532_
timestamp 1701859473
transform -1 0 9890 0 1 2870
box -12 -8 32 272
use FILL  FILL_7__2533_
timestamp 1701859473
transform -1 0 8970 0 1 4430
box -12 -8 32 272
use FILL  FILL_7__2535_
timestamp 1701859473
transform 1 0 150 0 -1 4950
box -12 -8 32 272
use FILL  FILL_7__2536_
timestamp 1701859473
transform 1 0 710 0 1 4950
box -12 -8 32 272
use FILL  FILL_7__2537_
timestamp 1701859473
transform 1 0 850 0 1 3390
box -12 -8 32 272
use FILL  FILL_7__2538_
timestamp 1701859473
transform -1 0 410 0 -1 3910
box -12 -8 32 272
use FILL  FILL_7__2539_
timestamp 1701859473
transform -1 0 170 0 1 4950
box -12 -8 32 272
use FILL  FILL_7__2540_
timestamp 1701859473
transform 1 0 3110 0 1 2350
box -12 -8 32 272
use FILL  FILL_7__2542_
timestamp 1701859473
transform -1 0 2370 0 -1 6510
box -12 -8 32 272
use FILL  FILL_7__2543_
timestamp 1701859473
transform 1 0 930 0 1 4950
box -12 -8 32 272
use FILL  FILL_7__2544_
timestamp 1701859473
transform 1 0 1490 0 1 4430
box -12 -8 32 272
use FILL  FILL_7__2545_
timestamp 1701859473
transform 1 0 1350 0 -1 5470
box -12 -8 32 272
use FILL  FILL_7__2546_
timestamp 1701859473
transform -1 0 2090 0 -1 5470
box -12 -8 32 272
use FILL  FILL_7__2547_
timestamp 1701859473
transform 1 0 2030 0 -1 4430
box -12 -8 32 272
use FILL  FILL_7__2549_
timestamp 1701859473
transform 1 0 1370 0 1 4950
box -12 -8 32 272
use FILL  FILL_7__2550_
timestamp 1701859473
transform -1 0 1850 0 -1 5470
box -12 -8 32 272
use FILL  FILL_7__2551_
timestamp 1701859473
transform 1 0 2630 0 -1 9630
box -12 -8 32 272
use FILL  FILL_7__2552_
timestamp 1701859473
transform 1 0 3470 0 -1 5470
box -12 -8 32 272
use FILL  FILL_7__2553_
timestamp 1701859473
transform -1 0 2850 0 -1 6510
box -12 -8 32 272
use FILL  FILL_7__2554_
timestamp 1701859473
transform -1 0 3310 0 1 6510
box -12 -8 32 272
use FILL  FILL_7__2556_
timestamp 1701859473
transform -1 0 2870 0 1 6510
box -12 -8 32 272
use FILL  FILL_7__2557_
timestamp 1701859473
transform 1 0 2570 0 -1 6510
box -12 -8 32 272
use FILL  FILL_7__2558_
timestamp 1701859473
transform 1 0 3310 0 -1 7550
box -12 -8 32 272
use FILL  FILL_7__2559_
timestamp 1701859473
transform 1 0 3510 0 -1 7550
box -12 -8 32 272
use FILL  FILL_7__2560_
timestamp 1701859473
transform -1 0 3570 0 1 7030
box -12 -8 32 272
use FILL  FILL_7__2561_
timestamp 1701859473
transform -1 0 1590 0 1 4950
box -12 -8 32 272
use FILL  FILL_7__2562_
timestamp 1701859473
transform 1 0 3310 0 1 7030
box -12 -8 32 272
use FILL  FILL_7__2564_
timestamp 1701859473
transform -1 0 3750 0 1 6510
box -12 -8 32 272
use FILL  FILL_7__2565_
timestamp 1701859473
transform 1 0 3810 0 1 7030
box -12 -8 32 272
use FILL  FILL_7__2566_
timestamp 1701859473
transform 1 0 3270 0 1 7550
box -12 -8 32 272
use FILL  FILL_7__2567_
timestamp 1701859473
transform 1 0 3230 0 -1 8070
box -12 -8 32 272
use FILL  FILL_7__2568_
timestamp 1701859473
transform -1 0 3050 0 -1 8590
box -12 -8 32 272
use FILL  FILL_7__2569_
timestamp 1701859473
transform 1 0 2810 0 -1 8590
box -12 -8 32 272
use FILL  FILL_7__2571_
timestamp 1701859473
transform -1 0 3950 0 -1 9630
box -12 -8 32 272
use FILL  FILL_7__2572_
timestamp 1701859473
transform -1 0 3970 0 -1 5990
box -12 -8 32 272
use FILL  FILL_7__2573_
timestamp 1701859473
transform -1 0 3830 0 -1 7030
box -12 -8 32 272
use FILL  FILL_7__2574_
timestamp 1701859473
transform 1 0 3550 0 -1 6510
box -12 -8 32 272
use FILL  FILL_7__2575_
timestamp 1701859473
transform 1 0 3450 0 -1 8070
box -12 -8 32 272
use FILL  FILL_7__2576_
timestamp 1701859473
transform -1 0 3490 0 -1 8590
box -12 -8 32 272
use FILL  FILL_7__2578_
timestamp 1701859473
transform 1 0 3870 0 1 9110
box -12 -8 32 272
use FILL  FILL_7__2579_
timestamp 1701859473
transform -1 0 2850 0 -1 9630
box -12 -8 32 272
use FILL  FILL_7__2580_
timestamp 1701859473
transform -1 0 4210 0 -1 9110
box -12 -8 32 272
use FILL  FILL_7__2581_
timestamp 1701859473
transform -1 0 4130 0 1 9110
box -12 -8 32 272
use FILL  FILL_7__2582_
timestamp 1701859473
transform 1 0 3630 0 1 9110
box -12 -8 32 272
use FILL  FILL_7__2583_
timestamp 1701859473
transform 1 0 3130 0 1 9110
box -12 -8 32 272
use FILL  FILL_7__2584_
timestamp 1701859473
transform 1 0 2890 0 1 9110
box -12 -8 32 272
use FILL  FILL_7__2586_
timestamp 1701859473
transform 1 0 3150 0 1 9630
box -12 -8 32 272
use FILL  FILL_7__2587_
timestamp 1701859473
transform 1 0 3730 0 -1 9110
box -12 -8 32 272
use FILL  FILL_7__2588_
timestamp 1701859473
transform 1 0 3330 0 1 8590
box -12 -8 32 272
use FILL  FILL_7__2589_
timestamp 1701859473
transform 1 0 3170 0 -1 10150
box -12 -8 32 272
use FILL  FILL_7__2590_
timestamp 1701859473
transform 1 0 2910 0 -1 10150
box -12 -8 32 272
use FILL  FILL_7__2591_
timestamp 1701859473
transform -1 0 3670 0 -1 11190
box -12 -8 32 272
use FILL  FILL_7__2593_
timestamp 1701859473
transform -1 0 3250 0 -1 9630
box -12 -8 32 272
use FILL  FILL_7__2594_
timestamp 1701859473
transform -1 0 3410 0 -1 10150
box -12 -8 32 272
use FILL  FILL_7__2595_
timestamp 1701859473
transform 1 0 3130 0 -1 11190
box -12 -8 32 272
use FILL  FILL_7__2596_
timestamp 1701859473
transform 1 0 3410 0 -1 11190
box -12 -8 32 272
use FILL  FILL_7__2597_
timestamp 1701859473
transform 1 0 2870 0 -1 10670
box -12 -8 32 272
use FILL  FILL_7__2598_
timestamp 1701859473
transform -1 0 3610 0 1 9630
box -12 -8 32 272
use FILL  FILL_7__2600_
timestamp 1701859473
transform -1 0 3110 0 1 10150
box -12 -8 32 272
use FILL  FILL_7__2601_
timestamp 1701859473
transform 1 0 3070 0 -1 10670
box -12 -8 32 272
use FILL  FILL_7__2602_
timestamp 1701859473
transform -1 0 3330 0 -1 10670
box -12 -8 32 272
use FILL  FILL_7__2603_
timestamp 1701859473
transform 1 0 3530 0 -1 10670
box -12 -8 32 272
use FILL  FILL_7__2604_
timestamp 1701859473
transform 1 0 3330 0 1 10150
box -12 -8 32 272
use FILL  FILL_7__2605_
timestamp 1701859473
transform 1 0 2450 0 1 10670
box -12 -8 32 272
use FILL  FILL_7__2607_
timestamp 1701859473
transform -1 0 2890 0 1 10670
box -12 -8 32 272
use FILL  FILL_7__2608_
timestamp 1701859473
transform -1 0 3850 0 1 9630
box -12 -8 32 272
use FILL  FILL_7__2609_
timestamp 1701859473
transform -1 0 2470 0 1 9630
box -12 -8 32 272
use FILL  FILL_7__2610_
timestamp 1701859473
transform -1 0 2690 0 -1 10150
box -12 -8 32 272
use FILL  FILL_7__2611_
timestamp 1701859473
transform -1 0 2410 0 -1 10670
box -12 -8 32 272
use FILL  FILL_7__2612_
timestamp 1701859473
transform 1 0 2630 0 -1 10670
box -12 -8 32 272
use FILL  FILL_7__2613_
timestamp 1701859473
transform 1 0 1950 0 1 10670
box -12 -8 32 272
use FILL  FILL_7__2615_
timestamp 1701859473
transform -1 0 2470 0 -1 11190
box -12 -8 32 272
use FILL  FILL_7__2616_
timestamp 1701859473
transform -1 0 3490 0 -1 9630
box -12 -8 32 272
use FILL  FILL_7__2617_
timestamp 1701859473
transform 1 0 2390 0 -1 9630
box -12 -8 32 272
use FILL  FILL_7__2618_
timestamp 1701859473
transform -1 0 2670 0 1 10150
box -12 -8 32 272
use FILL  FILL_7__2619_
timestamp 1701859473
transform 1 0 2170 0 1 10670
box -12 -8 32 272
use FILL  FILL_7__2620_
timestamp 1701859473
transform 1 0 2210 0 -1 11190
box -12 -8 32 272
use FILL  FILL_7__2622_
timestamp 1701859473
transform -1 0 1330 0 -1 5990
box -12 -8 32 272
use FILL  FILL_7__2623_
timestamp 1701859473
transform 1 0 2550 0 -1 5470
box -12 -8 32 272
use FILL  FILL_7__2624_
timestamp 1701859473
transform -1 0 2510 0 1 5470
box -12 -8 32 272
use FILL  FILL_7__2625_
timestamp 1701859473
transform 1 0 2310 0 -1 5470
box -12 -8 32 272
use FILL  FILL_7__2626_
timestamp 1701859473
transform -1 0 1050 0 -1 5470
box -12 -8 32 272
use FILL  FILL_7__2627_
timestamp 1701859473
transform -1 0 1570 0 1 3910
box -12 -8 32 272
use FILL  FILL_7__2629_
timestamp 1701859473
transform -1 0 850 0 -1 5470
box -12 -8 32 272
use FILL  FILL_7__2630_
timestamp 1701859473
transform 1 0 830 0 -1 5990
box -12 -8 32 272
use FILL  FILL_7__2631_
timestamp 1701859473
transform -1 0 830 0 1 5990
box -12 -8 32 272
use FILL  FILL_7__2632_
timestamp 1701859473
transform 1 0 2210 0 1 10150
box -12 -8 32 272
use FILL  FILL_7__2633_
timestamp 1701859473
transform -1 0 2450 0 1 10150
box -12 -8 32 272
use FILL  FILL_7__2634_
timestamp 1701859473
transform 1 0 2410 0 -1 10150
box -12 -8 32 272
use FILL  FILL_7__2635_
timestamp 1701859473
transform 1 0 2190 0 -1 10150
box -12 -8 32 272
use FILL  FILL_7__2637_
timestamp 1701859473
transform -1 0 630 0 1 6510
box -12 -8 32 272
use FILL  FILL_7__2638_
timestamp 1701859473
transform -1 0 410 0 1 6510
box -12 -8 32 272
use FILL  FILL_7__2639_
timestamp 1701859473
transform -1 0 390 0 -1 6510
box -12 -8 32 272
use FILL  FILL_7__2640_
timestamp 1701859473
transform -1 0 390 0 1 5990
box -12 -8 32 272
use FILL  FILL_7__2641_
timestamp 1701859473
transform 1 0 150 0 -1 7550
box -12 -8 32 272
use FILL  FILL_7__2642_
timestamp 1701859473
transform -1 0 490 0 1 4950
box -12 -8 32 272
use FILL  FILL_7__2644_
timestamp 1701859473
transform 1 0 2670 0 -1 7030
box -12 -8 32 272
use FILL  FILL_7__2645_
timestamp 1701859473
transform 1 0 2850 0 1 7030
box -12 -8 32 272
use FILL  FILL_7__2646_
timestamp 1701859473
transform 1 0 2150 0 1 7030
box -12 -8 32 272
use FILL  FILL_7__2647_
timestamp 1701859473
transform 1 0 830 0 1 7550
box -12 -8 32 272
use FILL  FILL_7__2648_
timestamp 1701859473
transform 1 0 370 0 1 7550
box -12 -8 32 272
use FILL  FILL_7__2649_
timestamp 1701859473
transform 1 0 350 0 -1 7550
box -12 -8 32 272
use FILL  FILL_7__2651_
timestamp 1701859473
transform 1 0 570 0 -1 7550
box -12 -8 32 272
use FILL  FILL_7__2652_
timestamp 1701859473
transform 1 0 570 0 1 7030
box -12 -8 32 272
use FILL  FILL_7__2653_
timestamp 1701859473
transform 1 0 150 0 1 7550
box -12 -8 32 272
use FILL  FILL_7__2654_
timestamp 1701859473
transform -1 0 630 0 1 7550
box -12 -8 32 272
use FILL  FILL_7__2655_
timestamp 1701859473
transform 1 0 1950 0 1 7030
box -12 -8 32 272
use FILL  FILL_7__2656_
timestamp 1701859473
transform 1 0 1590 0 -1 5470
box -12 -8 32 272
use FILL  FILL_7__2658_
timestamp 1701859473
transform -1 0 2270 0 1 5470
box -12 -8 32 272
use FILL  FILL_7__2659_
timestamp 1701859473
transform 1 0 2030 0 -1 5990
box -12 -8 32 272
use FILL  FILL_7__2660_
timestamp 1701859473
transform -1 0 2030 0 1 5470
box -12 -8 32 272
use FILL  FILL_7__2661_
timestamp 1701859473
transform -1 0 1710 0 1 5470
box -12 -8 32 272
use FILL  FILL_7__2662_
timestamp 1701859473
transform 1 0 810 0 1 5470
box -12 -8 32 272
use FILL  FILL_7__2663_
timestamp 1701859473
transform -1 0 1090 0 -1 5990
box -12 -8 32 272
use FILL  FILL_7__2664_
timestamp 1701859473
transform 1 0 810 0 -1 7030
box -12 -8 32 272
use FILL  FILL_7__2666_
timestamp 1701859473
transform 1 0 1470 0 1 7030
box -12 -8 32 272
use FILL  FILL_7__2667_
timestamp 1701859473
transform 1 0 1010 0 -1 7030
box -12 -8 32 272
use FILL  FILL_7__2668_
timestamp 1701859473
transform -1 0 2810 0 1 7550
box -12 -8 32 272
use FILL  FILL_7__2669_
timestamp 1701859473
transform 1 0 2750 0 -1 8070
box -12 -8 32 272
use FILL  FILL_7__2670_
timestamp 1701859473
transform 1 0 2010 0 -1 8070
box -12 -8 32 272
use FILL  FILL_7__2671_
timestamp 1701859473
transform -1 0 1510 0 1 7550
box -12 -8 32 272
use FILL  FILL_7__2673_
timestamp 1701859473
transform -1 0 1430 0 -1 7550
box -12 -8 32 272
use FILL  FILL_7__2674_
timestamp 1701859473
transform 1 0 1710 0 1 7030
box -12 -8 32 272
use FILL  FILL_7__2675_
timestamp 1701859473
transform 1 0 1650 0 -1 7550
box -12 -8 32 272
use FILL  FILL_7__2676_
timestamp 1701859473
transform -1 0 2090 0 -1 7550
box -12 -8 32 272
use FILL  FILL_7__2677_
timestamp 1701859473
transform 1 0 2490 0 -1 8070
box -12 -8 32 272
use FILL  FILL_7__2678_
timestamp 1701859473
transform -1 0 2270 0 -1 8070
box -12 -8 32 272
use FILL  FILL_7__2680_
timestamp 1701859473
transform -1 0 390 0 -1 8590
box -12 -8 32 272
use FILL  FILL_7__2681_
timestamp 1701859473
transform 1 0 1010 0 -1 7550
box -12 -8 32 272
use FILL  FILL_7__2682_
timestamp 1701859473
transform -1 0 390 0 -1 8070
box -12 -8 32 272
use FILL  FILL_7__2683_
timestamp 1701859473
transform -1 0 170 0 -1 9630
box -12 -8 32 272
use FILL  FILL_7__2684_
timestamp 1701859473
transform -1 0 170 0 1 10150
box -12 -8 32 272
use FILL  FILL_7__2685_
timestamp 1701859473
transform 1 0 1050 0 1 5990
box -12 -8 32 272
use FILL  FILL_7__2687_
timestamp 1701859473
transform -1 0 1030 0 -1 10150
box -12 -8 32 272
use FILL  FILL_7__2688_
timestamp 1701859473
transform 1 0 150 0 -1 10150
box -12 -8 32 272
use FILL  FILL_7__2689_
timestamp 1701859473
transform 1 0 370 0 -1 9630
box -12 -8 32 272
use FILL  FILL_7__2690_
timestamp 1701859473
transform 1 0 370 0 1 9110
box -12 -8 32 272
use FILL  FILL_7__2691_
timestamp 1701859473
transform 1 0 2830 0 1 8590
box -12 -8 32 272
use FILL  FILL_7__2692_
timestamp 1701859473
transform 1 0 2590 0 1 8590
box -12 -8 32 272
use FILL  FILL_7__2693_
timestamp 1701859473
transform -1 0 1250 0 -1 9630
box -12 -8 32 272
use FILL  FILL_7__2695_
timestamp 1701859473
transform 1 0 150 0 1 9630
box -12 -8 32 272
use FILL  FILL_7__2696_
timestamp 1701859473
transform -1 0 630 0 -1 10150
box -12 -8 32 272
use FILL  FILL_7__2697_
timestamp 1701859473
transform 1 0 370 0 -1 10150
box -12 -8 32 272
use FILL  FILL_7__2698_
timestamp 1701859473
transform 1 0 390 0 1 9630
box -12 -8 32 272
use FILL  FILL_7__2699_
timestamp 1701859473
transform 1 0 610 0 -1 9630
box -12 -8 32 272
use FILL  FILL_7__2700_
timestamp 1701859473
transform 1 0 630 0 1 9630
box -12 -8 32 272
use FILL  FILL_7__2702_
timestamp 1701859473
transform 1 0 3570 0 1 8590
box -12 -8 32 272
use FILL  FILL_7__2703_
timestamp 1701859473
transform -1 0 3110 0 1 8590
box -12 -8 32 272
use FILL  FILL_7__2704_
timestamp 1701859473
transform -1 0 1590 0 1 9630
box -12 -8 32 272
use FILL  FILL_7__2705_
timestamp 1701859473
transform 1 0 1330 0 1 9630
box -12 -8 32 272
use FILL  FILL_7__2706_
timestamp 1701859473
transform 1 0 350 0 1 10150
box -12 -8 32 272
use FILL  FILL_7__2707_
timestamp 1701859473
transform -1 0 590 0 1 10150
box -12 -8 32 272
use FILL  FILL_7__2709_
timestamp 1701859473
transform -1 0 610 0 -1 10670
box -12 -8 32 272
use FILL  FILL_7__2710_
timestamp 1701859473
transform 1 0 1790 0 1 10150
box -12 -8 32 272
use FILL  FILL_7__2711_
timestamp 1701859473
transform 1 0 2330 0 1 8590
box -12 -8 32 272
use FILL  FILL_7__2712_
timestamp 1701859473
transform -1 0 2110 0 1 8590
box -12 -8 32 272
use FILL  FILL_7__2713_
timestamp 1701859473
transform -1 0 1970 0 -1 9630
box -12 -8 32 272
use FILL  FILL_7__2714_
timestamp 1701859473
transform 1 0 1730 0 -1 10150
box -12 -8 32 272
use FILL  FILL_7__2715_
timestamp 1701859473
transform 1 0 1050 0 1 10150
box -12 -8 32 272
use FILL  FILL_7__2717_
timestamp 1701859473
transform 1 0 1550 0 1 10150
box -12 -8 32 272
use FILL  FILL_7__2718_
timestamp 1701859473
transform -1 0 10130 0 1 4950
box -12 -8 32 272
use FILL  FILL_7__2719_
timestamp 1701859473
transform -1 0 9890 0 1 4950
box -12 -8 32 272
use FILL  FILL_7__2720_
timestamp 1701859473
transform -1 0 4670 0 1 4950
box -12 -8 32 272
use FILL  FILL_7__2721_
timestamp 1701859473
transform -1 0 7430 0 -1 2350
box -12 -8 32 272
use FILL  FILL_7__2722_
timestamp 1701859473
transform 1 0 10070 0 -1 790
box -12 -8 32 272
use FILL  FILL_7__2724_
timestamp 1701859473
transform -1 0 7190 0 -1 2350
box -12 -8 32 272
use FILL  FILL_7__2725_
timestamp 1701859473
transform 1 0 7050 0 1 3390
box -12 -8 32 272
use FILL  FILL_7__2726_
timestamp 1701859473
transform -1 0 7290 0 1 3390
box -12 -8 32 272
use FILL  FILL_7__2727_
timestamp 1701859473
transform -1 0 5510 0 1 3390
box -12 -8 32 272
use FILL  FILL_7__2728_
timestamp 1701859473
transform -1 0 5730 0 1 3390
box -12 -8 32 272
use FILL  FILL_7__2729_
timestamp 1701859473
transform -1 0 6830 0 -1 3910
box -12 -8 32 272
use FILL  FILL_7__2731_
timestamp 1701859473
transform 1 0 9350 0 1 1830
box -12 -8 32 272
use FILL  FILL_7__2732_
timestamp 1701859473
transform 1 0 7790 0 1 1830
box -12 -8 32 272
use FILL  FILL_7__2733_
timestamp 1701859473
transform 1 0 8670 0 1 2350
box -12 -8 32 272
use FILL  FILL_7__2734_
timestamp 1701859473
transform 1 0 7250 0 -1 5470
box -12 -8 32 272
use FILL  FILL_7__2735_
timestamp 1701859473
transform 1 0 7330 0 -1 2870
box -12 -8 32 272
use FILL  FILL_7__2736_
timestamp 1701859473
transform -1 0 7610 0 1 1310
box -12 -8 32 272
use FILL  FILL_7__2738_
timestamp 1701859473
transform -1 0 8050 0 -1 2870
box -12 -8 32 272
use FILL  FILL_7__2739_
timestamp 1701859473
transform -1 0 7870 0 1 2870
box -12 -8 32 272
use FILL  FILL_7__2740_
timestamp 1701859473
transform -1 0 6650 0 -1 1830
box -12 -8 32 272
use FILL  FILL_7__2741_
timestamp 1701859473
transform 1 0 6850 0 -1 1830
box -12 -8 32 272
use FILL  FILL_7__2742_
timestamp 1701859473
transform -1 0 8290 0 -1 2870
box -12 -8 32 272
use FILL  FILL_7__2743_
timestamp 1701859473
transform -1 0 8310 0 1 2870
box -12 -8 32 272
use FILL  FILL_7__2744_
timestamp 1701859473
transform -1 0 7430 0 -1 270
box -12 -8 32 272
use FILL  FILL_7__2746_
timestamp 1701859473
transform 1 0 8050 0 1 2870
box -12 -8 32 272
use FILL  FILL_7__2747_
timestamp 1701859473
transform -1 0 7850 0 -1 2350
box -12 -8 32 272
use FILL  FILL_7__2748_
timestamp 1701859473
transform 1 0 8030 0 -1 2350
box -12 -8 32 272
use FILL  FILL_7__2749_
timestamp 1701859473
transform 1 0 5990 0 1 1830
box -12 -8 32 272
use FILL  FILL_7__2750_
timestamp 1701859473
transform -1 0 6750 0 -1 1310
box -12 -8 32 272
use FILL  FILL_7__2751_
timestamp 1701859473
transform -1 0 6470 0 1 1830
box -12 -8 32 272
use FILL  FILL_7__2753_
timestamp 1701859473
transform -1 0 7570 0 1 2350
box -12 -8 32 272
use FILL  FILL_7__2754_
timestamp 1701859473
transform 1 0 8910 0 -1 4950
box -12 -8 32 272
use FILL  FILL_7__2755_
timestamp 1701859473
transform 1 0 9810 0 1 790
box -12 -8 32 272
use FILL  FILL_7__2756_
timestamp 1701859473
transform -1 0 10050 0 1 790
box -12 -8 32 272
use FILL  FILL_7__2757_
timestamp 1701859473
transform 1 0 10750 0 -1 2870
box -12 -8 32 272
use FILL  FILL_7__2758_
timestamp 1701859473
transform -1 0 9250 0 -1 2870
box -12 -8 32 272
use FILL  FILL_7__2760_
timestamp 1701859473
transform 1 0 10510 0 -1 790
box -12 -8 32 272
use FILL  FILL_7__2761_
timestamp 1701859473
transform 1 0 10270 0 -1 790
box -12 -8 32 272
use FILL  FILL_7__2762_
timestamp 1701859473
transform -1 0 10950 0 -1 1830
box -12 -8 32 272
use FILL  FILL_7__2763_
timestamp 1701859473
transform 1 0 6690 0 1 1830
box -12 -8 32 272
use FILL  FILL_7__2764_
timestamp 1701859473
transform -1 0 6950 0 1 1830
box -12 -8 32 272
use FILL  FILL_7__2765_
timestamp 1701859473
transform -1 0 10250 0 1 1830
box -12 -8 32 272
use FILL  FILL_7__2766_
timestamp 1701859473
transform -1 0 10070 0 -1 1830
box -12 -8 32 272
use FILL  FILL_7__2768_
timestamp 1701859473
transform -1 0 10470 0 1 1830
box -12 -8 32 272
use FILL  FILL_7__2769_
timestamp 1701859473
transform -1 0 10930 0 1 2350
box -12 -8 32 272
use FILL  FILL_7__2770_
timestamp 1701859473
transform -1 0 10710 0 -1 1830
box -12 -8 32 272
use FILL  FILL_7__2771_
timestamp 1701859473
transform 1 0 11130 0 1 2350
box -12 -8 32 272
use FILL  FILL_7__2772_
timestamp 1701859473
transform -1 0 10790 0 1 4950
box -12 -8 32 272
use FILL  FILL_7__2773_
timestamp 1701859473
transform 1 0 10530 0 -1 3910
box -12 -8 32 272
use FILL  FILL_7__2775_
timestamp 1701859473
transform -1 0 9190 0 -1 1310
box -12 -8 32 272
use FILL  FILL_7__2776_
timestamp 1701859473
transform 1 0 10730 0 -1 790
box -12 -8 32 272
use FILL  FILL_7__2777_
timestamp 1701859473
transform -1 0 8490 0 -1 270
box -12 -8 32 272
use FILL  FILL_7__2778_
timestamp 1701859473
transform 1 0 11030 0 1 270
box -12 -8 32 272
use FILL  FILL_7__2779_
timestamp 1701859473
transform 1 0 9110 0 -1 1830
box -12 -8 32 272
use FILL  FILL_7__2780_
timestamp 1701859473
transform -1 0 10130 0 1 1310
box -12 -8 32 272
use FILL  FILL_7__2782_
timestamp 1701859473
transform 1 0 8890 0 1 1830
box -12 -8 32 272
use FILL  FILL_7__2783_
timestamp 1701859473
transform 1 0 8450 0 -1 1310
box -12 -8 32 272
use FILL  FILL_7__2784_
timestamp 1701859473
transform 1 0 8690 0 -1 1310
box -12 -8 32 272
use FILL  FILL_7__2785_
timestamp 1701859473
transform 1 0 8910 0 -1 1830
box -12 -8 32 272
use FILL  FILL_7__2786_
timestamp 1701859473
transform -1 0 9390 0 -1 1310
box -12 -8 32 272
use FILL  FILL_7__2787_
timestamp 1701859473
transform -1 0 9590 0 -1 1830
box -12 -8 32 272
use FILL  FILL_7__2789_
timestamp 1701859473
transform 1 0 10350 0 1 1310
box -12 -8 32 272
use FILL  FILL_7__2790_
timestamp 1701859473
transform -1 0 10150 0 -1 2350
box -12 -8 32 272
use FILL  FILL_7__2791_
timestamp 1701859473
transform 1 0 9910 0 -1 2350
box -12 -8 32 272
use FILL  FILL_7__2792_
timestamp 1701859473
transform -1 0 10370 0 -1 2350
box -12 -8 32 272
use FILL  FILL_7__2793_
timestamp 1701859473
transform -1 0 10610 0 -1 2350
box -12 -8 32 272
use FILL  FILL_7__2794_
timestamp 1701859473
transform -1 0 11030 0 -1 2350
box -12 -8 32 272
use FILL  FILL_7__2795_
timestamp 1701859473
transform -1 0 10990 0 -1 2870
box -12 -8 32 272
use FILL  FILL_7__2797_
timestamp 1701859473
transform -1 0 9830 0 -1 1830
box -12 -8 32 272
use FILL  FILL_7__2798_
timestamp 1701859473
transform -1 0 10710 0 1 2350
box -12 -8 32 272
use FILL  FILL_7__2799_
timestamp 1701859473
transform 1 0 10490 0 -1 2870
box -12 -8 32 272
use FILL  FILL_7__2800_
timestamp 1701859473
transform -1 0 10510 0 -1 4430
box -12 -8 32 272
use FILL  FILL_7__2801_
timestamp 1701859473
transform -1 0 9470 0 -1 2870
box -12 -8 32 272
use FILL  FILL_7__2802_
timestamp 1701859473
transform -1 0 7330 0 -1 1830
box -12 -8 32 272
use FILL  FILL_7__2804_
timestamp 1701859473
transform -1 0 9590 0 -1 3390
box -12 -8 32 272
use FILL  FILL_7__2805_
timestamp 1701859473
transform -1 0 9890 0 -1 2870
box -12 -8 32 272
use FILL  FILL_7__2806_
timestamp 1701859473
transform 1 0 9650 0 -1 2870
box -12 -8 32 272
use FILL  FILL_7__2807_
timestamp 1701859473
transform 1 0 8990 0 -1 2350
box -12 -8 32 272
use FILL  FILL_7__2808_
timestamp 1701859473
transform 1 0 8750 0 -1 2350
box -12 -8 32 272
use FILL  FILL_7__2809_
timestamp 1701859473
transform 1 0 10470 0 1 2350
box -12 -8 32 272
use FILL  FILL_7__2811_
timestamp 1701859473
transform 1 0 5030 0 -1 4430
box -12 -8 32 272
use FILL  FILL_7__2812_
timestamp 1701859473
transform -1 0 8990 0 1 4950
box -12 -8 32 272
use FILL  FILL_7__2813_
timestamp 1701859473
transform 1 0 9090 0 1 3390
box -12 -8 32 272
use FILL  FILL_7__2814_
timestamp 1701859473
transform -1 0 8910 0 -1 4430
box -12 -8 32 272
use FILL  FILL_7__2815_
timestamp 1701859473
transform -1 0 8690 0 1 3910
box -12 -8 32 272
use FILL  FILL_7__2816_
timestamp 1701859473
transform -1 0 8310 0 1 4950
box -12 -8 32 272
use FILL  FILL_7__2818_
timestamp 1701859473
transform 1 0 8450 0 -1 4430
box -12 -8 32 272
use FILL  FILL_7__2819_
timestamp 1701859473
transform 1 0 8650 0 -1 4430
box -12 -8 32 272
use FILL  FILL_7__2820_
timestamp 1701859473
transform -1 0 9610 0 1 2350
box -12 -8 32 272
use FILL  FILL_7__2821_
timestamp 1701859473
transform 1 0 9130 0 1 2350
box -12 -8 32 272
use FILL  FILL_7__2822_
timestamp 1701859473
transform -1 0 9130 0 1 1830
box -12 -8 32 272
use FILL  FILL_7__2823_
timestamp 1701859473
transform -1 0 8910 0 1 2350
box -12 -8 32 272
use FILL  FILL_7__2824_
timestamp 1701859473
transform 1 0 10030 0 -1 3390
box -12 -8 32 272
use FILL  FILL_7__2826_
timestamp 1701859473
transform 1 0 9610 0 1 790
box -12 -8 32 272
use FILL  FILL_7__2827_
timestamp 1701859473
transform -1 0 9350 0 -1 1830
box -12 -8 32 272
use FILL  FILL_7__2828_
timestamp 1701859473
transform 1 0 7070 0 -1 1830
box -12 -8 32 272
use FILL  FILL_7__2829_
timestamp 1701859473
transform -1 0 10090 0 1 2870
box -12 -8 32 272
use FILL  FILL_7__2830_
timestamp 1701859473
transform 1 0 8390 0 -1 3390
box -12 -8 32 272
use FILL  FILL_7__2831_
timestamp 1701859473
transform 1 0 8430 0 1 3910
box -12 -8 32 272
use FILL  FILL_7__2833_
timestamp 1701859473
transform -1 0 9350 0 -1 3390
box -12 -8 32 272
use FILL  FILL_7__2834_
timestamp 1701859473
transform -1 0 9110 0 -1 3390
box -12 -8 32 272
use FILL  FILL_7__2835_
timestamp 1701859473
transform -1 0 9410 0 1 790
box -12 -8 32 272
use FILL  FILL_7__2836_
timestamp 1701859473
transform 1 0 8990 0 1 1310
box -12 -8 32 272
use FILL  FILL_7__2837_
timestamp 1701859473
transform -1 0 9670 0 1 1310
box -12 -8 32 272
use FILL  FILL_7__2838_
timestamp 1701859473
transform -1 0 9790 0 1 3390
box -12 -8 32 272
use FILL  FILL_7__2840_
timestamp 1701859473
transform 1 0 9150 0 -1 270
box -12 -8 32 272
use FILL  FILL_7__2841_
timestamp 1701859473
transform -1 0 8950 0 -1 270
box -12 -8 32 272
use FILL  FILL_7__2842_
timestamp 1701859473
transform 1 0 9370 0 -1 270
box -12 -8 32 272
use FILL  FILL_7__2843_
timestamp 1701859473
transform 1 0 9610 0 -1 270
box -12 -8 32 272
use FILL  FILL_7__2844_
timestamp 1701859473
transform 1 0 9410 0 1 270
box -12 -8 32 272
use FILL  FILL_7__2845_
timestamp 1701859473
transform -1 0 10090 0 1 270
box -12 -8 32 272
use FILL  FILL_7__2846_
timestamp 1701859473
transform 1 0 9830 0 1 270
box -12 -8 32 272
use FILL  FILL_7__2848_
timestamp 1701859473
transform -1 0 10710 0 -1 1310
box -12 -8 32 272
use FILL  FILL_7__2849_
timestamp 1701859473
transform -1 0 11050 0 1 1310
box -12 -8 32 272
use FILL  FILL_7__2850_
timestamp 1701859473
transform -1 0 11190 0 -1 1830
box -12 -8 32 272
use FILL  FILL_7__2851_
timestamp 1701859473
transform 1 0 10790 0 -1 3910
box -12 -8 32 272
use FILL  FILL_7__2852_
timestamp 1701859473
transform -1 0 8990 0 1 270
box -12 -8 32 272
use FILL  FILL_7__2853_
timestamp 1701859473
transform -1 0 9210 0 1 270
box -12 -8 32 272
use FILL  FILL_7__2855_
timestamp 1701859473
transform -1 0 9910 0 1 1310
box -12 -8 32 272
use FILL  FILL_7__2856_
timestamp 1701859473
transform -1 0 10570 0 1 1310
box -12 -8 32 272
use FILL  FILL_7__2857_
timestamp 1701859473
transform -1 0 10810 0 1 1310
box -12 -8 32 272
use FILL  FILL_7__2858_
timestamp 1701859473
transform -1 0 11170 0 1 1830
box -12 -8 32 272
use FILL  FILL_7__2859_
timestamp 1701859473
transform 1 0 11030 0 -1 3910
box -12 -8 32 272
use FILL  FILL_7__2860_
timestamp 1701859473
transform 1 0 10950 0 -1 3390
box -12 -8 32 272
use FILL  FILL_7__2862_
timestamp 1701859473
transform 1 0 8690 0 -1 270
box -12 -8 32 272
use FILL  FILL_7__2863_
timestamp 1701859473
transform -1 0 10330 0 1 270
box -12 -8 32 272
use FILL  FILL_7__2864_
timestamp 1701859473
transform 1 0 10570 0 1 270
box -12 -8 32 272
use FILL  FILL_7__2865_
timestamp 1701859473
transform -1 0 10810 0 1 270
box -12 -8 32 272
use FILL  FILL_7__2866_
timestamp 1701859473
transform -1 0 11190 0 -1 790
box -12 -8 32 272
use FILL  FILL_7__2867_
timestamp 1701859473
transform 1 0 11150 0 -1 3390
box -12 -8 32 272
use FILL  FILL_7__2869_
timestamp 1701859473
transform 1 0 10250 0 1 790
box -12 -8 32 272
use FILL  FILL_7__2870_
timestamp 1701859473
transform -1 0 10470 0 1 790
box -12 -8 32 272
use FILL  FILL_7__2871_
timestamp 1701859473
transform -1 0 10910 0 1 790
box -12 -8 32 272
use FILL  FILL_7__2872_
timestamp 1701859473
transform -1 0 11250 0 1 1310
box -12 -8 32 272
use FILL  FILL_7__2873_
timestamp 1701859473
transform -1 0 10030 0 1 3390
box -12 -8 32 272
use FILL  FILL_7__2874_
timestamp 1701859473
transform -1 0 10270 0 1 3390
box -12 -8 32 272
use FILL  FILL_7__2875_
timestamp 1701859473
transform -1 0 10850 0 -1 4950
box -12 -8 32 272
use FILL  FILL_7__2877_
timestamp 1701859473
transform 1 0 9990 0 1 1830
box -12 -8 32 272
use FILL  FILL_7__2878_
timestamp 1701859473
transform 1 0 9810 0 -1 1310
box -12 -8 32 272
use FILL  FILL_7__2879_
timestamp 1701859473
transform -1 0 10050 0 -1 1310
box -12 -8 32 272
use FILL  FILL_7__2880_
timestamp 1701859473
transform 1 0 9550 0 1 1830
box -12 -8 32 272
use FILL  FILL_7__2881_
timestamp 1701859473
transform 1 0 10930 0 -1 790
box -12 -8 32 272
use FILL  FILL_7__2882_
timestamp 1701859473
transform -1 0 9610 0 -1 1310
box -12 -8 32 272
use FILL  FILL_7__2884_
timestamp 1701859473
transform 1 0 11150 0 -1 1310
box -12 -8 32 272
use FILL  FILL_7__2885_
timestamp 1701859473
transform -1 0 10930 0 -1 1310
box -12 -8 32 272
use FILL  FILL_7__2886_
timestamp 1701859473
transform 1 0 10690 0 1 1830
box -12 -8 32 272
use FILL  FILL_7__2887_
timestamp 1701859473
transform 1 0 10250 0 -1 4430
box -12 -8 32 272
use FILL  FILL_7__2888_
timestamp 1701859473
transform -1 0 4070 0 1 5470
box -12 -8 32 272
use FILL  FILL_7__2889_
timestamp 1701859473
transform 1 0 6190 0 1 2350
box -12 -8 32 272
use FILL  FILL_7__2891_
timestamp 1701859473
transform -1 0 8270 0 1 5990
box -12 -8 32 272
use FILL  FILL_7__2892_
timestamp 1701859473
transform 1 0 7490 0 -1 5470
box -12 -8 32 272
use FILL  FILL_7__2893_
timestamp 1701859473
transform 1 0 7310 0 1 5470
box -12 -8 32 272
use FILL  FILL_7__2894_
timestamp 1701859473
transform 1 0 6590 0 -1 6510
box -12 -8 32 272
use FILL  FILL_7__2895_
timestamp 1701859473
transform 1 0 6730 0 1 6510
box -12 -8 32 272
use FILL  FILL_7__2896_
timestamp 1701859473
transform -1 0 7990 0 -1 5470
box -12 -8 32 272
use FILL  FILL_7__2898_
timestamp 1701859473
transform 1 0 7310 0 -1 6510
box -12 -8 32 272
use FILL  FILL_7__2899_
timestamp 1701859473
transform 1 0 6830 0 -1 6510
box -12 -8 32 272
use FILL  FILL_7__2900_
timestamp 1701859473
transform -1 0 6370 0 -1 6510
box -12 -8 32 272
use FILL  FILL_7__2901_
timestamp 1701859473
transform 1 0 6110 0 -1 6510
box -12 -8 32 272
use FILL  FILL_7__2902_
timestamp 1701859473
transform -1 0 8030 0 1 5990
box -12 -8 32 272
use FILL  FILL_7__2903_
timestamp 1701859473
transform 1 0 7310 0 1 5990
box -12 -8 32 272
use FILL  FILL_7__2904_
timestamp 1701859473
transform 1 0 8430 0 -1 5470
box -12 -8 32 272
use FILL  FILL_7__2906_
timestamp 1701859473
transform 1 0 8190 0 -1 5990
box -12 -8 32 272
use FILL  FILL_7__2907_
timestamp 1701859473
transform -1 0 7970 0 -1 5990
box -12 -8 32 272
use FILL  FILL_7__2908_
timestamp 1701859473
transform -1 0 8290 0 -1 4950
box -12 -8 32 272
use FILL  FILL_7__2909_
timestamp 1701859473
transform 1 0 3430 0 -1 4430
box -12 -8 32 272
use FILL  FILL_7__2910_
timestamp 1701859473
transform -1 0 6590 0 -1 4430
box -12 -8 32 272
use FILL  FILL_7__2911_
timestamp 1701859473
transform -1 0 6930 0 1 4430
box -12 -8 32 272
use FILL  FILL_7__2913_
timestamp 1701859473
transform -1 0 6890 0 -1 4950
box -12 -8 32 272
use FILL  FILL_7__2914_
timestamp 1701859473
transform 1 0 7150 0 -1 8070
box -12 -8 32 272
use FILL  FILL_7__2915_
timestamp 1701859473
transform 1 0 7270 0 -1 5990
box -12 -8 32 272
use FILL  FILL_7__2916_
timestamp 1701859473
transform 1 0 7030 0 -1 5990
box -12 -8 32 272
use FILL  FILL_7__2917_
timestamp 1701859473
transform -1 0 6410 0 -1 5990
box -12 -8 32 272
use FILL  FILL_7__2918_
timestamp 1701859473
transform 1 0 6330 0 1 5470
box -12 -8 32 272
use FILL  FILL_7__2920_
timestamp 1701859473
transform 1 0 6010 0 1 4950
box -12 -8 32 272
use FILL  FILL_7__2921_
timestamp 1701859473
transform -1 0 7470 0 -1 3910
box -12 -8 32 272
use FILL  FILL_7__2922_
timestamp 1701859473
transform -1 0 7510 0 1 3910
box -12 -8 32 272
use FILL  FILL_7__2923_
timestamp 1701859473
transform -1 0 6830 0 -1 4430
box -12 -8 32 272
use FILL  FILL_7__2924_
timestamp 1701859473
transform 1 0 6450 0 1 4950
box -12 -8 32 272
use FILL  FILL_7__2925_
timestamp 1701859473
transform 1 0 7350 0 1 7550
box -12 -8 32 272
use FILL  FILL_7__2926_
timestamp 1701859473
transform -1 0 7590 0 1 4430
box -12 -8 32 272
use FILL  FILL_7__2928_
timestamp 1701859473
transform 1 0 7110 0 -1 4950
box -12 -8 32 272
use FILL  FILL_7__2929_
timestamp 1701859473
transform -1 0 6690 0 1 4950
box -12 -8 32 272
use FILL  FILL_7__2930_
timestamp 1701859473
transform 1 0 6230 0 1 1830
box -12 -8 32 272
use FILL  FILL_7__2931_
timestamp 1701859473
transform 1 0 7110 0 -1 2870
box -12 -8 32 272
use FILL  FILL_7__2932_
timestamp 1701859473
transform 1 0 5270 0 -1 4430
box -12 -8 32 272
use FILL  FILL_7__2933_
timestamp 1701859473
transform 1 0 5470 0 -1 4430
box -12 -8 32 272
use FILL  FILL_7__2935_
timestamp 1701859473
transform 1 0 6530 0 1 6510
box -12 -8 32 272
use FILL  FILL_7__2936_
timestamp 1701859473
transform 1 0 6410 0 -1 4950
box -12 -8 32 272
use FILL  FILL_7__2937_
timestamp 1701859473
transform 1 0 6630 0 -1 4950
box -12 -8 32 272
use FILL  FILL_7__2938_
timestamp 1701859473
transform 1 0 5110 0 1 4950
box -12 -8 32 272
use FILL  FILL_7__2939_
timestamp 1701859473
transform 1 0 4890 0 1 4950
box -12 -8 32 272
use FILL  FILL_7__2940_
timestamp 1701859473
transform -1 0 5950 0 -1 5470
box -12 -8 32 272
use FILL  FILL_7__2942_
timestamp 1701859473
transform -1 0 9410 0 1 4430
box -12 -8 32 272
use FILL  FILL_7__2943_
timestamp 1701859473
transform 1 0 6370 0 -1 4430
box -12 -8 32 272
use FILL  FILL_7__2944_
timestamp 1701859473
transform -1 0 6390 0 1 3910
box -12 -8 32 272
use FILL  FILL_7__2945_
timestamp 1701859473
transform -1 0 6470 0 1 4430
box -12 -8 32 272
use FILL  FILL_7__2946_
timestamp 1701859473
transform 1 0 6230 0 1 4430
box -12 -8 32 272
use FILL  FILL_7__2947_
timestamp 1701859473
transform -1 0 6630 0 -1 5990
box -12 -8 32 272
use FILL  FILL_7__2949_
timestamp 1701859473
transform -1 0 5990 0 -1 5990
box -12 -8 32 272
use FILL  FILL_7__2950_
timestamp 1701859473
transform 1 0 5850 0 1 5470
box -12 -8 32 272
use FILL  FILL_7__2951_
timestamp 1701859473
transform -1 0 6110 0 1 5470
box -12 -8 32 272
use FILL  FILL_7__2952_
timestamp 1701859473
transform -1 0 6190 0 -1 4950
box -12 -8 32 272
use FILL  FILL_7__2953_
timestamp 1701859473
transform -1 0 4470 0 1 4950
box -12 -8 32 272
use FILL  FILL_7__2954_
timestamp 1701859473
transform -1 0 6730 0 1 4430
box -12 -8 32 272
use FILL  FILL_7__2955_
timestamp 1701859473
transform -1 0 6010 0 1 4430
box -12 -8 32 272
use FILL  FILL_7__2957_
timestamp 1701859473
transform 1 0 5230 0 -1 4950
box -12 -8 32 272
use FILL  FILL_7__2958_
timestamp 1701859473
transform -1 0 5550 0 1 4430
box -12 -8 32 272
use FILL  FILL_7__2959_
timestamp 1701859473
transform 1 0 7050 0 -1 5470
box -12 -8 32 272
use FILL  FILL_7__2960_
timestamp 1701859473
transform -1 0 6590 0 1 5470
box -12 -8 32 272
use FILL  FILL_7__2961_
timestamp 1701859473
transform 1 0 6350 0 -1 5470
box -12 -8 32 272
use FILL  FILL_7__2962_
timestamp 1701859473
transform -1 0 6610 0 -1 5470
box -12 -8 32 272
use FILL  FILL_7__2964_
timestamp 1701859473
transform -1 0 5490 0 -1 4950
box -12 -8 32 272
use FILL  FILL_7__2965_
timestamp 1701859473
transform 1 0 4990 0 -1 4950
box -12 -8 32 272
use FILL  FILL_7__2966_
timestamp 1701859473
transform -1 0 6450 0 1 2350
box -12 -8 32 272
use FILL  FILL_7__2967_
timestamp 1701859473
transform 1 0 7710 0 1 3910
box -12 -8 32 272
use FILL  FILL_7__2968_
timestamp 1701859473
transform -1 0 7030 0 -1 3910
box -12 -8 32 272
use FILL  FILL_7__2969_
timestamp 1701859473
transform -1 0 7250 0 -1 3910
box -12 -8 32 272
use FILL  FILL_7__2971_
timestamp 1701859473
transform -1 0 6810 0 1 3910
box -12 -8 32 272
use FILL  FILL_7__2972_
timestamp 1701859473
transform 1 0 7030 0 1 3910
box -12 -8 32 272
use FILL  FILL_7__2973_
timestamp 1701859473
transform -1 0 7150 0 1 4430
box -12 -8 32 272
use FILL  FILL_7__2974_
timestamp 1701859473
transform 1 0 7050 0 -1 4430
box -12 -8 32 272
use FILL  FILL_7__2975_
timestamp 1701859473
transform -1 0 7810 0 -1 4430
box -12 -8 32 272
use FILL  FILL_7__2976_
timestamp 1701859473
transform -1 0 7570 0 -1 4430
box -12 -8 32 272
use FILL  FILL_7__2977_
timestamp 1701859473
transform 1 0 7290 0 -1 4430
box -12 -8 32 272
use FILL  FILL_7__2979_
timestamp 1701859473
transform -1 0 3690 0 -1 4950
box -12 -8 32 272
use FILL  FILL_7__2980_
timestamp 1701859473
transform -1 0 3070 0 1 7550
box -12 -8 32 272
use FILL  FILL_7__2981_
timestamp 1701859473
transform 1 0 3590 0 1 4950
box -12 -8 32 272
use FILL  FILL_7__2982_
timestamp 1701859473
transform 1 0 9650 0 1 6510
box -12 -8 32 272
use FILL  FILL_7__2983_
timestamp 1701859473
transform 1 0 1970 0 1 4430
box -12 -8 32 272
use FILL  FILL_7__2984_
timestamp 1701859473
transform -1 0 3590 0 -1 3910
box -12 -8 32 272
use FILL  FILL_7__2986_
timestamp 1701859473
transform -1 0 5950 0 -1 4430
box -12 -8 32 272
use FILL  FILL_7__2987_
timestamp 1701859473
transform -1 0 5770 0 1 4430
box -12 -8 32 272
use FILL  FILL_7__2988_
timestamp 1701859473
transform 1 0 9430 0 1 6510
box -12 -8 32 272
use FILL  FILL_7__2989_
timestamp 1701859473
transform 1 0 6050 0 1 6510
box -12 -8 32 272
use FILL  FILL_7__2990_
timestamp 1701859473
transform -1 0 6310 0 1 6510
box -12 -8 32 272
use FILL  FILL_7__2991_
timestamp 1701859473
transform 1 0 7210 0 1 6510
box -12 -8 32 272
use FILL  FILL_7__2993_
timestamp 1701859473
transform 1 0 9930 0 1 7030
box -12 -8 32 272
use FILL  FILL_7__2994_
timestamp 1701859473
transform -1 0 10850 0 -1 7550
box -12 -8 32 272
use FILL  FILL_7__2995_
timestamp 1701859473
transform -1 0 7650 0 -1 7550
box -12 -8 32 272
use FILL  FILL_7__2996_
timestamp 1701859473
transform 1 0 7550 0 1 7550
box -12 -8 32 272
use FILL  FILL_7__2997_
timestamp 1701859473
transform -1 0 7430 0 -1 7550
box -12 -8 32 272
use FILL  FILL_7__2998_
timestamp 1701859473
transform -1 0 6490 0 -1 7550
box -12 -8 32 272
use FILL  FILL_7__3000_
timestamp 1701859473
transform -1 0 6050 0 -1 7550
box -12 -8 32 272
use FILL  FILL_7__3001_
timestamp 1701859473
transform -1 0 5830 0 -1 7550
box -12 -8 32 272
use FILL  FILL_7__3002_
timestamp 1701859473
transform -1 0 6250 0 -1 7550
box -12 -8 32 272
use FILL  FILL_7__3003_
timestamp 1701859473
transform -1 0 6430 0 1 7550
box -12 -8 32 272
use FILL  FILL_7__3004_
timestamp 1701859473
transform 1 0 8230 0 1 7550
box -12 -8 32 272
use FILL  FILL_7__3005_
timestamp 1701859473
transform 1 0 11050 0 -1 7550
box -12 -8 32 272
use FILL  FILL_7__3006_
timestamp 1701859473
transform -1 0 10530 0 1 7550
box -12 -8 32 272
use FILL  FILL_7__3008_
timestamp 1701859473
transform -1 0 6610 0 1 7030
box -12 -8 32 272
use FILL  FILL_7__3009_
timestamp 1701859473
transform -1 0 6010 0 -1 7030
box -12 -8 32 272
use FILL  FILL_7__3010_
timestamp 1701859473
transform 1 0 6230 0 -1 7030
box -12 -8 32 272
use FILL  FILL_7__3011_
timestamp 1701859473
transform 1 0 6810 0 1 7030
box -12 -8 32 272
use FILL  FILL_7__3012_
timestamp 1701859473
transform -1 0 7930 0 -1 7030
box -12 -8 32 272
use FILL  FILL_7__3013_
timestamp 1701859473
transform 1 0 8370 0 -1 7030
box -12 -8 32 272
use FILL  FILL_7__3015_
timestamp 1701859473
transform -1 0 6450 0 -1 7030
box -12 -8 32 272
use FILL  FILL_7__3016_
timestamp 1701859473
transform -1 0 7330 0 1 7030
box -12 -8 32 272
use FILL  FILL_7__3017_
timestamp 1701859473
transform 1 0 6670 0 -1 7030
box -12 -8 32 272
use FILL  FILL_7__3018_
timestamp 1701859473
transform -1 0 6970 0 -1 7030
box -12 -8 32 272
use FILL  FILL_7__3019_
timestamp 1701859473
transform -1 0 7210 0 -1 7030
box -12 -8 32 272
use FILL  FILL_7__3020_
timestamp 1701859473
transform 1 0 8370 0 1 7030
box -12 -8 32 272
use FILL  FILL_7__3022_
timestamp 1701859473
transform 1 0 9610 0 -1 8070
box -12 -8 32 272
use FILL  FILL_7__3023_
timestamp 1701859473
transform -1 0 5830 0 1 6510
box -12 -8 32 272
use FILL  FILL_7__3024_
timestamp 1701859473
transform 1 0 5570 0 1 6510
box -12 -8 32 272
use FILL  FILL_7__3025_
timestamp 1701859473
transform -1 0 5590 0 -1 6510
box -12 -8 32 272
use FILL  FILL_7__3026_
timestamp 1701859473
transform 1 0 11010 0 -1 5990
box -12 -8 32 272
use FILL  FILL_7__3027_
timestamp 1701859473
transform -1 0 11250 0 -1 5990
box -12 -8 32 272
use FILL  FILL_7__3029_
timestamp 1701859473
transform -1 0 7190 0 -1 7550
box -12 -8 32 272
use FILL  FILL_7__3030_
timestamp 1701859473
transform -1 0 8170 0 -1 7030
box -12 -8 32 272
use FILL  FILL_7__3031_
timestamp 1701859473
transform 1 0 8150 0 1 7030
box -12 -8 32 272
use FILL  FILL_7__3032_
timestamp 1701859473
transform 1 0 7770 0 1 7550
box -12 -8 32 272
use FILL  FILL_7__3033_
timestamp 1701859473
transform -1 0 6850 0 1 8070
box -12 -8 32 272
use FILL  FILL_7__3034_
timestamp 1701859473
transform -1 0 7830 0 -1 8070
box -12 -8 32 272
use FILL  FILL_7__3035_
timestamp 1701859473
transform 1 0 7570 0 -1 8070
box -12 -8 32 272
use FILL  FILL_7__3037_
timestamp 1701859473
transform -1 0 6610 0 1 8070
box -12 -8 32 272
use FILL  FILL_7__3038_
timestamp 1701859473
transform -1 0 7230 0 1 8070
box -12 -8 32 272
use FILL  FILL_7__3039_
timestamp 1701859473
transform 1 0 7450 0 1 8070
box -12 -8 32 272
use FILL  FILL_7__3040_
timestamp 1701859473
transform 1 0 9790 0 1 7550
box -12 -8 32 272
use FILL  FILL_7__3041_
timestamp 1701859473
transform -1 0 9650 0 -1 6510
box -12 -8 32 272
use FILL  FILL_7__3042_
timestamp 1701859473
transform 1 0 7350 0 -1 8070
box -12 -8 32 272
use FILL  FILL_7__3044_
timestamp 1701859473
transform -1 0 6710 0 -1 7550
box -12 -8 32 272
use FILL  FILL_7__3045_
timestamp 1701859473
transform 1 0 6930 0 -1 7550
box -12 -8 32 272
use FILL  FILL_7__3046_
timestamp 1701859473
transform -1 0 7890 0 1 6510
box -12 -8 32 272
use FILL  FILL_7__3047_
timestamp 1701859473
transform 1 0 9230 0 1 6510
box -12 -8 32 272
use FILL  FILL_7__3048_
timestamp 1701859473
transform 1 0 9850 0 -1 6510
box -12 -8 32 272
use FILL  FILL_7__3049_
timestamp 1701859473
transform -1 0 6930 0 1 7550
box -12 -8 32 272
use FILL  FILL_7__3051_
timestamp 1701859473
transform -1 0 7890 0 1 7030
box -12 -8 32 272
use FILL  FILL_7__3052_
timestamp 1701859473
transform 1 0 7590 0 1 7030
box -12 -8 32 272
use FILL  FILL_7__3053_
timestamp 1701859473
transform 1 0 7430 0 -1 7030
box -12 -8 32 272
use FILL  FILL_7__3054_
timestamp 1701859473
transform -1 0 7690 0 -1 7030
box -12 -8 32 272
use FILL  FILL_7__3055_
timestamp 1701859473
transform 1 0 8110 0 1 6510
box -12 -8 32 272
use FILL  FILL_7__3056_
timestamp 1701859473
transform -1 0 9630 0 1 5470
box -12 -8 32 272
use FILL  FILL_7__3057_
timestamp 1701859473
transform -1 0 9390 0 1 5470
box -12 -8 32 272
use FILL  FILL_7__3059_
timestamp 1701859473
transform -1 0 8690 0 -1 5990
box -12 -8 32 272
use FILL  FILL_7__3060_
timestamp 1701859473
transform 1 0 9870 0 1 6510
box -12 -8 32 272
use FILL  FILL_7__3061_
timestamp 1701859473
transform 1 0 10110 0 1 6510
box -12 -8 32 272
use FILL  FILL_7__3062_
timestamp 1701859473
transform -1 0 9730 0 -1 7550
box -12 -8 32 272
use FILL  FILL_7__3063_
timestamp 1701859473
transform 1 0 9470 0 -1 7550
box -12 -8 32 272
use FILL  FILL_7__3064_
timestamp 1701859473
transform -1 0 10430 0 -1 7030
box -12 -8 32 272
use FILL  FILL_7__3066_
timestamp 1701859473
transform -1 0 8590 0 -1 7550
box -12 -8 32 272
use FILL  FILL_7__3067_
timestamp 1701859473
transform 1 0 8330 0 -1 7550
box -12 -8 32 272
use FILL  FILL_7__3068_
timestamp 1701859473
transform 1 0 10290 0 -1 5990
box -12 -8 32 272
use FILL  FILL_7__3069_
timestamp 1701859473
transform 1 0 10530 0 -1 5990
box -12 -8 32 272
use FILL  FILL_7__3070_
timestamp 1701859473
transform 1 0 8990 0 -1 7550
box -12 -8 32 272
use FILL  FILL_7__3071_
timestamp 1701859473
transform -1 0 9250 0 -1 7550
box -12 -8 32 272
use FILL  FILL_7__3073_
timestamp 1701859473
transform -1 0 10090 0 1 5990
box -12 -8 32 272
use FILL  FILL_7__3074_
timestamp 1701859473
transform 1 0 8910 0 1 5990
box -12 -8 32 272
use FILL  FILL_7__3075_
timestamp 1701859473
transform 1 0 8910 0 -1 5990
box -12 -8 32 272
use FILL  FILL_7__3076_
timestamp 1701859473
transform 1 0 10810 0 1 6510
box -12 -8 32 272
use FILL  FILL_7__3077_
timestamp 1701859473
transform 1 0 11010 0 1 6510
box -12 -8 32 272
use FILL  FILL_7__3078_
timestamp 1701859473
transform -1 0 8810 0 -1 7030
box -12 -8 32 272
use FILL  FILL_7__3080_
timestamp 1701859473
transform 1 0 11070 0 -1 8590
box -12 -8 32 272
use FILL  FILL_7__3081_
timestamp 1701859473
transform -1 0 11070 0 -1 270
box -12 -8 32 272
use FILL  FILL_7__3082_
timestamp 1701859473
transform 1 0 10170 0 -1 8590
box -12 -8 32 272
use FILL  FILL_7__3083_
timestamp 1701859473
transform -1 0 9950 0 -1 8590
box -12 -8 32 272
use FILL  FILL_7__3084_
timestamp 1701859473
transform -1 0 9130 0 1 7550
box -12 -8 32 272
use FILL  FILL_7__3085_
timestamp 1701859473
transform 1 0 9030 0 1 7030
box -12 -8 32 272
use FILL  FILL_7__3086_
timestamp 1701859473
transform -1 0 10790 0 1 5990
box -12 -8 32 272
use FILL  FILL_7__3088_
timestamp 1701859473
transform 1 0 8350 0 1 8070
box -12 -8 32 272
use FILL  FILL_7__3089_
timestamp 1701859473
transform -1 0 8130 0 1 8070
box -12 -8 32 272
use FILL  FILL_7__3090_
timestamp 1701859473
transform -1 0 11230 0 1 4950
box -12 -8 32 272
use FILL  FILL_7__3091_
timestamp 1701859473
transform 1 0 10970 0 1 4950
box -12 -8 32 272
use FILL  FILL_7__3092_
timestamp 1701859473
transform 1 0 8890 0 -1 5470
box -12 -8 32 272
use FILL  FILL_7__3093_
timestamp 1701859473
transform -1 0 9130 0 -1 5470
box -12 -8 32 272
use FILL  FILL_7__3095_
timestamp 1701859473
transform 1 0 10270 0 1 5470
box -12 -8 32 272
use FILL  FILL_7__3096_
timestamp 1701859473
transform 1 0 9010 0 1 6510
box -12 -8 32 272
use FILL  FILL_7__3097_
timestamp 1701859473
transform -1 0 8790 0 1 6510
box -12 -8 32 272
use FILL  FILL_7__3098_
timestamp 1701859473
transform -1 0 10490 0 1 8070
box -12 -8 32 272
use FILL  FILL_7__3099_
timestamp 1701859473
transform -1 0 11250 0 -1 8070
box -12 -8 32 272
use FILL  FILL_7__3100_
timestamp 1701859473
transform 1 0 10250 0 1 8070
box -12 -8 32 272
use FILL  FILL_7__3102_
timestamp 1701859473
transform 1 0 8470 0 -1 8070
box -12 -8 32 272
use FILL  FILL_7__3103_
timestamp 1701859473
transform -1 0 8450 0 1 7550
box -12 -8 32 272
use FILL  FILL_7__3104_
timestamp 1701859473
transform -1 0 11250 0 1 6510
box -12 -8 32 272
use FILL  FILL_7__3105_
timestamp 1701859473
transform -1 0 11050 0 -1 4950
box -12 -8 32 272
use FILL  FILL_7__3106_
timestamp 1701859473
transform 1 0 9470 0 -1 8590
box -12 -8 32 272
use FILL  FILL_7__3107_
timestamp 1701859473
transform -1 0 9710 0 -1 8590
box -12 -8 32 272
use FILL  FILL_7__3109_
timestamp 1701859473
transform -1 0 9850 0 1 5470
box -12 -8 32 272
use FILL  FILL_7__3110_
timestamp 1701859473
transform 1 0 8490 0 -1 6510
box -12 -8 32 272
use FILL  FILL_7__3111_
timestamp 1701859473
transform -1 0 8270 0 -1 6510
box -12 -8 32 272
use FILL  FILL_7__3112_
timestamp 1701859473
transform 1 0 610 0 -1 2870
box -12 -8 32 272
use FILL  FILL_7__3113_
timestamp 1701859473
transform 1 0 150 0 -1 2870
box -12 -8 32 272
use FILL  FILL_7__3114_
timestamp 1701859473
transform -1 0 410 0 -1 2870
box -12 -8 32 272
use FILL  FILL_7__3115_
timestamp 1701859473
transform -1 0 1290 0 1 2350
box -12 -8 32 272
use FILL  FILL_7__3117_
timestamp 1701859473
transform 1 0 2130 0 -1 1310
box -12 -8 32 272
use FILL  FILL_7__3118_
timestamp 1701859473
transform -1 0 1510 0 -1 2350
box -12 -8 32 272
use FILL  FILL_7__3119_
timestamp 1701859473
transform -1 0 1270 0 -1 2350
box -12 -8 32 272
use FILL  FILL_7__3120_
timestamp 1701859473
transform -1 0 570 0 1 2350
box -12 -8 32 272
use FILL  FILL_7__3121_
timestamp 1701859473
transform 1 0 350 0 1 2870
box -12 -8 32 272
use FILL  FILL_7__3122_
timestamp 1701859473
transform 1 0 2610 0 -1 3390
box -12 -8 32 272
use FILL  FILL_7__3124_
timestamp 1701859473
transform -1 0 410 0 1 3390
box -12 -8 32 272
use FILL  FILL_7__3125_
timestamp 1701859473
transform -1 0 830 0 -1 2350
box -12 -8 32 272
use FILL  FILL_7__3126_
timestamp 1701859473
transform -1 0 1530 0 1 2350
box -12 -8 32 272
use FILL  FILL_7__3127_
timestamp 1701859473
transform -1 0 1050 0 1 2350
box -12 -8 32 272
use FILL  FILL_7__3128_
timestamp 1701859473
transform -1 0 1990 0 1 2350
box -12 -8 32 272
use FILL  FILL_7__3129_
timestamp 1701859473
transform -1 0 1750 0 -1 2350
box -12 -8 32 272
use FILL  FILL_7__3131_
timestamp 1701859473
transform -1 0 810 0 1 2350
box -12 -8 32 272
use FILL  FILL_7__3132_
timestamp 1701859473
transform 1 0 570 0 1 2870
box -12 -8 32 272
use FILL  FILL_7__3133_
timestamp 1701859473
transform 1 0 630 0 -1 3910
box -12 -8 32 272
use FILL  FILL_7__3134_
timestamp 1701859473
transform -1 0 1310 0 1 3390
box -12 -8 32 272
use FILL  FILL_7__3135_
timestamp 1701859473
transform 1 0 1070 0 1 3390
box -12 -8 32 272
use FILL  FILL_7__3136_
timestamp 1701859473
transform -1 0 650 0 -1 3390
box -12 -8 32 272
use FILL  FILL_7__3137_
timestamp 1701859473
transform 1 0 370 0 -1 3390
box -12 -8 32 272
use FILL  FILL_7__3139_
timestamp 1701859473
transform -1 0 1970 0 -1 3390
box -12 -8 32 272
use FILL  FILL_7__3140_
timestamp 1701859473
transform -1 0 390 0 1 3910
box -12 -8 32 272
use FILL  FILL_7__3141_
timestamp 1701859473
transform 1 0 830 0 1 4430
box -12 -8 32 272
use FILL  FILL_7__3142_
timestamp 1701859473
transform 1 0 1070 0 1 4430
box -12 -8 32 272
use FILL  FILL_7__3143_
timestamp 1701859473
transform 1 0 1090 0 -1 4430
box -12 -8 32 272
use FILL  FILL_7__3144_
timestamp 1701859473
transform -1 0 1330 0 -1 4430
box -12 -8 32 272
use FILL  FILL_7__3146_
timestamp 1701859473
transform -1 0 830 0 1 3910
box -12 -8 32 272
use FILL  FILL_7__3147_
timestamp 1701859473
transform 1 0 610 0 -1 4430
box -12 -8 32 272
use FILL  FILL_7__3148_
timestamp 1701859473
transform -1 0 870 0 -1 4430
box -12 -8 32 272
use FILL  FILL_7__3149_
timestamp 1701859473
transform -1 0 170 0 -1 3910
box -12 -8 32 272
use FILL  FILL_7__3150_
timestamp 1701859473
transform -1 0 1030 0 1 3910
box -12 -8 32 272
use FILL  FILL_7__3151_
timestamp 1701859473
transform 1 0 150 0 1 3910
box -12 -8 32 272
use FILL  FILL_7__3153_
timestamp 1701859473
transform -1 0 390 0 -1 4430
box -12 -8 32 272
use FILL  FILL_7__3154_
timestamp 1701859473
transform -1 0 890 0 -1 3390
box -12 -8 32 272
use FILL  FILL_7__3155_
timestamp 1701859473
transform -1 0 170 0 1 2870
box -12 -8 32 272
use FILL  FILL_7__3156_
timestamp 1701859473
transform 1 0 150 0 -1 3390
box -12 -8 32 272
use FILL  FILL_7__3157_
timestamp 1701859473
transform -1 0 170 0 1 3390
box -12 -8 32 272
use FILL  FILL_7__3158_
timestamp 1701859473
transform 1 0 150 0 1 4430
box -12 -8 32 272
use FILL  FILL_7__3160_
timestamp 1701859473
transform -1 0 610 0 1 4430
box -12 -8 32 272
use FILL  FILL_7__3161_
timestamp 1701859473
transform 1 0 4250 0 -1 7030
box -12 -8 32 272
use FILL  FILL_7__3162_
timestamp 1701859473
transform -1 0 4490 0 -1 7030
box -12 -8 32 272
use FILL  FILL_7__3163_
timestamp 1701859473
transform 1 0 4710 0 -1 7030
box -12 -8 32 272
use FILL  FILL_7__3164_
timestamp 1701859473
transform 1 0 4950 0 1 7030
box -12 -8 32 272
use FILL  FILL_7__3165_
timestamp 1701859473
transform 1 0 4210 0 1 7550
box -12 -8 32 272
use FILL  FILL_7__3166_
timestamp 1701859473
transform -1 0 4450 0 1 7550
box -12 -8 32 272
use FILL  FILL_7__3168_
timestamp 1701859473
transform 1 0 5130 0 -1 10150
box -12 -8 32 272
use FILL  FILL_7__3169_
timestamp 1701859473
transform -1 0 3770 0 -1 10670
box -12 -8 32 272
use FILL  FILL_7__3170_
timestamp 1701859473
transform -1 0 3990 0 -1 10670
box -12 -8 32 272
use FILL  FILL_7__3171_
timestamp 1701859473
transform 1 0 4410 0 -1 10670
box -12 -8 32 272
use FILL  FILL_7__3172_
timestamp 1701859473
transform -1 0 4650 0 -1 10670
box -12 -8 32 272
use FILL  FILL_7__3173_
timestamp 1701859473
transform 1 0 4250 0 1 10150
box -12 -8 32 272
use FILL  FILL_7__3175_
timestamp 1701859473
transform 1 0 5590 0 1 10150
box -12 -8 32 272
use FILL  FILL_7__3176_
timestamp 1701859473
transform 1 0 5350 0 1 10150
box -12 -8 32 272
use FILL  FILL_7__3177_
timestamp 1701859473
transform -1 0 1830 0 -1 5990
box -12 -8 32 272
use FILL  FILL_7__3178_
timestamp 1701859473
transform 1 0 2270 0 -1 5990
box -12 -8 32 272
use FILL  FILL_7__3179_
timestamp 1701859473
transform -1 0 1550 0 1 6510
box -12 -8 32 272
use FILL  FILL_7__3180_
timestamp 1701859473
transform -1 0 1770 0 1 6510
box -12 -8 32 272
use FILL  FILL_7__3182_
timestamp 1701859473
transform -1 0 1030 0 -1 6510
box -12 -8 32 272
use FILL  FILL_7__3183_
timestamp 1701859473
transform 1 0 390 0 1 8070
box -12 -8 32 272
use FILL  FILL_7__3184_
timestamp 1701859473
transform -1 0 630 0 1 8070
box -12 -8 32 272
use FILL  FILL_7__3185_
timestamp 1701859473
transform -1 0 170 0 -1 8590
box -12 -8 32 272
use FILL  FILL_7__3186_
timestamp 1701859473
transform -1 0 170 0 1 8070
box -12 -8 32 272
use FILL  FILL_7__3187_
timestamp 1701859473
transform 1 0 790 0 -1 9110
box -12 -8 32 272
use FILL  FILL_7__3188_
timestamp 1701859473
transform 1 0 1010 0 -1 9110
box -12 -8 32 272
use FILL  FILL_7__3190_
timestamp 1701859473
transform 1 0 2430 0 1 9110
box -12 -8 32 272
use FILL  FILL_7__3191_
timestamp 1701859473
transform 1 0 1490 0 -1 9110
box -12 -8 32 272
use FILL  FILL_7__3192_
timestamp 1701859473
transform -1 0 1730 0 -1 9110
box -12 -8 32 272
use FILL  FILL_7__3324_
timestamp 1701859473
transform 1 0 5670 0 1 8070
box -12 -8 32 272
use FILL  FILL_7__3325_
timestamp 1701859473
transform -1 0 6390 0 1 8070
box -12 -8 32 272
use FILL  FILL_7__3326_
timestamp 1701859473
transform -1 0 6290 0 -1 8070
box -12 -8 32 272
use FILL  FILL_7__3328_
timestamp 1701859473
transform -1 0 6150 0 1 8070
box -12 -8 32 272
use FILL  FILL_7__3329_
timestamp 1701859473
transform 1 0 5910 0 1 8070
box -12 -8 32 272
use FILL  FILL_7__3330_
timestamp 1701859473
transform -1 0 7090 0 1 8590
box -12 -8 32 272
use FILL  FILL_7__3331_
timestamp 1701859473
transform 1 0 7370 0 -1 8590
box -12 -8 32 272
use FILL  FILL_7__3332_
timestamp 1701859473
transform 1 0 7090 0 -1 8590
box -12 -8 32 272
use FILL  FILL_7__3333_
timestamp 1701859473
transform 1 0 10290 0 1 8590
box -12 -8 32 272
use FILL  FILL_7__3335_
timestamp 1701859473
transform 1 0 7950 0 -1 10150
box -12 -8 32 272
use FILL  FILL_7__3336_
timestamp 1701859473
transform -1 0 6790 0 1 9630
box -12 -8 32 272
use FILL  FILL_7__3337_
timestamp 1701859473
transform -1 0 6310 0 1 9630
box -12 -8 32 272
use FILL  FILL_7__3338_
timestamp 1701859473
transform 1 0 7270 0 -1 10150
box -12 -8 32 272
use FILL  FILL_7__3339_
timestamp 1701859473
transform -1 0 8150 0 1 10150
box -12 -8 32 272
use FILL  FILL_7__3340_
timestamp 1701859473
transform 1 0 7910 0 1 10150
box -12 -8 32 272
use FILL  FILL_7__3342_
timestamp 1701859473
transform 1 0 6890 0 -1 11190
box -12 -8 32 272
use FILL  FILL_7__3343_
timestamp 1701859473
transform -1 0 7490 0 -1 10150
box -12 -8 32 272
use FILL  FILL_7__3344_
timestamp 1701859473
transform 1 0 7710 0 -1 10150
box -12 -8 32 272
use FILL  FILL_7__3345_
timestamp 1701859473
transform -1 0 9090 0 1 9630
box -12 -8 32 272
use FILL  FILL_7__3346_
timestamp 1701859473
transform 1 0 8610 0 1 10150
box -12 -8 32 272
use FILL  FILL_7__3347_
timestamp 1701859473
transform -1 0 8390 0 1 10150
box -12 -8 32 272
use FILL  FILL_7__3348_
timestamp 1701859473
transform 1 0 9210 0 -1 10670
box -12 -8 32 272
use FILL  FILL_7__3350_
timestamp 1701859473
transform 1 0 7650 0 -1 8590
box -12 -8 32 272
use FILL  FILL_7__3351_
timestamp 1701859473
transform -1 0 7830 0 1 8590
box -12 -8 32 272
use FILL  FILL_7__3352_
timestamp 1701859473
transform -1 0 8290 0 -1 9110
box -12 -8 32 272
use FILL  FILL_7__3353_
timestamp 1701859473
transform 1 0 8170 0 -1 10150
box -12 -8 32 272
use FILL  FILL_7__3354_
timestamp 1701859473
transform 1 0 7850 0 -1 10670
box -12 -8 32 272
use FILL  FILL_7__3355_
timestamp 1701859473
transform -1 0 7630 0 -1 10670
box -12 -8 32 272
use FILL  FILL_7__3357_
timestamp 1701859473
transform 1 0 7230 0 1 10670
box -12 -8 32 272
use FILL  FILL_7__3358_
timestamp 1701859473
transform 1 0 7490 0 1 10670
box -12 -8 32 272
use FILL  FILL_7__3359_
timestamp 1701859473
transform 1 0 7730 0 1 10670
box -12 -8 32 272
use FILL  FILL_7__3360_
timestamp 1701859473
transform -1 0 7990 0 1 10670
box -12 -8 32 272
use FILL  FILL_7__3361_
timestamp 1701859473
transform 1 0 9010 0 -1 10670
box -12 -8 32 272
use FILL  FILL_7__3362_
timestamp 1701859473
transform 1 0 8070 0 -1 10670
box -12 -8 32 272
use FILL  FILL_7__3364_
timestamp 1701859473
transform 1 0 8030 0 -1 11190
box -12 -8 32 272
use FILL  FILL_7__3365_
timestamp 1701859473
transform -1 0 7570 0 -1 11190
box -12 -8 32 272
use FILL  FILL_7__3366_
timestamp 1701859473
transform 1 0 7090 0 -1 11190
box -12 -8 32 272
use FILL  FILL_7__3367_
timestamp 1701859473
transform 1 0 6970 0 1 10670
box -12 -8 32 272
use FILL  FILL_7__3368_
timestamp 1701859473
transform 1 0 7310 0 -1 11190
box -12 -8 32 272
use FILL  FILL_7__3369_
timestamp 1701859473
transform 1 0 7790 0 -1 11190
box -12 -8 32 272
use FILL  FILL_7__3371_
timestamp 1701859473
transform 1 0 8410 0 1 10670
box -12 -8 32 272
use FILL  FILL_7__3372_
timestamp 1701859473
transform 1 0 9590 0 1 10670
box -12 -8 32 272
use FILL  FILL_7__3373_
timestamp 1701859473
transform -1 0 6690 0 -1 11190
box -12 -8 32 272
use FILL  FILL_7__3374_
timestamp 1701859473
transform 1 0 5790 0 1 10670
box -12 -8 32 272
use FILL  FILL_7__3375_
timestamp 1701859473
transform -1 0 6050 0 1 10670
box -12 -8 32 272
use FILL  FILL_7__3376_
timestamp 1701859473
transform -1 0 6270 0 1 10670
box -12 -8 32 272
use FILL  FILL_7__3377_
timestamp 1701859473
transform 1 0 6510 0 1 10670
box -12 -8 32 272
use FILL  FILL_7__3379_
timestamp 1701859473
transform 1 0 8770 0 -1 10670
box -12 -8 32 272
use FILL  FILL_7__3380_
timestamp 1701859473
transform 1 0 8890 0 1 10670
box -12 -8 32 272
use FILL  FILL_7__3381_
timestamp 1701859473
transform -1 0 6770 0 1 10670
box -12 -8 32 272
use FILL  FILL_7__3382_
timestamp 1701859473
transform 1 0 6230 0 -1 10670
box -12 -8 32 272
use FILL  FILL_7__3383_
timestamp 1701859473
transform -1 0 6490 0 -1 10670
box -12 -8 32 272
use FILL  FILL_7__3384_
timestamp 1701859473
transform -1 0 6930 0 -1 10670
box -12 -8 32 272
use FILL  FILL_7__3386_
timestamp 1701859473
transform 1 0 7170 0 -1 10670
box -12 -8 32 272
use FILL  FILL_7__3387_
timestamp 1701859473
transform 1 0 8530 0 -1 10670
box -12 -8 32 272
use FILL  FILL_7__3388_
timestamp 1701859473
transform 1 0 8650 0 1 10670
box -12 -8 32 272
use FILL  FILL_7__3389_
timestamp 1701859473
transform 1 0 10310 0 -1 10670
box -12 -8 32 272
use FILL  FILL_7__3390_
timestamp 1701859473
transform 1 0 9870 0 -1 10670
box -12 -8 32 272
use FILL  FILL_7__3391_
timestamp 1701859473
transform 1 0 10070 0 -1 10670
box -12 -8 32 272
use FILL  FILL_7__3393_
timestamp 1701859473
transform -1 0 11270 0 -1 10150
box -12 -8 32 272
use FILL  FILL_7__3394_
timestamp 1701859473
transform 1 0 7450 0 1 10150
box -12 -8 32 272
use FILL  FILL_7__3395_
timestamp 1701859473
transform 1 0 6510 0 1 10150
box -12 -8 32 272
use FILL  FILL_7__3396_
timestamp 1701859473
transform -1 0 6770 0 1 10150
box -12 -8 32 272
use FILL  FILL_7__3397_
timestamp 1701859473
transform -1 0 7090 0 -1 10150
box -12 -8 32 272
use FILL  FILL_7__3398_
timestamp 1701859473
transform 1 0 6370 0 -1 10150
box -12 -8 32 272
use FILL  FILL_7__3399_
timestamp 1701859473
transform -1 0 6850 0 -1 10150
box -12 -8 32 272
use FILL  FILL_7__3401_
timestamp 1701859473
transform 1 0 7210 0 1 10150
box -12 -8 32 272
use FILL  FILL_7__3402_
timestamp 1701859473
transform -1 0 9150 0 1 10150
box -12 -8 32 272
use FILL  FILL_7__3403_
timestamp 1701859473
transform 1 0 9590 0 1 10150
box -12 -8 32 272
use FILL  FILL_7__3404_
timestamp 1701859473
transform -1 0 5850 0 1 9630
box -12 -8 32 272
use FILL  FILL_7__3405_
timestamp 1701859473
transform -1 0 6130 0 -1 10150
box -12 -8 32 272
use FILL  FILL_7__3406_
timestamp 1701859473
transform 1 0 6490 0 -1 9630
box -12 -8 32 272
use FILL  FILL_7__3408_
timestamp 1701859473
transform 1 0 6970 0 1 9630
box -12 -8 32 272
use FILL  FILL_7__3409_
timestamp 1701859473
transform -1 0 6590 0 -1 10150
box -12 -8 32 272
use FILL  FILL_7__3410_
timestamp 1701859473
transform 1 0 9330 0 -1 10150
box -12 -8 32 272
use FILL  FILL_7__3411_
timestamp 1701859473
transform 1 0 9350 0 1 10150
box -12 -8 32 272
use FILL  FILL_7__3412_
timestamp 1701859473
transform 1 0 10070 0 1 10150
box -12 -8 32 272
use FILL  FILL_7__3413_
timestamp 1701859473
transform -1 0 6090 0 1 9630
box -12 -8 32 272
use FILL  FILL_7__3415_
timestamp 1701859473
transform 1 0 6510 0 1 9630
box -12 -8 32 272
use FILL  FILL_7__3416_
timestamp 1701859473
transform 1 0 7350 0 1 8590
box -12 -8 32 272
use FILL  FILL_7__3417_
timestamp 1701859473
transform 1 0 7430 0 -1 9110
box -12 -8 32 272
use FILL  FILL_7__3418_
timestamp 1701859473
transform -1 0 7570 0 -1 9630
box -12 -8 32 272
use FILL  FILL_7__3419_
timestamp 1701859473
transform 1 0 7330 0 -1 9630
box -12 -8 32 272
use FILL  FILL_7__3420_
timestamp 1701859473
transform -1 0 6910 0 -1 9630
box -12 -8 32 272
use FILL  FILL_7__3422_
timestamp 1701859473
transform -1 0 7230 0 1 9630
box -12 -8 32 272
use FILL  FILL_7__3423_
timestamp 1701859473
transform -1 0 8290 0 -1 9630
box -12 -8 32 272
use FILL  FILL_7__3424_
timestamp 1701859473
transform -1 0 7810 0 -1 9630
box -12 -8 32 272
use FILL  FILL_7__3425_
timestamp 1701859473
transform -1 0 7470 0 1 9630
box -12 -8 32 272
use FILL  FILL_7__3426_
timestamp 1701859473
transform -1 0 9110 0 -1 10150
box -12 -8 32 272
use FILL  FILL_7__3427_
timestamp 1701859473
transform 1 0 8870 0 -1 10150
box -12 -8 32 272
use FILL  FILL_7__3428_
timestamp 1701859473
transform 1 0 7550 0 1 8590
box -12 -8 32 272
use FILL  FILL_7__3430_
timestamp 1701859473
transform -1 0 7850 0 -1 9110
box -12 -8 32 272
use FILL  FILL_7__3431_
timestamp 1701859473
transform 1 0 7770 0 1 9110
box -12 -8 32 272
use FILL  FILL_7__3432_
timestamp 1701859473
transform 1 0 8010 0 1 9110
box -12 -8 32 272
use FILL  FILL_7__3433_
timestamp 1701859473
transform -1 0 8050 0 -1 9630
box -12 -8 32 272
use FILL  FILL_7__3434_
timestamp 1701859473
transform 1 0 7690 0 1 9630
box -12 -8 32 272
use FILL  FILL_7__3435_
timestamp 1701859473
transform 1 0 10310 0 1 10150
box -12 -8 32 272
use FILL  FILL_7__3437_
timestamp 1701859473
transform 1 0 10750 0 1 10150
box -12 -8 32 272
use FILL  FILL_7__3438_
timestamp 1701859473
transform 1 0 10530 0 1 10150
box -12 -8 32 272
use FILL  FILL_7__3439_
timestamp 1701859473
transform 1 0 10970 0 1 10150
box -12 -8 32 272
use FILL  FILL_7__3440_
timestamp 1701859473
transform -1 0 10790 0 -1 10150
box -12 -8 32 272
use FILL  FILL_7__3441_
timestamp 1701859473
transform -1 0 10650 0 1 9630
box -12 -8 32 272
use FILL  FILL_7__3442_
timestamp 1701859473
transform -1 0 10530 0 -1 10150
box -12 -8 32 272
use FILL  FILL_7__3444_
timestamp 1701859473
transform -1 0 8490 0 -1 9630
box -12 -8 32 272
use FILL  FILL_7__3445_
timestamp 1701859473
transform -1 0 8190 0 1 9630
box -12 -8 32 272
use FILL  FILL_7__3446_
timestamp 1701859473
transform 1 0 8630 0 1 9630
box -12 -8 32 272
use FILL  FILL_7__3447_
timestamp 1701859473
transform 1 0 8410 0 1 9630
box -12 -8 32 272
use FILL  FILL_7__3448_
timestamp 1701859473
transform -1 0 8850 0 1 9630
box -12 -8 32 272
use FILL  FILL_7__3449_
timestamp 1701859473
transform -1 0 9890 0 1 10150
box -12 -8 32 272
use FILL  FILL_7__3451_
timestamp 1701859473
transform 1 0 9570 0 -1 10150
box -12 -8 32 272
use FILL  FILL_7__3452_
timestamp 1701859473
transform -1 0 9310 0 1 9630
box -12 -8 32 272
use FILL  FILL_7__3453_
timestamp 1701859473
transform -1 0 10070 0 -1 10150
box -12 -8 32 272
use FILL  FILL_7__3454_
timestamp 1701859473
transform 1 0 9510 0 1 9630
box -12 -8 32 272
use FILL  FILL_7__3455_
timestamp 1701859473
transform 1 0 9730 0 1 9630
box -12 -8 32 272
use FILL  FILL_7__3456_
timestamp 1701859473
transform -1 0 10430 0 1 9630
box -12 -8 32 272
use FILL  FILL_7__3457_
timestamp 1701859473
transform -1 0 9970 0 1 9630
box -12 -8 32 272
use FILL  FILL_7__3459_
timestamp 1701859473
transform -1 0 10350 0 -1 9630
box -12 -8 32 272
use FILL  FILL_7__3460_
timestamp 1701859473
transform 1 0 11010 0 -1 10150
box -12 -8 32 272
use FILL  FILL_7__3461_
timestamp 1701859473
transform -1 0 11250 0 -1 9630
box -12 -8 32 272
use FILL  FILL_7__3462_
timestamp 1701859473
transform -1 0 10790 0 -1 9630
box -12 -8 32 272
use FILL  FILL_7__3463_
timestamp 1701859473
transform 1 0 10470 0 -1 11190
box -12 -8 32 272
use FILL  FILL_7__3464_
timestamp 1701859473
transform 1 0 9810 0 -1 11190
box -12 -8 32 272
use FILL  FILL_7__3466_
timestamp 1701859473
transform 1 0 10230 0 -1 11190
box -12 -8 32 272
use FILL  FILL_7__3467_
timestamp 1701859473
transform -1 0 11210 0 1 10670
box -12 -8 32 272
use FILL  FILL_7__3468_
timestamp 1701859473
transform 1 0 10710 0 1 10670
box -12 -8 32 272
use FILL  FILL_7__3469_
timestamp 1701859473
transform 1 0 9430 0 -1 10670
box -12 -8 32 272
use FILL  FILL_7__3470_
timestamp 1701859473
transform 1 0 9670 0 -1 10670
box -12 -8 32 272
use FILL  FILL_7__3471_
timestamp 1701859473
transform 1 0 9810 0 1 10670
box -12 -8 32 272
use FILL  FILL_7__3473_
timestamp 1701859473
transform 1 0 8690 0 -1 11190
box -12 -8 32 272
use FILL  FILL_7__3474_
timestamp 1701859473
transform 1 0 8250 0 -1 11190
box -12 -8 32 272
use FILL  FILL_7__3475_
timestamp 1701859473
transform 1 0 8490 0 -1 11190
box -12 -8 32 272
use FILL  FILL_7__3476_
timestamp 1701859473
transform -1 0 8930 0 -1 11190
box -12 -8 32 272
use FILL  FILL_7__3477_
timestamp 1701859473
transform 1 0 9150 0 -1 11190
box -12 -8 32 272
use FILL  FILL_7__3478_
timestamp 1701859473
transform 1 0 9130 0 1 10670
box -12 -8 32 272
use FILL  FILL_7__3479_
timestamp 1701859473
transform 1 0 8410 0 -1 10150
box -12 -8 32 272
use FILL  FILL_7__3481_
timestamp 1701859473
transform -1 0 8450 0 1 9110
box -12 -8 32 272
use FILL  FILL_7__3482_
timestamp 1701859473
transform -1 0 8670 0 1 9110
box -12 -8 32 272
use FILL  FILL_7__3483_
timestamp 1701859473
transform 1 0 8850 0 1 10150
box -12 -8 32 272
use FILL  FILL_7__3484_
timestamp 1701859473
transform -1 0 10150 0 -1 9630
box -12 -8 32 272
use FILL  FILL_7__3485_
timestamp 1701859473
transform 1 0 11170 0 1 10150
box -12 -8 32 272
use FILL  FILL_7__3486_
timestamp 1701859473
transform 1 0 10510 0 1 9110
box -12 -8 32 272
use FILL  FILL_7__3488_
timestamp 1701859473
transform -1 0 10850 0 1 9630
box -12 -8 32 272
use FILL  FILL_7__3489_
timestamp 1701859473
transform 1 0 10690 0 -1 11190
box -12 -8 32 272
use FILL  FILL_7__3490_
timestamp 1701859473
transform 1 0 11150 0 -1 11190
box -12 -8 32 272
use FILL  FILL_7__3491_
timestamp 1701859473
transform -1 0 10950 0 -1 11190
box -12 -8 32 272
use FILL  FILL_7__3492_
timestamp 1701859473
transform -1 0 10510 0 1 10670
box -12 -8 32 272
use FILL  FILL_7__3493_
timestamp 1701859473
transform -1 0 10290 0 1 10670
box -12 -8 32 272
use FILL  FILL_7__3495_
timestamp 1701859473
transform -1 0 9590 0 -1 11190
box -12 -8 32 272
use FILL  FILL_7__3496_
timestamp 1701859473
transform 1 0 9350 0 -1 11190
box -12 -8 32 272
use FILL  FILL_7__3497_
timestamp 1701859473
transform -1 0 9450 0 -1 9630
box -12 -8 32 272
use FILL  FILL_7__3498_
timestamp 1701859473
transform -1 0 8950 0 1 9110
box -12 -8 32 272
use FILL  FILL_7__3499_
timestamp 1701859473
transform 1 0 8470 0 -1 9110
box -12 -8 32 272
use FILL  FILL_7__3500_
timestamp 1701859473
transform 1 0 9850 0 1 9110
box -12 -8 32 272
use FILL  FILL_7__3502_
timestamp 1701859473
transform -1 0 8350 0 -1 8590
box -12 -8 32 272
use FILL  FILL_7__3503_
timestamp 1701859473
transform -1 0 8730 0 -1 9630
box -12 -8 32 272
use FILL  FILL_7__3504_
timestamp 1701859473
transform 1 0 8950 0 -1 9630
box -12 -8 32 272
use FILL  FILL_7__3505_
timestamp 1701859473
transform -1 0 9210 0 -1 9630
box -12 -8 32 272
use FILL  FILL_7__3506_
timestamp 1701859473
transform -1 0 8730 0 1 8590
box -12 -8 32 272
use FILL  FILL_7__3507_
timestamp 1701859473
transform 1 0 10810 0 -1 9110
box -12 -8 32 272
use FILL  FILL_7__3508_
timestamp 1701859473
transform 1 0 10570 0 -1 9110
box -12 -8 32 272
use FILL  FILL_7__3510_
timestamp 1701859473
transform -1 0 8970 0 1 8590
box -12 -8 32 272
use FILL  FILL_7__3511_
timestamp 1701859473
transform 1 0 10030 0 -1 270
box -12 -8 32 272
use FILL  FILL_7__3512_
timestamp 1701859473
transform 1 0 11030 0 -1 9110
box -12 -8 32 272
use FILL  FILL_7__3513_
timestamp 1701859473
transform 1 0 11010 0 -1 9630
box -12 -8 32 272
use FILL  FILL_7__3514_
timestamp 1701859473
transform 1 0 10970 0 1 10670
box -12 -8 32 272
use FILL  FILL_7__3515_
timestamp 1701859473
transform -1 0 10770 0 -1 10670
box -12 -8 32 272
use FILL  FILL_7__3517_
timestamp 1701859473
transform 1 0 9670 0 -1 9630
box -12 -8 32 272
use FILL  FILL_7__3518_
timestamp 1701859473
transform 1 0 9890 0 -1 9630
box -12 -8 32 272
use FILL  FILL_7__3519_
timestamp 1701859473
transform 1 0 9170 0 1 9110
box -12 -8 32 272
use FILL  FILL_7__3520_
timestamp 1701859473
transform -1 0 9410 0 1 9110
box -12 -8 32 272
use FILL  FILL_7__3521_
timestamp 1701859473
transform 1 0 6650 0 1 8590
box -12 -8 32 272
use FILL  FILL_7__3522_
timestamp 1701859473
transform 1 0 8050 0 -1 9110
box -12 -8 32 272
use FILL  FILL_7__3524_
timestamp 1701859473
transform 1 0 7570 0 1 9110
box -12 -8 32 272
use FILL  FILL_7__3525_
timestamp 1701859473
transform 1 0 7110 0 1 9110
box -12 -8 32 272
use FILL  FILL_7__3526_
timestamp 1701859473
transform -1 0 7350 0 1 9110
box -12 -8 32 272
use FILL  FILL_7__3539_
timestamp 1701859473
transform 1 0 11210 0 -1 7030
box -12 -8 32 272
use FILL  FILL_7__3540_
timestamp 1701859473
transform 1 0 4710 0 1 10670
box -12 -8 32 272
use FILL  FILL_7__3541_
timestamp 1701859473
transform -1 0 170 0 1 5990
box -12 -8 32 272
use FILL  FILL_7__3542_
timestamp 1701859473
transform -1 0 170 0 -1 8070
box -12 -8 32 272
use FILL  FILL_7__3544_
timestamp 1701859473
transform -1 0 170 0 1 9110
box -12 -8 32 272
use FILL  FILL_7__3545_
timestamp 1701859473
transform -1 0 2010 0 -1 11190
box -12 -8 32 272
use FILL  FILL_7__3546_
timestamp 1701859473
transform -1 0 630 0 1 9110
box -12 -8 32 272
use FILL  FILL_7__3547_
timestamp 1701859473
transform 1 0 4750 0 -1 11190
box -12 -8 32 272
use FILL  FILL_7__3548_
timestamp 1701859473
transform 1 0 5350 0 1 10670
box -12 -8 32 272
use FILL  FILL_7__3549_
timestamp 1701859473
transform -1 0 4350 0 -1 11190
box -12 -8 32 272
use FILL  FILL_7__3551_
timestamp 1701859473
transform 1 0 5590 0 -1 11190
box -12 -8 32 272
use FILL  FILL_7__3552_
timestamp 1701859473
transform 1 0 5370 0 -1 11190
box -12 -8 32 272
use FILL  FILL_7__3553_
timestamp 1701859473
transform -1 0 170 0 -1 5990
box -12 -8 32 272
use FILL  FILL_7__3554_
timestamp 1701859473
transform -1 0 370 0 1 7030
box -12 -8 32 272
use FILL  FILL_7__3555_
timestamp 1701859473
transform -1 0 5150 0 1 10670
box -12 -8 32 272
use FILL  FILL_7__3556_
timestamp 1701859473
transform 1 0 6290 0 1 10150
box -12 -8 32 272
use FILL  FILL_7__3558_
timestamp 1701859473
transform 1 0 6230 0 -1 11190
box -12 -8 32 272
use FILL  FILL_7__3559_
timestamp 1701859473
transform -1 0 4890 0 -1 10670
box -12 -8 32 272
use FILL  FILL_7__3560_
timestamp 1701859473
transform 1 0 5570 0 1 10670
box -12 -8 32 272
use FILL  FILL_7__3561_
timestamp 1701859473
transform 1 0 6010 0 -1 11190
box -12 -8 32 272
use FILL  FILL_7__3562_
timestamp 1701859473
transform 1 0 5810 0 1 10150
box -12 -8 32 272
use FILL  FILL_7__3563_
timestamp 1701859473
transform 1 0 5270 0 1 3390
box -12 -8 32 272
use FILL  FILL_7_BUFX2_insert0
timestamp 1701859473
transform 1 0 5890 0 -1 10150
box -12 -8 32 272
use FILL  FILL_7_BUFX2_insert1
timestamp 1701859473
transform 1 0 6650 0 1 2350
box -12 -8 32 272
use FILL  FILL_7_BUFX2_insert2
timestamp 1701859473
transform 1 0 5490 0 -1 1830
box -12 -8 32 272
use FILL  FILL_7_BUFX2_insert3
timestamp 1701859473
transform -1 0 630 0 -1 5470
box -12 -8 32 272
use FILL  FILL_7_BUFX2_insert4
timestamp 1701859473
transform 1 0 3370 0 1 4950
box -12 -8 32 272
use FILL  FILL_7_BUFX2_insert5
timestamp 1701859473
transform 1 0 1430 0 -1 1830
box -12 -8 32 272
use FILL  FILL_7_BUFX2_insert7
timestamp 1701859473
transform 1 0 1730 0 1 10670
box -12 -8 32 272
use FILL  FILL_7_BUFX2_insert8
timestamp 1701859473
transform 1 0 1690 0 1 1830
box -12 -8 32 272
use FILL  FILL_7_BUFX2_insert9
timestamp 1701859473
transform 1 0 1990 0 -1 3910
box -12 -8 32 272
use FILL  FILL_7_BUFX2_insert10
timestamp 1701859473
transform 1 0 1810 0 -1 4430
box -12 -8 32 272
use FILL  FILL_7_BUFX2_insert11
timestamp 1701859473
transform -1 0 1790 0 -1 3910
box -12 -8 32 272
use FILL  FILL_7_BUFX2_insert12
timestamp 1701859473
transform -1 0 1570 0 -1 3910
box -12 -8 32 272
use FILL  FILL_7_BUFX2_insert13
timestamp 1701859473
transform -1 0 1470 0 -1 1310
box -12 -8 32 272
use FILL  FILL_7_BUFX2_insert15
timestamp 1701859473
transform 1 0 4590 0 -1 5470
box -12 -8 32 272
use FILL  FILL_7_BUFX2_insert16
timestamp 1701859473
transform 1 0 1390 0 -1 4950
box -12 -8 32 272
use FILL  FILL_7_BUFX2_insert17
timestamp 1701859473
transform 1 0 3670 0 1 1310
box -12 -8 32 272
use FILL  FILL_7_BUFX2_insert18
timestamp 1701859473
transform -1 0 9810 0 1 2350
box -12 -8 32 272
use FILL  FILL_7_BUFX2_insert19
timestamp 1701859473
transform -1 0 8550 0 -1 790
box -12 -8 32 272
use FILL  FILL_7_BUFX2_insert20
timestamp 1701859473
transform 1 0 10010 0 1 2350
box -12 -8 32 272
use FILL  FILL_7_BUFX2_insert22
timestamp 1701859473
transform -1 0 3250 0 -1 2870
box -12 -8 32 272
use FILL  FILL_7_BUFX2_insert23
timestamp 1701859473
transform -1 0 2790 0 -1 4950
box -12 -8 32 272
use FILL  FILL_7_BUFX2_insert24
timestamp 1701859473
transform -1 0 3690 0 -1 4430
box -12 -8 32 272
use FILL  FILL_7_BUFX2_insert25
timestamp 1701859473
transform 1 0 4430 0 1 4430
box -12 -8 32 272
use FILL  FILL_7_BUFX2_insert26
timestamp 1701859473
transform 1 0 4250 0 1 2870
box -12 -8 32 272
use FILL  FILL_7_BUFX2_insert27
timestamp 1701859473
transform 1 0 9650 0 1 4950
box -12 -8 32 272
use FILL  FILL_7_BUFX2_insert29
timestamp 1701859473
transform -1 0 1330 0 1 6510
box -12 -8 32 272
use FILL  FILL_7_BUFX2_insert30
timestamp 1701859473
transform -1 0 8830 0 -1 3910
box -12 -8 32 272
use FILL  FILL_7_BUFX2_insert31
timestamp 1701859473
transform -1 0 9610 0 1 3910
box -12 -8 32 272
use FILL  FILL_7_BUFX2_insert32
timestamp 1701859473
transform 1 0 5910 0 -1 3910
box -12 -8 32 272
use FILL  FILL_7_BUFX2_insert33
timestamp 1701859473
transform -1 0 9590 0 -1 4950
box -12 -8 32 272
use FILL  FILL_7_BUFX2_insert34
timestamp 1701859473
transform 1 0 5250 0 1 8590
box -12 -8 32 272
use FILL  FILL_7_BUFX2_insert35
timestamp 1701859473
transform -1 0 6010 0 1 7550
box -12 -8 32 272
use FILL  FILL_7_BUFX2_insert37
timestamp 1701859473
transform -1 0 9630 0 1 8590
box -12 -8 32 272
use FILL  FILL_7_BUFX2_insert49
timestamp 1701859473
transform -1 0 3090 0 1 6510
box -12 -8 32 272
use FILL  FILL_7_BUFX2_insert51
timestamp 1701859473
transform 1 0 3250 0 -1 8590
box -12 -8 32 272
use FILL  FILL_7_BUFX2_insert52
timestamp 1701859473
transform 1 0 3430 0 1 5470
box -12 -8 32 272
use FILL  FILL_7_BUFX2_insert53
timestamp 1701859473
transform -1 0 11270 0 1 9110
box -12 -8 32 272
use FILL  FILL_7_BUFX2_insert54
timestamp 1701859473
transform -1 0 9210 0 1 8590
box -12 -8 32 272
use FILL  FILL_7_BUFX2_insert55
timestamp 1701859473
transform -1 0 9650 0 1 9110
box -12 -8 32 272
use FILL  FILL_7_BUFX2_insert56
timestamp 1701859473
transform -1 0 10310 0 1 9110
box -12 -8 32 272
use FILL  FILL_7_BUFX2_insert58
timestamp 1701859473
transform -1 0 9010 0 1 2870
box -12 -8 32 272
use FILL  FILL_7_BUFX2_insert59
timestamp 1701859473
transform -1 0 7590 0 1 1830
box -12 -8 32 272
use FILL  FILL_7_BUFX2_insert60
timestamp 1701859473
transform 1 0 10930 0 1 1830
box -12 -8 32 272
use FILL  FILL_7_BUFX2_insert61
timestamp 1701859473
transform -1 0 11210 0 1 2870
box -12 -8 32 272
use FILL  FILL_7_BUFX2_insert62
timestamp 1701859473
transform 1 0 2250 0 1 3910
box -12 -8 32 272
use FILL  FILL_7_BUFX2_insert63
timestamp 1701859473
transform 1 0 2170 0 1 3390
box -12 -8 32 272
use FILL  FILL_7_BUFX2_insert64
timestamp 1701859473
transform -1 0 1830 0 1 3910
box -12 -8 32 272
use FILL  FILL_7_BUFX2_insert66
timestamp 1701859473
transform -1 0 4350 0 1 1310
box -12 -8 32 272
use FILL  FILL_7_BUFX2_insert67
timestamp 1701859473
transform -1 0 3650 0 -1 10150
box -12 -8 32 272
use FILL  FILL_7_BUFX2_insert68
timestamp 1701859473
transform -1 0 7210 0 1 2870
box -12 -8 32 272
use FILL  FILL_7_BUFX2_insert69
timestamp 1701859473
transform -1 0 5690 0 -1 3390
box -12 -8 32 272
use FILL  FILL_7_BUFX2_insert70
timestamp 1701859473
transform -1 0 3710 0 -1 1830
box -12 -8 32 272
use FILL  FILL_7_BUFX2_insert71
timestamp 1701859473
transform -1 0 7350 0 1 2350
box -12 -8 32 272
use FILL  FILL_7_BUFX2_insert73
timestamp 1701859473
transform 1 0 3650 0 1 5470
box -12 -8 32 272
use FILL  FILL_7_BUFX2_insert74
timestamp 1701859473
transform 1 0 7610 0 -1 2350
box -12 -8 32 272
use FILL  FILL_7_BUFX2_insert75
timestamp 1701859473
transform 1 0 7630 0 1 2870
box -12 -8 32 272
use FILL  FILL_7_BUFX2_insert76
timestamp 1701859473
transform 1 0 7410 0 1 2870
box -12 -8 32 272
use FILL  FILL_7_BUFX2_insert77
timestamp 1701859473
transform -1 0 3470 0 -1 2870
box -12 -8 32 272
use FILL  FILL_7_BUFX2_insert78
timestamp 1701859473
transform 1 0 1970 0 -1 2870
box -12 -8 32 272
use FILL  FILL_7_BUFX2_insert80
timestamp 1701859473
transform 1 0 2450 0 1 4430
box -12 -8 32 272
use FILL  FILL_7_BUFX2_insert81
timestamp 1701859473
transform -1 0 2050 0 1 3910
box -12 -8 32 272
use FILL  FILL_7_BUFX2_insert82
timestamp 1701859473
transform -1 0 370 0 1 8590
box -12 -8 32 272
use FILL  FILL_7_BUFX2_insert83
timestamp 1701859473
transform 1 0 4250 0 -1 10150
box -12 -8 32 272
use FILL  FILL_7_BUFX2_insert84
timestamp 1701859473
transform 1 0 4210 0 -1 7550
box -12 -8 32 272
use FILL  FILL_7_BUFX2_insert85
timestamp 1701859473
transform -1 0 170 0 -1 6510
box -12 -8 32 272
use FILL  FILL_7_BUFX2_insert86
timestamp 1701859473
transform 1 0 1970 0 -1 10150
box -12 -8 32 272
use FILL  FILL_7_CLKBUF1_insert38
timestamp 1701859473
transform 1 0 2970 0 -1 7550
box -12 -8 32 272
use FILL  FILL_7_CLKBUF1_insert39
timestamp 1701859473
transform -1 0 4770 0 -1 6510
box -12 -8 32 272
use FILL  FILL_7_CLKBUF1_insert40
timestamp 1701859473
transform -1 0 1070 0 -1 4950
box -12 -8 32 272
use FILL  FILL_7_CLKBUF1_insert41
timestamp 1701859473
transform -1 0 10730 0 -1 270
box -12 -8 32 272
use FILL  FILL_7_CLKBUF1_insert42
timestamp 1701859473
transform 1 0 9790 0 -1 4950
box -12 -8 32 272
use FILL  FILL_7_CLKBUF1_insert44
timestamp 1701859473
transform -1 0 10850 0 1 4430
box -12 -8 32 272
use FILL  FILL_7_CLKBUF1_insert45
timestamp 1701859473
transform 1 0 5770 0 -1 6510
box -12 -8 32 272
use FILL  FILL_7_CLKBUF1_insert46
timestamp 1701859473
transform 1 0 4090 0 1 5990
box -12 -8 32 272
use FILL  FILL_7_CLKBUF1_insert47
timestamp 1701859473
transform -1 0 2210 0 1 7550
box -12 -8 32 272
use FILL  FILL_7_CLKBUF1_insert48
timestamp 1701859473
transform -1 0 10890 0 -1 7030
box -12 -8 32 272
<< labels >>
flabel metal1 s 11343 2 11403 2 3 FreeSans 16 270 0 0 gnd
port 0 nsew
flabel metal1 s -63 2 -3 2 7 FreeSans 16 270 0 0 vdd
port 1 nsew
flabel metal2 s 5357 11237 5363 11243 3 FreeSans 16 90 0 0 AB[7]
port 10 nsew
flabel metal2 s 4797 11237 4803 11243 3 FreeSans 16 90 0 0 AB[2]
port 15 nsew
flabel metal2 s 4717 11237 4723 11243 3 FreeSans 16 90 0 0 AB[1]
port 16 nsew
flabel metal2 s 1737 11237 1743 11243 3 FreeSans 16 90 0 0 DI[6]
port 19 nsew
flabel metal2 s 6897 -23 6903 -17 7 FreeSans 16 270 0 0 DI[0]
port 25 nsew
flabel metal2 s 5797 11237 5803 11243 3 FreeSans 16 90 0 0 DO[2]
port 31 nsew
flabel metal2 s 5337 -23 5343 -17 7 FreeSans 16 270 0 0 WE
port 37 nsew
flabel metal3 s 11395 5096 11403 5104 3 FreeSans 16 0 0 0 NMI
port 35 nsew
flabel metal3 s 11395 6076 11403 6084 3 FreeSans 16 0 0 0 IRQ
port 34 nsew
flabel metal3 s 11395 6636 11403 6644 3 FreeSans 16 0 0 0 reset
port 39 nsew
flabel metal3 s 11395 6896 11403 6904 3 FreeSans 16 0 0 0 AB[0]
port 17 nsew
flabel metal2 s 6397 11237 6403 11243 3 FreeSans 16 90 0 0 DO[1]
port 32 nsew
flabel metal2 s 6297 11237 6303 11243 3 FreeSans 16 90 0 0 DO[3]
port 30 nsew
flabel metal2 s 6077 11237 6083 11243 3 FreeSans 16 90 0 0 DO[6]
port 27 nsew
flabel metal2 s 5977 11237 5983 11243 3 FreeSans 16 90 0 0 DI[1]
port 24 nsew
flabel metal2 s 5897 11237 5903 11243 3 FreeSans 16 90 0 0 DO[7]
port 26 nsew
flabel metal2 s 5657 11237 5663 11243 3 FreeSans 16 90 0 0 AB[6]
port 11 nsew
flabel metal2 s 5700 11237 5706 11243 3 FreeSans 16 90 0 0 DO[5]
port 28 nsew
flabel metal2 s 5458 11237 5464 11243 3 FreeSans 16 90 0 0 AB[3]
port 14 nsew
flabel metal2 s 5097 11237 5103 11243 3 FreeSans 16 90 0 0 DO[0]
port 33 nsew
flabel metal2 s 5178 11237 5184 11243 3 FreeSans 16 90 0 0 AB[5]
port 12 nsew
flabel metal2 s 4857 11237 4863 11243 3 FreeSans 16 90 0 0 DO[4]
port 29 nsew
flabel metal2 s 4357 11237 4363 11243 3 FreeSans 16 90 0 0 AB[4]
port 13 nsew
flabel metal2 s 2117 11237 2123 11243 3 FreeSans 16 90 0 0 DI[7]
port 18 nsew
flabel metal2 s 1997 11237 2003 11243 3 FreeSans 16 90 0 0 AB[14]
port 3 nsew
flabel metal2 s 1397 11237 1403 11243 3 FreeSans 16 90 0 0 DI[5]
port 20 nsew
flabel metal2 s 377 11237 383 11243 3 FreeSans 16 90 0 0 DI[3]
port 22 nsew
flabel metal3 s -63 11097 -55 11105 7 FreeSans 16 0 0 0 RDY
port 36 nsew
flabel metal3 s -63 9256 -55 9264 7 FreeSans 16 0 0 0 AB[13]
port 4 nsew
flabel metal3 s -63 9307 -55 9315 7 FreeSans 16 0 0 0 AB[15]
port 2 nsew
flabel metal3 s -63 8716 -55 8724 7 FreeSans 16 0 0 0 AB[12]
port 5 nsew
flabel metal3 s -63 7936 -55 7944 7 FreeSans 16 0 0 0 AB[11]
port 6 nsew
flabel metal3 s -63 7216 -55 7224 7 FreeSans 16 0 0 0 AB[9]
port 8 nsew
flabel metal3 s -63 7156 -55 7164 7 FreeSans 16 0 0 0 DI[4]
port 21 nsew
flabel metal3 s -63 6116 -55 6124 7 FreeSans 16 0 0 0 AB[10]
port 7 nsew
flabel metal3 s -63 5856 -55 5864 7 FreeSans 16 0 0 0 AB[8]
port 9 nsew
flabel metal3 s -63 5296 -55 5304 7 FreeSans 16 0 0 0 DI[2]
port 23 nsew
flabel metal3 s 11395 7156 11403 7164 3 FreeSans 16 0 0 0 clk
port 38 nsew
<< properties >>
string FIXED_BBOX -40 -40 11380 11240
<< end >>
